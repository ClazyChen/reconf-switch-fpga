module SRAM(
  input         clock,
  input         io_w_en,
  input  [7:0]  io_w_addr,
  input  [63:0] io_w_data,
  input  [7:0]  io_r_addr,
  output [63:0] io_r_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mem [0:255]; // @[sram.scala 30:26]
  wire [63:0] mem_io_r_data_MPORT_data; // @[sram.scala 30:26]
  wire [7:0] mem_io_r_data_MPORT_addr; // @[sram.scala 30:26]
  wire [63:0] mem_MPORT_data; // @[sram.scala 30:26]
  wire [7:0] mem_MPORT_addr; // @[sram.scala 30:26]
  wire  mem_MPORT_mask; // @[sram.scala 30:26]
  wire  mem_MPORT_en; // @[sram.scala 30:26]
  reg  mem_io_r_data_MPORT_en_pipe_0;
  reg [7:0] mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_addr = mem_io_r_data_MPORT_addr_pipe_0;
  assign mem_io_r_data_MPORT_data = mem[mem_io_r_data_MPORT_addr]; // @[sram.scala 30:26]
  assign mem_MPORT_data = io_w_data;
  assign mem_MPORT_addr = io_w_addr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_w_en;
  assign io_r_data = mem_io_r_data_MPORT_data; // @[sram.scala 37:24 sram.scala 38:23]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[sram.scala 30:26]
    end
    if (io_w_en) begin
      mem_io_r_data_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      mem_io_r_data_MPORT_en_pipe_0 <= 1'h1;
    end
    if (io_w_en ? 1'h0 : 1'h1) begin
      mem_io_r_data_MPORT_addr_pipe_0 <= io_r_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_r_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_r_data_MPORT_addr_pipe_0 = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ActionReader(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  input         io_hit,
  input  [63:0] io_match_value,
  output [7:0]  io_args_out_0,
  output [7:0]  io_args_out_1,
  output [7:0]  io_args_out_2,
  output [7:0]  io_args_out_3,
  output [7:0]  io_args_out_4,
  output [7:0]  io_args_out_5,
  output [7:0]  io_args_out_6,
  output [31:0] io_vliw_out_0,
  output [31:0] io_vliw_out_1,
  output [31:0] io_vliw_out_2,
  output [31:0] io_vliw_out_3,
  input         io_action_mod_en,
  input  [7:0]  io_action_mod_addr,
  input  [63:0] io_action_mod_data_0,
  input  [63:0] io_action_mod_data_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [63:0] _RAND_116;
`endif // RANDOMIZE_REG_INIT
  wire  sram_0_clock; // @[executor.scala 40:29]
  wire  sram_0_io_w_en; // @[executor.scala 40:29]
  wire [7:0] sram_0_io_w_addr; // @[executor.scala 40:29]
  wire [63:0] sram_0_io_w_data; // @[executor.scala 40:29]
  wire [7:0] sram_0_io_r_addr; // @[executor.scala 40:29]
  wire [63:0] sram_0_io_r_data; // @[executor.scala 40:29]
  wire  sram_1_clock; // @[executor.scala 40:29]
  wire  sram_1_io_w_en; // @[executor.scala 40:29]
  wire [7:0] sram_1_io_w_addr; // @[executor.scala 40:29]
  wire [63:0] sram_1_io_w_data; // @[executor.scala 40:29]
  wire [7:0] sram_1_io_r_addr; // @[executor.scala 40:29]
  wire [63:0] sram_1_io_r_data; // @[executor.scala 40:29]
  reg [7:0] phv_data_0; // @[executor.scala 28:22]
  reg [7:0] phv_data_1; // @[executor.scala 28:22]
  reg [7:0] phv_data_2; // @[executor.scala 28:22]
  reg [7:0] phv_data_3; // @[executor.scala 28:22]
  reg [7:0] phv_data_4; // @[executor.scala 28:22]
  reg [7:0] phv_data_5; // @[executor.scala 28:22]
  reg [7:0] phv_data_6; // @[executor.scala 28:22]
  reg [7:0] phv_data_7; // @[executor.scala 28:22]
  reg [7:0] phv_data_8; // @[executor.scala 28:22]
  reg [7:0] phv_data_9; // @[executor.scala 28:22]
  reg [7:0] phv_data_10; // @[executor.scala 28:22]
  reg [7:0] phv_data_11; // @[executor.scala 28:22]
  reg [7:0] phv_data_12; // @[executor.scala 28:22]
  reg [7:0] phv_data_13; // @[executor.scala 28:22]
  reg [7:0] phv_data_14; // @[executor.scala 28:22]
  reg [7:0] phv_data_15; // @[executor.scala 28:22]
  reg [7:0] phv_data_16; // @[executor.scala 28:22]
  reg [7:0] phv_data_17; // @[executor.scala 28:22]
  reg [7:0] phv_data_18; // @[executor.scala 28:22]
  reg [7:0] phv_data_19; // @[executor.scala 28:22]
  reg [7:0] phv_data_20; // @[executor.scala 28:22]
  reg [7:0] phv_data_21; // @[executor.scala 28:22]
  reg [7:0] phv_data_22; // @[executor.scala 28:22]
  reg [7:0] phv_data_23; // @[executor.scala 28:22]
  reg [7:0] phv_data_24; // @[executor.scala 28:22]
  reg [7:0] phv_data_25; // @[executor.scala 28:22]
  reg [7:0] phv_data_26; // @[executor.scala 28:22]
  reg [7:0] phv_data_27; // @[executor.scala 28:22]
  reg [7:0] phv_data_28; // @[executor.scala 28:22]
  reg [7:0] phv_data_29; // @[executor.scala 28:22]
  reg [7:0] phv_data_30; // @[executor.scala 28:22]
  reg [7:0] phv_data_31; // @[executor.scala 28:22]
  reg [7:0] phv_data_32; // @[executor.scala 28:22]
  reg [7:0] phv_data_33; // @[executor.scala 28:22]
  reg [7:0] phv_data_34; // @[executor.scala 28:22]
  reg [7:0] phv_data_35; // @[executor.scala 28:22]
  reg [7:0] phv_data_36; // @[executor.scala 28:22]
  reg [7:0] phv_data_37; // @[executor.scala 28:22]
  reg [7:0] phv_data_38; // @[executor.scala 28:22]
  reg [7:0] phv_data_39; // @[executor.scala 28:22]
  reg [7:0] phv_data_40; // @[executor.scala 28:22]
  reg [7:0] phv_data_41; // @[executor.scala 28:22]
  reg [7:0] phv_data_42; // @[executor.scala 28:22]
  reg [7:0] phv_data_43; // @[executor.scala 28:22]
  reg [7:0] phv_data_44; // @[executor.scala 28:22]
  reg [7:0] phv_data_45; // @[executor.scala 28:22]
  reg [7:0] phv_data_46; // @[executor.scala 28:22]
  reg [7:0] phv_data_47; // @[executor.scala 28:22]
  reg [7:0] phv_data_48; // @[executor.scala 28:22]
  reg [7:0] phv_data_49; // @[executor.scala 28:22]
  reg [7:0] phv_data_50; // @[executor.scala 28:22]
  reg [7:0] phv_data_51; // @[executor.scala 28:22]
  reg [7:0] phv_data_52; // @[executor.scala 28:22]
  reg [7:0] phv_data_53; // @[executor.scala 28:22]
  reg [7:0] phv_data_54; // @[executor.scala 28:22]
  reg [7:0] phv_data_55; // @[executor.scala 28:22]
  reg [7:0] phv_data_56; // @[executor.scala 28:22]
  reg [7:0] phv_data_57; // @[executor.scala 28:22]
  reg [7:0] phv_data_58; // @[executor.scala 28:22]
  reg [7:0] phv_data_59; // @[executor.scala 28:22]
  reg [7:0] phv_data_60; // @[executor.scala 28:22]
  reg [7:0] phv_data_61; // @[executor.scala 28:22]
  reg [7:0] phv_data_62; // @[executor.scala 28:22]
  reg [7:0] phv_data_63; // @[executor.scala 28:22]
  reg [7:0] phv_data_64; // @[executor.scala 28:22]
  reg [7:0] phv_data_65; // @[executor.scala 28:22]
  reg [7:0] phv_data_66; // @[executor.scala 28:22]
  reg [7:0] phv_data_67; // @[executor.scala 28:22]
  reg [7:0] phv_data_68; // @[executor.scala 28:22]
  reg [7:0] phv_data_69; // @[executor.scala 28:22]
  reg [7:0] phv_data_70; // @[executor.scala 28:22]
  reg [7:0] phv_data_71; // @[executor.scala 28:22]
  reg [7:0] phv_data_72; // @[executor.scala 28:22]
  reg [7:0] phv_data_73; // @[executor.scala 28:22]
  reg [7:0] phv_data_74; // @[executor.scala 28:22]
  reg [7:0] phv_data_75; // @[executor.scala 28:22]
  reg [7:0] phv_data_76; // @[executor.scala 28:22]
  reg [7:0] phv_data_77; // @[executor.scala 28:22]
  reg [7:0] phv_data_78; // @[executor.scala 28:22]
  reg [7:0] phv_data_79; // @[executor.scala 28:22]
  reg [7:0] phv_data_80; // @[executor.scala 28:22]
  reg [7:0] phv_data_81; // @[executor.scala 28:22]
  reg [7:0] phv_data_82; // @[executor.scala 28:22]
  reg [7:0] phv_data_83; // @[executor.scala 28:22]
  reg [7:0] phv_data_84; // @[executor.scala 28:22]
  reg [7:0] phv_data_85; // @[executor.scala 28:22]
  reg [7:0] phv_data_86; // @[executor.scala 28:22]
  reg [7:0] phv_data_87; // @[executor.scala 28:22]
  reg [7:0] phv_data_88; // @[executor.scala 28:22]
  reg [7:0] phv_data_89; // @[executor.scala 28:22]
  reg [7:0] phv_data_90; // @[executor.scala 28:22]
  reg [7:0] phv_data_91; // @[executor.scala 28:22]
  reg [7:0] phv_data_92; // @[executor.scala 28:22]
  reg [7:0] phv_data_93; // @[executor.scala 28:22]
  reg [7:0] phv_data_94; // @[executor.scala 28:22]
  reg [7:0] phv_data_95; // @[executor.scala 28:22]
  reg [15:0] phv_header_0; // @[executor.scala 28:22]
  reg [15:0] phv_header_1; // @[executor.scala 28:22]
  reg [15:0] phv_header_2; // @[executor.scala 28:22]
  reg [15:0] phv_header_3; // @[executor.scala 28:22]
  reg [15:0] phv_header_4; // @[executor.scala 28:22]
  reg [15:0] phv_header_5; // @[executor.scala 28:22]
  reg [15:0] phv_header_6; // @[executor.scala 28:22]
  reg [15:0] phv_header_7; // @[executor.scala 28:22]
  reg [15:0] phv_header_8; // @[executor.scala 28:22]
  reg [15:0] phv_header_9; // @[executor.scala 28:22]
  reg [15:0] phv_header_10; // @[executor.scala 28:22]
  reg [15:0] phv_header_11; // @[executor.scala 28:22]
  reg [15:0] phv_header_12; // @[executor.scala 28:22]
  reg [15:0] phv_header_13; // @[executor.scala 28:22]
  reg [15:0] phv_header_14; // @[executor.scala 28:22]
  reg [15:0] phv_header_15; // @[executor.scala 28:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 28:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 28:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 28:22]
  reg [1:0] phv_next_processor_id; // @[executor.scala 28:22]
  reg [55:0] args; // @[executor.scala 33:23]
  SRAM sram_0 ( // @[executor.scala 40:29]
    .clock(sram_0_clock),
    .io_w_en(sram_0_io_w_en),
    .io_w_addr(sram_0_io_w_addr),
    .io_w_data(sram_0_io_w_data),
    .io_r_addr(sram_0_io_r_addr),
    .io_r_data(sram_0_io_r_data)
  );
  SRAM sram_1 ( // @[executor.scala 40:29]
    .clock(sram_1_clock),
    .io_w_en(sram_1_io_w_en),
    .io_w_addr(sram_1_io_w_addr),
    .io_w_data(sram_1_io_w_data),
    .io_r_addr(sram_1_io_r_addr),
    .io_r_data(sram_1_io_r_data)
  );
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 30:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 30:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 30:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 30:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 30:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 30:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 30:25]
  assign io_args_out_0 = args[55:48]; // @[executor.scala 36:35]
  assign io_args_out_1 = args[47:40]; // @[executor.scala 36:35]
  assign io_args_out_2 = args[39:32]; // @[executor.scala 36:35]
  assign io_args_out_3 = args[31:24]; // @[executor.scala 36:35]
  assign io_args_out_4 = args[23:16]; // @[executor.scala 36:35]
  assign io_args_out_5 = args[15:8]; // @[executor.scala 36:35]
  assign io_args_out_6 = args[7:0]; // @[executor.scala 36:35]
  assign io_vliw_out_0 = sram_0_io_r_data[63:32]; // @[executor.scala 51:93]
  assign io_vliw_out_1 = sram_0_io_r_data[31:0]; // @[executor.scala 51:93]
  assign io_vliw_out_2 = sram_1_io_r_data[63:32]; // @[executor.scala 51:93]
  assign io_vliw_out_3 = sram_1_io_r_data[31:0]; // @[executor.scala 51:93]
  assign sram_0_clock = clock;
  assign sram_0_io_w_en = io_action_mod_en; // @[executor.scala 43:27]
  assign sram_0_io_w_addr = io_action_mod_addr; // @[executor.scala 44:27]
  assign sram_0_io_w_data = io_action_mod_data_0; // @[executor.scala 45:27]
  assign sram_0_io_r_addr = io_hit ? 8'h0 : io_match_value[63:56]; // @[executor.scala 32:28]
  assign sram_1_clock = clock;
  assign sram_1_io_w_en = io_action_mod_en; // @[executor.scala 43:27]
  assign sram_1_io_w_addr = io_action_mod_addr; // @[executor.scala 44:27]
  assign sram_1_io_w_data = io_action_mod_data_1; // @[executor.scala 45:27]
  assign sram_1_io_r_addr = io_hit ? 8'h0 : io_match_value[63:56]; // @[executor.scala 32:28]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 29:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 29:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 29:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 29:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 29:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 29:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 29:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 29:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 29:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 29:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 29:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 29:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 29:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 29:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 29:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 29:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 29:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 29:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 29:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 29:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 29:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 29:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 29:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 29:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 29:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 29:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 29:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 29:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 29:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 29:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 29:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 29:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 29:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 29:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 29:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 29:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 29:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 29:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 29:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 29:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 29:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 29:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 29:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 29:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 29:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 29:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 29:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 29:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 29:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 29:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 29:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 29:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 29:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 29:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 29:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 29:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 29:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 29:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 29:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 29:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 29:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 29:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 29:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 29:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 29:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 29:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 29:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 29:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 29:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 29:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 29:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 29:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 29:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 29:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 29:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 29:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 29:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 29:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 29:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 29:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 29:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 29:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 29:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 29:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 29:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 29:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 29:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 29:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 29:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 29:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 29:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 29:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 29:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 29:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 29:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 29:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 29:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 29:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 29:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 29:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 29:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 29:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 29:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 29:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 29:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 29:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 29:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 29:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 29:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 29:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 29:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 29:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 29:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 29:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 29:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 29:13]
    args <= io_match_value[55:0]; // @[executor.scala 34:31]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {2{`RANDOM}};
  args = _RAND_116[55:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PrimitiveGetOffset(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  output [7:0]  io_args_out_0,
  output [7:0]  io_args_out_1,
  output [7:0]  io_args_out_2,
  output [7:0]  io_args_out_3,
  output [7:0]  io_args_out_4,
  output [7:0]  io_args_out_5,
  output [7:0]  io_args_out_6,
  output [31:0] io_vliw_out_0,
  output [31:0] io_vliw_out_1,
  output [31:0] io_vliw_out_2,
  output [31:0] io_vliw_out_3,
  output [7:0]  io_offset_out_0,
  output [7:0]  io_offset_out_1,
  output [7:0]  io_offset_out_2,
  output [7:0]  io_offset_out_3,
  output [7:0]  io_length_out_0,
  output [7:0]  io_length_out_1,
  output [7:0]  io_length_out_2,
  output [7:0]  io_length_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 69:22]
  reg [7:0] phv_data_1; // @[executor.scala 69:22]
  reg [7:0] phv_data_2; // @[executor.scala 69:22]
  reg [7:0] phv_data_3; // @[executor.scala 69:22]
  reg [7:0] phv_data_4; // @[executor.scala 69:22]
  reg [7:0] phv_data_5; // @[executor.scala 69:22]
  reg [7:0] phv_data_6; // @[executor.scala 69:22]
  reg [7:0] phv_data_7; // @[executor.scala 69:22]
  reg [7:0] phv_data_8; // @[executor.scala 69:22]
  reg [7:0] phv_data_9; // @[executor.scala 69:22]
  reg [7:0] phv_data_10; // @[executor.scala 69:22]
  reg [7:0] phv_data_11; // @[executor.scala 69:22]
  reg [7:0] phv_data_12; // @[executor.scala 69:22]
  reg [7:0] phv_data_13; // @[executor.scala 69:22]
  reg [7:0] phv_data_14; // @[executor.scala 69:22]
  reg [7:0] phv_data_15; // @[executor.scala 69:22]
  reg [7:0] phv_data_16; // @[executor.scala 69:22]
  reg [7:0] phv_data_17; // @[executor.scala 69:22]
  reg [7:0] phv_data_18; // @[executor.scala 69:22]
  reg [7:0] phv_data_19; // @[executor.scala 69:22]
  reg [7:0] phv_data_20; // @[executor.scala 69:22]
  reg [7:0] phv_data_21; // @[executor.scala 69:22]
  reg [7:0] phv_data_22; // @[executor.scala 69:22]
  reg [7:0] phv_data_23; // @[executor.scala 69:22]
  reg [7:0] phv_data_24; // @[executor.scala 69:22]
  reg [7:0] phv_data_25; // @[executor.scala 69:22]
  reg [7:0] phv_data_26; // @[executor.scala 69:22]
  reg [7:0] phv_data_27; // @[executor.scala 69:22]
  reg [7:0] phv_data_28; // @[executor.scala 69:22]
  reg [7:0] phv_data_29; // @[executor.scala 69:22]
  reg [7:0] phv_data_30; // @[executor.scala 69:22]
  reg [7:0] phv_data_31; // @[executor.scala 69:22]
  reg [7:0] phv_data_32; // @[executor.scala 69:22]
  reg [7:0] phv_data_33; // @[executor.scala 69:22]
  reg [7:0] phv_data_34; // @[executor.scala 69:22]
  reg [7:0] phv_data_35; // @[executor.scala 69:22]
  reg [7:0] phv_data_36; // @[executor.scala 69:22]
  reg [7:0] phv_data_37; // @[executor.scala 69:22]
  reg [7:0] phv_data_38; // @[executor.scala 69:22]
  reg [7:0] phv_data_39; // @[executor.scala 69:22]
  reg [7:0] phv_data_40; // @[executor.scala 69:22]
  reg [7:0] phv_data_41; // @[executor.scala 69:22]
  reg [7:0] phv_data_42; // @[executor.scala 69:22]
  reg [7:0] phv_data_43; // @[executor.scala 69:22]
  reg [7:0] phv_data_44; // @[executor.scala 69:22]
  reg [7:0] phv_data_45; // @[executor.scala 69:22]
  reg [7:0] phv_data_46; // @[executor.scala 69:22]
  reg [7:0] phv_data_47; // @[executor.scala 69:22]
  reg [7:0] phv_data_48; // @[executor.scala 69:22]
  reg [7:0] phv_data_49; // @[executor.scala 69:22]
  reg [7:0] phv_data_50; // @[executor.scala 69:22]
  reg [7:0] phv_data_51; // @[executor.scala 69:22]
  reg [7:0] phv_data_52; // @[executor.scala 69:22]
  reg [7:0] phv_data_53; // @[executor.scala 69:22]
  reg [7:0] phv_data_54; // @[executor.scala 69:22]
  reg [7:0] phv_data_55; // @[executor.scala 69:22]
  reg [7:0] phv_data_56; // @[executor.scala 69:22]
  reg [7:0] phv_data_57; // @[executor.scala 69:22]
  reg [7:0] phv_data_58; // @[executor.scala 69:22]
  reg [7:0] phv_data_59; // @[executor.scala 69:22]
  reg [7:0] phv_data_60; // @[executor.scala 69:22]
  reg [7:0] phv_data_61; // @[executor.scala 69:22]
  reg [7:0] phv_data_62; // @[executor.scala 69:22]
  reg [7:0] phv_data_63; // @[executor.scala 69:22]
  reg [7:0] phv_data_64; // @[executor.scala 69:22]
  reg [7:0] phv_data_65; // @[executor.scala 69:22]
  reg [7:0] phv_data_66; // @[executor.scala 69:22]
  reg [7:0] phv_data_67; // @[executor.scala 69:22]
  reg [7:0] phv_data_68; // @[executor.scala 69:22]
  reg [7:0] phv_data_69; // @[executor.scala 69:22]
  reg [7:0] phv_data_70; // @[executor.scala 69:22]
  reg [7:0] phv_data_71; // @[executor.scala 69:22]
  reg [7:0] phv_data_72; // @[executor.scala 69:22]
  reg [7:0] phv_data_73; // @[executor.scala 69:22]
  reg [7:0] phv_data_74; // @[executor.scala 69:22]
  reg [7:0] phv_data_75; // @[executor.scala 69:22]
  reg [7:0] phv_data_76; // @[executor.scala 69:22]
  reg [7:0] phv_data_77; // @[executor.scala 69:22]
  reg [7:0] phv_data_78; // @[executor.scala 69:22]
  reg [7:0] phv_data_79; // @[executor.scala 69:22]
  reg [7:0] phv_data_80; // @[executor.scala 69:22]
  reg [7:0] phv_data_81; // @[executor.scala 69:22]
  reg [7:0] phv_data_82; // @[executor.scala 69:22]
  reg [7:0] phv_data_83; // @[executor.scala 69:22]
  reg [7:0] phv_data_84; // @[executor.scala 69:22]
  reg [7:0] phv_data_85; // @[executor.scala 69:22]
  reg [7:0] phv_data_86; // @[executor.scala 69:22]
  reg [7:0] phv_data_87; // @[executor.scala 69:22]
  reg [7:0] phv_data_88; // @[executor.scala 69:22]
  reg [7:0] phv_data_89; // @[executor.scala 69:22]
  reg [7:0] phv_data_90; // @[executor.scala 69:22]
  reg [7:0] phv_data_91; // @[executor.scala 69:22]
  reg [7:0] phv_data_92; // @[executor.scala 69:22]
  reg [7:0] phv_data_93; // @[executor.scala 69:22]
  reg [7:0] phv_data_94; // @[executor.scala 69:22]
  reg [7:0] phv_data_95; // @[executor.scala 69:22]
  reg [15:0] phv_header_0; // @[executor.scala 69:22]
  reg [15:0] phv_header_1; // @[executor.scala 69:22]
  reg [15:0] phv_header_2; // @[executor.scala 69:22]
  reg [15:0] phv_header_3; // @[executor.scala 69:22]
  reg [15:0] phv_header_4; // @[executor.scala 69:22]
  reg [15:0] phv_header_5; // @[executor.scala 69:22]
  reg [15:0] phv_header_6; // @[executor.scala 69:22]
  reg [15:0] phv_header_7; // @[executor.scala 69:22]
  reg [15:0] phv_header_8; // @[executor.scala 69:22]
  reg [15:0] phv_header_9; // @[executor.scala 69:22]
  reg [15:0] phv_header_10; // @[executor.scala 69:22]
  reg [15:0] phv_header_11; // @[executor.scala 69:22]
  reg [15:0] phv_header_12; // @[executor.scala 69:22]
  reg [15:0] phv_header_13; // @[executor.scala 69:22]
  reg [15:0] phv_header_14; // @[executor.scala 69:22]
  reg [15:0] phv_header_15; // @[executor.scala 69:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 69:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 69:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 69:22]
  reg [1:0] phv_next_processor_id; // @[executor.scala 69:22]
  reg [7:0] args_0; // @[executor.scala 73:23]
  reg [7:0] args_1; // @[executor.scala 73:23]
  reg [7:0] args_2; // @[executor.scala 73:23]
  reg [7:0] args_3; // @[executor.scala 73:23]
  reg [7:0] args_4; // @[executor.scala 73:23]
  reg [7:0] args_5; // @[executor.scala 73:23]
  reg [7:0] args_6; // @[executor.scala 73:23]
  reg [31:0] vliw_0; // @[executor.scala 77:23]
  reg [31:0] vliw_1; // @[executor.scala 77:23]
  reg [31:0] vliw_2; // @[executor.scala 77:23]
  reg [31:0] vliw_3; // @[executor.scala 77:23]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1 = vliw_0[27:14]; // @[primitive.scala 10:44]
  wire [13:0] parameter_2 = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire  is_addi = 4'h8 == opcode; // @[executor.scala 86:48]
  wire  is_copy = 4'h9 == opcode; // @[executor.scala 87:48]
  wire [13:0] dst = is_addi ? parameter_1 : parameter_2; // @[executor.scala 90:30]
  wire [3:0] header_id = dst[13:10]; // @[primitive.scala 27:52]
  wire [4:0] internal_offset = dst[9:5]; // @[primitive.scala 28:52]
  wire [4:0] length = dst[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_1 = 4'h1 == header_id ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_2 = 4'h2 == header_id ? phv_header_2 : _GEN_1; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_3 = 4'h3 == header_id ? phv_header_3 : _GEN_2; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_4 = 4'h4 == header_id ? phv_header_4 : _GEN_3; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_5 = 4'h5 == header_id ? phv_header_5 : _GEN_4; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_6 = 4'h6 == header_id ? phv_header_6 : _GEN_5; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_7 = 4'h7 == header_id ? phv_header_7 : _GEN_6; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_8 = 4'h8 == header_id ? phv_header_8 : _GEN_7; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_9 = 4'h9 == header_id ? phv_header_9 : _GEN_8; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_10 = 4'ha == header_id ? phv_header_10 : _GEN_9; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_11 = 4'hb == header_id ? phv_header_11 : _GEN_10; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_12 = 4'hc == header_id ? phv_header_12 : _GEN_11; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_13 = 4'hd == header_id ? phv_header_13 : _GEN_12; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_14 = 4'he == header_id ? phv_header_14 : _GEN_13; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_15 = 4'hf == header_id ? phv_header_15 : _GEN_14; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] header_offset = _GEN_15[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_72 = {{3'd0}, internal_offset}; // @[executor.scala 95:53]
  wire [7:0] offset = header_offset + _GEN_72; // @[executor.scala 95:53]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_1 = vliw_1[27:14]; // @[primitive.scala 10:44]
  wire [13:0] parameter_2_1 = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire  is_addi_1 = 4'h8 == opcode_1; // @[executor.scala 86:48]
  wire  is_copy_1 = 4'h9 == opcode_1; // @[executor.scala 87:48]
  wire [13:0] dst_1 = is_addi_1 ? parameter_1_1 : parameter_2_1; // @[executor.scala 90:30]
  wire [3:0] header_id_1 = dst_1[13:10]; // @[primitive.scala 27:52]
  wire [4:0] internal_offset_1 = dst_1[9:5]; // @[primitive.scala 28:52]
  wire [4:0] length_1 = dst_1[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_19 = 4'h1 == header_id_1 ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_20 = 4'h2 == header_id_1 ? phv_header_2 : _GEN_19; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_21 = 4'h3 == header_id_1 ? phv_header_3 : _GEN_20; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_22 = 4'h4 == header_id_1 ? phv_header_4 : _GEN_21; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_23 = 4'h5 == header_id_1 ? phv_header_5 : _GEN_22; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_24 = 4'h6 == header_id_1 ? phv_header_6 : _GEN_23; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_25 = 4'h7 == header_id_1 ? phv_header_7 : _GEN_24; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_26 = 4'h8 == header_id_1 ? phv_header_8 : _GEN_25; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_27 = 4'h9 == header_id_1 ? phv_header_9 : _GEN_26; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_28 = 4'ha == header_id_1 ? phv_header_10 : _GEN_27; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_29 = 4'hb == header_id_1 ? phv_header_11 : _GEN_28; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_30 = 4'hc == header_id_1 ? phv_header_12 : _GEN_29; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_31 = 4'hd == header_id_1 ? phv_header_13 : _GEN_30; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_32 = 4'he == header_id_1 ? phv_header_14 : _GEN_31; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_33 = 4'hf == header_id_1 ? phv_header_15 : _GEN_32; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] header_offset_1 = _GEN_33[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_73 = {{3'd0}, internal_offset_1}; // @[executor.scala 95:53]
  wire [7:0] offset_1 = header_offset_1 + _GEN_73; // @[executor.scala 95:53]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_2 = vliw_2[27:14]; // @[primitive.scala 10:44]
  wire [13:0] parameter_2_2 = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire  is_addi_2 = 4'h8 == opcode_2; // @[executor.scala 86:48]
  wire  is_copy_2 = 4'h9 == opcode_2; // @[executor.scala 87:48]
  wire [13:0] dst_2 = is_addi_2 ? parameter_1_2 : parameter_2_2; // @[executor.scala 90:30]
  wire [3:0] header_id_2 = dst_2[13:10]; // @[primitive.scala 27:52]
  wire [4:0] internal_offset_2 = dst_2[9:5]; // @[primitive.scala 28:52]
  wire [4:0] length_2 = dst_2[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_37 = 4'h1 == header_id_2 ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_38 = 4'h2 == header_id_2 ? phv_header_2 : _GEN_37; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_39 = 4'h3 == header_id_2 ? phv_header_3 : _GEN_38; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_40 = 4'h4 == header_id_2 ? phv_header_4 : _GEN_39; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_41 = 4'h5 == header_id_2 ? phv_header_5 : _GEN_40; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_42 = 4'h6 == header_id_2 ? phv_header_6 : _GEN_41; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_43 = 4'h7 == header_id_2 ? phv_header_7 : _GEN_42; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_44 = 4'h8 == header_id_2 ? phv_header_8 : _GEN_43; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_45 = 4'h9 == header_id_2 ? phv_header_9 : _GEN_44; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_46 = 4'ha == header_id_2 ? phv_header_10 : _GEN_45; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_47 = 4'hb == header_id_2 ? phv_header_11 : _GEN_46; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_48 = 4'hc == header_id_2 ? phv_header_12 : _GEN_47; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_49 = 4'hd == header_id_2 ? phv_header_13 : _GEN_48; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_50 = 4'he == header_id_2 ? phv_header_14 : _GEN_49; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_51 = 4'hf == header_id_2 ? phv_header_15 : _GEN_50; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] header_offset_2 = _GEN_51[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_74 = {{3'd0}, internal_offset_2}; // @[executor.scala 95:53]
  wire [7:0] offset_2 = header_offset_2 + _GEN_74; // @[executor.scala 95:53]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_3 = vliw_3[27:14]; // @[primitive.scala 10:44]
  wire [13:0] parameter_2_3 = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire  is_addi_3 = 4'h8 == opcode_3; // @[executor.scala 86:48]
  wire  is_copy_3 = 4'h9 == opcode_3; // @[executor.scala 87:48]
  wire [13:0] dst_3 = is_addi_3 ? parameter_1_3 : parameter_2_3; // @[executor.scala 90:30]
  wire [3:0] header_id_3 = dst_3[13:10]; // @[primitive.scala 27:52]
  wire [4:0] internal_offset_3 = dst_3[9:5]; // @[primitive.scala 28:52]
  wire [4:0] length_3 = dst_3[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_55 = 4'h1 == header_id_3 ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_56 = 4'h2 == header_id_3 ? phv_header_2 : _GEN_55; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_57 = 4'h3 == header_id_3 ? phv_header_3 : _GEN_56; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_58 = 4'h4 == header_id_3 ? phv_header_4 : _GEN_57; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_59 = 4'h5 == header_id_3 ? phv_header_5 : _GEN_58; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_60 = 4'h6 == header_id_3 ? phv_header_6 : _GEN_59; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_61 = 4'h7 == header_id_3 ? phv_header_7 : _GEN_60; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_62 = 4'h8 == header_id_3 ? phv_header_8 : _GEN_61; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_63 = 4'h9 == header_id_3 ? phv_header_9 : _GEN_62; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_64 = 4'ha == header_id_3 ? phv_header_10 : _GEN_63; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_65 = 4'hb == header_id_3 ? phv_header_11 : _GEN_64; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_66 = 4'hc == header_id_3 ? phv_header_12 : _GEN_65; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_67 = 4'hd == header_id_3 ? phv_header_13 : _GEN_66; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_68 = 4'he == header_id_3 ? phv_header_14 : _GEN_67; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_69 = 4'hf == header_id_3 ? phv_header_15 : _GEN_68; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] header_offset_3 = _GEN_69[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_75 = {{3'd0}, internal_offset_3}; // @[executor.scala 95:53]
  wire [7:0] offset_3 = header_offset_3 + _GEN_75; // @[executor.scala 95:53]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 71:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 71:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 71:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 71:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 71:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 71:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 71:25]
  assign io_args_out_0 = args_0; // @[executor.scala 75:21]
  assign io_args_out_1 = args_1; // @[executor.scala 75:21]
  assign io_args_out_2 = args_2; // @[executor.scala 75:21]
  assign io_args_out_3 = args_3; // @[executor.scala 75:21]
  assign io_args_out_4 = args_4; // @[executor.scala 75:21]
  assign io_args_out_5 = args_5; // @[executor.scala 75:21]
  assign io_args_out_6 = args_6; // @[executor.scala 75:21]
  assign io_vliw_out_0 = vliw_0; // @[executor.scala 79:21]
  assign io_vliw_out_1 = vliw_1; // @[executor.scala 79:21]
  assign io_vliw_out_2 = vliw_2; // @[executor.scala 79:21]
  assign io_vliw_out_3 = vliw_3; // @[executor.scala 79:21]
  assign io_offset_out_0 = is_addi | is_copy ? offset : 8'h0; // @[executor.scala 89:39 executor.scala 96:37 executor.scala 99:37]
  assign io_offset_out_1 = is_addi_1 | is_copy_1 ? offset_1 : 8'h0; // @[executor.scala 89:39 executor.scala 96:37 executor.scala 99:37]
  assign io_offset_out_2 = is_addi_2 | is_copy_2 ? offset_2 : 8'h0; // @[executor.scala 89:39 executor.scala 96:37 executor.scala 99:37]
  assign io_offset_out_3 = is_addi_3 | is_copy_3 ? offset_3 : 8'h0; // @[executor.scala 89:39 executor.scala 96:37 executor.scala 99:37]
  assign io_length_out_0 = is_addi | is_copy ? {{3'd0}, length} : 8'h0; // @[executor.scala 89:39 executor.scala 97:37 executor.scala 100:37]
  assign io_length_out_1 = is_addi_1 | is_copy_1 ? {{3'd0}, length_1} : 8'h0; // @[executor.scala 89:39 executor.scala 97:37 executor.scala 100:37]
  assign io_length_out_2 = is_addi_2 | is_copy_2 ? {{3'd0}, length_2} : 8'h0; // @[executor.scala 89:39 executor.scala 97:37 executor.scala 100:37]
  assign io_length_out_3 = is_addi_3 | is_copy_3 ? {{3'd0}, length_3} : 8'h0; // @[executor.scala 89:39 executor.scala 97:37 executor.scala 100:37]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 70:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 70:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 70:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 70:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 70:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 70:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 70:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 70:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 70:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 70:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 70:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 70:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 70:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 70:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 70:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 70:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 70:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 70:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 70:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 70:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 70:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 70:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 70:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 70:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 70:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 70:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 70:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 70:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 70:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 70:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 70:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 70:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 70:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 70:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 70:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 70:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 70:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 70:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 70:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 70:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 70:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 70:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 70:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 70:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 70:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 70:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 70:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 70:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 70:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 70:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 70:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 70:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 70:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 70:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 70:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 70:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 70:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 70:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 70:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 70:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 70:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 70:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 70:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 70:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 70:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 70:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 70:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 70:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 70:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 70:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 70:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 70:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 70:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 70:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 70:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 70:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 70:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 70:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 70:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 70:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 70:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 70:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 70:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 70:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 70:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 70:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 70:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 70:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 70:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 70:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 70:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 70:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 70:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 70:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 70:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 70:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 70:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 70:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 70:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 70:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 70:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 70:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 70:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 70:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 70:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 70:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 70:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 70:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 70:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 70:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 70:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 70:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 70:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 70:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 70:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 70:13]
    args_0 <= io_args_in_0; // @[executor.scala 74:14]
    args_1 <= io_args_in_1; // @[executor.scala 74:14]
    args_2 <= io_args_in_2; // @[executor.scala 74:14]
    args_3 <= io_args_in_3; // @[executor.scala 74:14]
    args_4 <= io_args_in_4; // @[executor.scala 74:14]
    args_5 <= io_args_in_5; // @[executor.scala 74:14]
    args_6 <= io_args_in_6; // @[executor.scala 74:14]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 78:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 78:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 78:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 78:14]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  args_0 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  args_1 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  args_2 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  args_3 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  args_4 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  args_5 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  args_6 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  vliw_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  vliw_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  vliw_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  vliw_3 = _RAND_126[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PrimitiveGetSource(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [7:0]  io_offset_in_0,
  input  [7:0]  io_offset_in_1,
  input  [7:0]  io_offset_in_2,
  input  [7:0]  io_offset_in_3,
  input  [7:0]  io_length_in_0,
  input  [7:0]  io_length_in_1,
  input  [7:0]  io_length_in_2,
  input  [7:0]  io_length_in_3,
  output [31:0] io_vliw_out_0,
  output [31:0] io_vliw_out_1,
  output [31:0] io_vliw_out_2,
  output [31:0] io_vliw_out_3,
  output [63:0] io_field_out_0,
  output [63:0] io_field_out_1,
  output [63:0] io_field_out_2,
  output [63:0] io_field_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 119:22]
  reg [7:0] phv_data_1; // @[executor.scala 119:22]
  reg [7:0] phv_data_2; // @[executor.scala 119:22]
  reg [7:0] phv_data_3; // @[executor.scala 119:22]
  reg [7:0] phv_data_4; // @[executor.scala 119:22]
  reg [7:0] phv_data_5; // @[executor.scala 119:22]
  reg [7:0] phv_data_6; // @[executor.scala 119:22]
  reg [7:0] phv_data_7; // @[executor.scala 119:22]
  reg [7:0] phv_data_8; // @[executor.scala 119:22]
  reg [7:0] phv_data_9; // @[executor.scala 119:22]
  reg [7:0] phv_data_10; // @[executor.scala 119:22]
  reg [7:0] phv_data_11; // @[executor.scala 119:22]
  reg [7:0] phv_data_12; // @[executor.scala 119:22]
  reg [7:0] phv_data_13; // @[executor.scala 119:22]
  reg [7:0] phv_data_14; // @[executor.scala 119:22]
  reg [7:0] phv_data_15; // @[executor.scala 119:22]
  reg [7:0] phv_data_16; // @[executor.scala 119:22]
  reg [7:0] phv_data_17; // @[executor.scala 119:22]
  reg [7:0] phv_data_18; // @[executor.scala 119:22]
  reg [7:0] phv_data_19; // @[executor.scala 119:22]
  reg [7:0] phv_data_20; // @[executor.scala 119:22]
  reg [7:0] phv_data_21; // @[executor.scala 119:22]
  reg [7:0] phv_data_22; // @[executor.scala 119:22]
  reg [7:0] phv_data_23; // @[executor.scala 119:22]
  reg [7:0] phv_data_24; // @[executor.scala 119:22]
  reg [7:0] phv_data_25; // @[executor.scala 119:22]
  reg [7:0] phv_data_26; // @[executor.scala 119:22]
  reg [7:0] phv_data_27; // @[executor.scala 119:22]
  reg [7:0] phv_data_28; // @[executor.scala 119:22]
  reg [7:0] phv_data_29; // @[executor.scala 119:22]
  reg [7:0] phv_data_30; // @[executor.scala 119:22]
  reg [7:0] phv_data_31; // @[executor.scala 119:22]
  reg [7:0] phv_data_32; // @[executor.scala 119:22]
  reg [7:0] phv_data_33; // @[executor.scala 119:22]
  reg [7:0] phv_data_34; // @[executor.scala 119:22]
  reg [7:0] phv_data_35; // @[executor.scala 119:22]
  reg [7:0] phv_data_36; // @[executor.scala 119:22]
  reg [7:0] phv_data_37; // @[executor.scala 119:22]
  reg [7:0] phv_data_38; // @[executor.scala 119:22]
  reg [7:0] phv_data_39; // @[executor.scala 119:22]
  reg [7:0] phv_data_40; // @[executor.scala 119:22]
  reg [7:0] phv_data_41; // @[executor.scala 119:22]
  reg [7:0] phv_data_42; // @[executor.scala 119:22]
  reg [7:0] phv_data_43; // @[executor.scala 119:22]
  reg [7:0] phv_data_44; // @[executor.scala 119:22]
  reg [7:0] phv_data_45; // @[executor.scala 119:22]
  reg [7:0] phv_data_46; // @[executor.scala 119:22]
  reg [7:0] phv_data_47; // @[executor.scala 119:22]
  reg [7:0] phv_data_48; // @[executor.scala 119:22]
  reg [7:0] phv_data_49; // @[executor.scala 119:22]
  reg [7:0] phv_data_50; // @[executor.scala 119:22]
  reg [7:0] phv_data_51; // @[executor.scala 119:22]
  reg [7:0] phv_data_52; // @[executor.scala 119:22]
  reg [7:0] phv_data_53; // @[executor.scala 119:22]
  reg [7:0] phv_data_54; // @[executor.scala 119:22]
  reg [7:0] phv_data_55; // @[executor.scala 119:22]
  reg [7:0] phv_data_56; // @[executor.scala 119:22]
  reg [7:0] phv_data_57; // @[executor.scala 119:22]
  reg [7:0] phv_data_58; // @[executor.scala 119:22]
  reg [7:0] phv_data_59; // @[executor.scala 119:22]
  reg [7:0] phv_data_60; // @[executor.scala 119:22]
  reg [7:0] phv_data_61; // @[executor.scala 119:22]
  reg [7:0] phv_data_62; // @[executor.scala 119:22]
  reg [7:0] phv_data_63; // @[executor.scala 119:22]
  reg [7:0] phv_data_64; // @[executor.scala 119:22]
  reg [7:0] phv_data_65; // @[executor.scala 119:22]
  reg [7:0] phv_data_66; // @[executor.scala 119:22]
  reg [7:0] phv_data_67; // @[executor.scala 119:22]
  reg [7:0] phv_data_68; // @[executor.scala 119:22]
  reg [7:0] phv_data_69; // @[executor.scala 119:22]
  reg [7:0] phv_data_70; // @[executor.scala 119:22]
  reg [7:0] phv_data_71; // @[executor.scala 119:22]
  reg [7:0] phv_data_72; // @[executor.scala 119:22]
  reg [7:0] phv_data_73; // @[executor.scala 119:22]
  reg [7:0] phv_data_74; // @[executor.scala 119:22]
  reg [7:0] phv_data_75; // @[executor.scala 119:22]
  reg [7:0] phv_data_76; // @[executor.scala 119:22]
  reg [7:0] phv_data_77; // @[executor.scala 119:22]
  reg [7:0] phv_data_78; // @[executor.scala 119:22]
  reg [7:0] phv_data_79; // @[executor.scala 119:22]
  reg [7:0] phv_data_80; // @[executor.scala 119:22]
  reg [7:0] phv_data_81; // @[executor.scala 119:22]
  reg [7:0] phv_data_82; // @[executor.scala 119:22]
  reg [7:0] phv_data_83; // @[executor.scala 119:22]
  reg [7:0] phv_data_84; // @[executor.scala 119:22]
  reg [7:0] phv_data_85; // @[executor.scala 119:22]
  reg [7:0] phv_data_86; // @[executor.scala 119:22]
  reg [7:0] phv_data_87; // @[executor.scala 119:22]
  reg [7:0] phv_data_88; // @[executor.scala 119:22]
  reg [7:0] phv_data_89; // @[executor.scala 119:22]
  reg [7:0] phv_data_90; // @[executor.scala 119:22]
  reg [7:0] phv_data_91; // @[executor.scala 119:22]
  reg [7:0] phv_data_92; // @[executor.scala 119:22]
  reg [7:0] phv_data_93; // @[executor.scala 119:22]
  reg [7:0] phv_data_94; // @[executor.scala 119:22]
  reg [7:0] phv_data_95; // @[executor.scala 119:22]
  reg [15:0] phv_header_0; // @[executor.scala 119:22]
  reg [15:0] phv_header_1; // @[executor.scala 119:22]
  reg [15:0] phv_header_2; // @[executor.scala 119:22]
  reg [15:0] phv_header_3; // @[executor.scala 119:22]
  reg [15:0] phv_header_4; // @[executor.scala 119:22]
  reg [15:0] phv_header_5; // @[executor.scala 119:22]
  reg [15:0] phv_header_6; // @[executor.scala 119:22]
  reg [15:0] phv_header_7; // @[executor.scala 119:22]
  reg [15:0] phv_header_8; // @[executor.scala 119:22]
  reg [15:0] phv_header_9; // @[executor.scala 119:22]
  reg [15:0] phv_header_10; // @[executor.scala 119:22]
  reg [15:0] phv_header_11; // @[executor.scala 119:22]
  reg [15:0] phv_header_12; // @[executor.scala 119:22]
  reg [15:0] phv_header_13; // @[executor.scala 119:22]
  reg [15:0] phv_header_14; // @[executor.scala 119:22]
  reg [15:0] phv_header_15; // @[executor.scala 119:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 119:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 119:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 119:22]
  reg [1:0] phv_next_processor_id; // @[executor.scala 119:22]
  reg [7:0] args_0; // @[executor.scala 123:23]
  reg [7:0] args_1; // @[executor.scala 123:23]
  reg [7:0] args_2; // @[executor.scala 123:23]
  reg [7:0] args_3; // @[executor.scala 123:23]
  reg [7:0] args_4; // @[executor.scala 123:23]
  reg [7:0] args_5; // @[executor.scala 123:23]
  reg [7:0] args_6; // @[executor.scala 123:23]
  reg [31:0] vliw_0; // @[executor.scala 126:23]
  reg [31:0] vliw_1; // @[executor.scala 126:23]
  reg [31:0] vliw_2; // @[executor.scala 126:23]
  reg [31:0] vliw_3; // @[executor.scala 126:23]
  reg [7:0] offset_0; // @[executor.scala 130:25]
  reg [7:0] offset_1; // @[executor.scala 130:25]
  reg [7:0] offset_2; // @[executor.scala 130:25]
  reg [7:0] offset_3; // @[executor.scala 130:25]
  reg [7:0] length_0; // @[executor.scala 131:25]
  reg [7:0] length_1; // @[executor.scala 131:25]
  reg [7:0] length_2; // @[executor.scala 131:25]
  reg [7:0] length_3; // @[executor.scala 131:25]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_0_lo = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire  from_header = length_0 != 8'h0; // @[executor.scala 141:41]
  wire [8:0] _total_offset_T = {{1'd0}, offset_0}; // @[executor.scala 148:53]
  wire [7:0] total_offset = _total_offset_T[7:0]; // @[executor.scala 148:53]
  wire [7:0] _GEN_1 = 7'h1 == total_offset[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2 = 7'h2 == total_offset[6:0] ? phv_data_2 : _GEN_1; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3 = 7'h3 == total_offset[6:0] ? phv_data_3 : _GEN_2; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_4 = 7'h4 == total_offset[6:0] ? phv_data_4 : _GEN_3; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_5 = 7'h5 == total_offset[6:0] ? phv_data_5 : _GEN_4; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_6 = 7'h6 == total_offset[6:0] ? phv_data_6 : _GEN_5; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_7 = 7'h7 == total_offset[6:0] ? phv_data_7 : _GEN_6; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_8 = 7'h8 == total_offset[6:0] ? phv_data_8 : _GEN_7; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_9 = 7'h9 == total_offset[6:0] ? phv_data_9 : _GEN_8; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_10 = 7'ha == total_offset[6:0] ? phv_data_10 : _GEN_9; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_11 = 7'hb == total_offset[6:0] ? phv_data_11 : _GEN_10; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_12 = 7'hc == total_offset[6:0] ? phv_data_12 : _GEN_11; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_13 = 7'hd == total_offset[6:0] ? phv_data_13 : _GEN_12; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_14 = 7'he == total_offset[6:0] ? phv_data_14 : _GEN_13; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_15 = 7'hf == total_offset[6:0] ? phv_data_15 : _GEN_14; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_16 = 7'h10 == total_offset[6:0] ? phv_data_16 : _GEN_15; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_17 = 7'h11 == total_offset[6:0] ? phv_data_17 : _GEN_16; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_18 = 7'h12 == total_offset[6:0] ? phv_data_18 : _GEN_17; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_19 = 7'h13 == total_offset[6:0] ? phv_data_19 : _GEN_18; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_20 = 7'h14 == total_offset[6:0] ? phv_data_20 : _GEN_19; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_21 = 7'h15 == total_offset[6:0] ? phv_data_21 : _GEN_20; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_22 = 7'h16 == total_offset[6:0] ? phv_data_22 : _GEN_21; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_23 = 7'h17 == total_offset[6:0] ? phv_data_23 : _GEN_22; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_24 = 7'h18 == total_offset[6:0] ? phv_data_24 : _GEN_23; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_25 = 7'h19 == total_offset[6:0] ? phv_data_25 : _GEN_24; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_26 = 7'h1a == total_offset[6:0] ? phv_data_26 : _GEN_25; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_27 = 7'h1b == total_offset[6:0] ? phv_data_27 : _GEN_26; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_28 = 7'h1c == total_offset[6:0] ? phv_data_28 : _GEN_27; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_29 = 7'h1d == total_offset[6:0] ? phv_data_29 : _GEN_28; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_30 = 7'h1e == total_offset[6:0] ? phv_data_30 : _GEN_29; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_31 = 7'h1f == total_offset[6:0] ? phv_data_31 : _GEN_30; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_32 = 7'h20 == total_offset[6:0] ? phv_data_32 : _GEN_31; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_33 = 7'h21 == total_offset[6:0] ? phv_data_33 : _GEN_32; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_34 = 7'h22 == total_offset[6:0] ? phv_data_34 : _GEN_33; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_35 = 7'h23 == total_offset[6:0] ? phv_data_35 : _GEN_34; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_36 = 7'h24 == total_offset[6:0] ? phv_data_36 : _GEN_35; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_37 = 7'h25 == total_offset[6:0] ? phv_data_37 : _GEN_36; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_38 = 7'h26 == total_offset[6:0] ? phv_data_38 : _GEN_37; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_39 = 7'h27 == total_offset[6:0] ? phv_data_39 : _GEN_38; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_40 = 7'h28 == total_offset[6:0] ? phv_data_40 : _GEN_39; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_41 = 7'h29 == total_offset[6:0] ? phv_data_41 : _GEN_40; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_42 = 7'h2a == total_offset[6:0] ? phv_data_42 : _GEN_41; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_43 = 7'h2b == total_offset[6:0] ? phv_data_43 : _GEN_42; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_44 = 7'h2c == total_offset[6:0] ? phv_data_44 : _GEN_43; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_45 = 7'h2d == total_offset[6:0] ? phv_data_45 : _GEN_44; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_46 = 7'h2e == total_offset[6:0] ? phv_data_46 : _GEN_45; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_47 = 7'h2f == total_offset[6:0] ? phv_data_47 : _GEN_46; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_48 = 7'h30 == total_offset[6:0] ? phv_data_48 : _GEN_47; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_49 = 7'h31 == total_offset[6:0] ? phv_data_49 : _GEN_48; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_50 = 7'h32 == total_offset[6:0] ? phv_data_50 : _GEN_49; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_51 = 7'h33 == total_offset[6:0] ? phv_data_51 : _GEN_50; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_52 = 7'h34 == total_offset[6:0] ? phv_data_52 : _GEN_51; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_53 = 7'h35 == total_offset[6:0] ? phv_data_53 : _GEN_52; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_54 = 7'h36 == total_offset[6:0] ? phv_data_54 : _GEN_53; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_55 = 7'h37 == total_offset[6:0] ? phv_data_55 : _GEN_54; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_56 = 7'h38 == total_offset[6:0] ? phv_data_56 : _GEN_55; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_57 = 7'h39 == total_offset[6:0] ? phv_data_57 : _GEN_56; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_58 = 7'h3a == total_offset[6:0] ? phv_data_58 : _GEN_57; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_59 = 7'h3b == total_offset[6:0] ? phv_data_59 : _GEN_58; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_60 = 7'h3c == total_offset[6:0] ? phv_data_60 : _GEN_59; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_61 = 7'h3d == total_offset[6:0] ? phv_data_61 : _GEN_60; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_62 = 7'h3e == total_offset[6:0] ? phv_data_62 : _GEN_61; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_63 = 7'h3f == total_offset[6:0] ? phv_data_63 : _GEN_62; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_64 = 7'h40 == total_offset[6:0] ? phv_data_64 : _GEN_63; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_65 = 7'h41 == total_offset[6:0] ? phv_data_65 : _GEN_64; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_66 = 7'h42 == total_offset[6:0] ? phv_data_66 : _GEN_65; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_67 = 7'h43 == total_offset[6:0] ? phv_data_67 : _GEN_66; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_68 = 7'h44 == total_offset[6:0] ? phv_data_68 : _GEN_67; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_69 = 7'h45 == total_offset[6:0] ? phv_data_69 : _GEN_68; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_70 = 7'h46 == total_offset[6:0] ? phv_data_70 : _GEN_69; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_71 = 7'h47 == total_offset[6:0] ? phv_data_71 : _GEN_70; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_72 = 7'h48 == total_offset[6:0] ? phv_data_72 : _GEN_71; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_73 = 7'h49 == total_offset[6:0] ? phv_data_73 : _GEN_72; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_74 = 7'h4a == total_offset[6:0] ? phv_data_74 : _GEN_73; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_75 = 7'h4b == total_offset[6:0] ? phv_data_75 : _GEN_74; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_76 = 7'h4c == total_offset[6:0] ? phv_data_76 : _GEN_75; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_77 = 7'h4d == total_offset[6:0] ? phv_data_77 : _GEN_76; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_78 = 7'h4e == total_offset[6:0] ? phv_data_78 : _GEN_77; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_79 = 7'h4f == total_offset[6:0] ? phv_data_79 : _GEN_78; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_80 = 7'h50 == total_offset[6:0] ? phv_data_80 : _GEN_79; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_81 = 7'h51 == total_offset[6:0] ? phv_data_81 : _GEN_80; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_82 = 7'h52 == total_offset[6:0] ? phv_data_82 : _GEN_81; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_83 = 7'h53 == total_offset[6:0] ? phv_data_83 : _GEN_82; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_84 = 7'h54 == total_offset[6:0] ? phv_data_84 : _GEN_83; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_85 = 7'h55 == total_offset[6:0] ? phv_data_85 : _GEN_84; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_86 = 7'h56 == total_offset[6:0] ? phv_data_86 : _GEN_85; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_87 = 7'h57 == total_offset[6:0] ? phv_data_87 : _GEN_86; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_88 = 7'h58 == total_offset[6:0] ? phv_data_88 : _GEN_87; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_89 = 7'h59 == total_offset[6:0] ? phv_data_89 : _GEN_88; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_90 = 7'h5a == total_offset[6:0] ? phv_data_90 : _GEN_89; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_91 = 7'h5b == total_offset[6:0] ? phv_data_91 : _GEN_90; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_92 = 7'h5c == total_offset[6:0] ? phv_data_92 : _GEN_91; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_93 = 7'h5d == total_offset[6:0] ? phv_data_93 : _GEN_92; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_94 = 7'h5e == total_offset[6:0] ? phv_data_94 : _GEN_93; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_95 = 7'h5f == total_offset[6:0] ? phv_data_95 : _GEN_94; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__0 = 8'h0 < length_0 ? _GEN_95 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_1 = offset_0 + 8'h1; // @[executor.scala 148:53]
  wire [7:0] _GEN_98 = 7'h1 == total_offset_1[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_99 = 7'h2 == total_offset_1[6:0] ? phv_data_2 : _GEN_98; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_100 = 7'h3 == total_offset_1[6:0] ? phv_data_3 : _GEN_99; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_101 = 7'h4 == total_offset_1[6:0] ? phv_data_4 : _GEN_100; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_102 = 7'h5 == total_offset_1[6:0] ? phv_data_5 : _GEN_101; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_103 = 7'h6 == total_offset_1[6:0] ? phv_data_6 : _GEN_102; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_104 = 7'h7 == total_offset_1[6:0] ? phv_data_7 : _GEN_103; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_105 = 7'h8 == total_offset_1[6:0] ? phv_data_8 : _GEN_104; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_106 = 7'h9 == total_offset_1[6:0] ? phv_data_9 : _GEN_105; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_107 = 7'ha == total_offset_1[6:0] ? phv_data_10 : _GEN_106; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_108 = 7'hb == total_offset_1[6:0] ? phv_data_11 : _GEN_107; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_109 = 7'hc == total_offset_1[6:0] ? phv_data_12 : _GEN_108; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_110 = 7'hd == total_offset_1[6:0] ? phv_data_13 : _GEN_109; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_111 = 7'he == total_offset_1[6:0] ? phv_data_14 : _GEN_110; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_112 = 7'hf == total_offset_1[6:0] ? phv_data_15 : _GEN_111; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_113 = 7'h10 == total_offset_1[6:0] ? phv_data_16 : _GEN_112; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_114 = 7'h11 == total_offset_1[6:0] ? phv_data_17 : _GEN_113; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_115 = 7'h12 == total_offset_1[6:0] ? phv_data_18 : _GEN_114; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_116 = 7'h13 == total_offset_1[6:0] ? phv_data_19 : _GEN_115; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_117 = 7'h14 == total_offset_1[6:0] ? phv_data_20 : _GEN_116; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_118 = 7'h15 == total_offset_1[6:0] ? phv_data_21 : _GEN_117; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_119 = 7'h16 == total_offset_1[6:0] ? phv_data_22 : _GEN_118; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_120 = 7'h17 == total_offset_1[6:0] ? phv_data_23 : _GEN_119; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_121 = 7'h18 == total_offset_1[6:0] ? phv_data_24 : _GEN_120; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_122 = 7'h19 == total_offset_1[6:0] ? phv_data_25 : _GEN_121; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_123 = 7'h1a == total_offset_1[6:0] ? phv_data_26 : _GEN_122; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_124 = 7'h1b == total_offset_1[6:0] ? phv_data_27 : _GEN_123; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_125 = 7'h1c == total_offset_1[6:0] ? phv_data_28 : _GEN_124; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_126 = 7'h1d == total_offset_1[6:0] ? phv_data_29 : _GEN_125; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_127 = 7'h1e == total_offset_1[6:0] ? phv_data_30 : _GEN_126; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_128 = 7'h1f == total_offset_1[6:0] ? phv_data_31 : _GEN_127; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_129 = 7'h20 == total_offset_1[6:0] ? phv_data_32 : _GEN_128; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_130 = 7'h21 == total_offset_1[6:0] ? phv_data_33 : _GEN_129; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_131 = 7'h22 == total_offset_1[6:0] ? phv_data_34 : _GEN_130; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_132 = 7'h23 == total_offset_1[6:0] ? phv_data_35 : _GEN_131; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_133 = 7'h24 == total_offset_1[6:0] ? phv_data_36 : _GEN_132; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_134 = 7'h25 == total_offset_1[6:0] ? phv_data_37 : _GEN_133; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_135 = 7'h26 == total_offset_1[6:0] ? phv_data_38 : _GEN_134; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_136 = 7'h27 == total_offset_1[6:0] ? phv_data_39 : _GEN_135; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_137 = 7'h28 == total_offset_1[6:0] ? phv_data_40 : _GEN_136; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_138 = 7'h29 == total_offset_1[6:0] ? phv_data_41 : _GEN_137; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_139 = 7'h2a == total_offset_1[6:0] ? phv_data_42 : _GEN_138; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_140 = 7'h2b == total_offset_1[6:0] ? phv_data_43 : _GEN_139; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_141 = 7'h2c == total_offset_1[6:0] ? phv_data_44 : _GEN_140; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_142 = 7'h2d == total_offset_1[6:0] ? phv_data_45 : _GEN_141; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_143 = 7'h2e == total_offset_1[6:0] ? phv_data_46 : _GEN_142; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_144 = 7'h2f == total_offset_1[6:0] ? phv_data_47 : _GEN_143; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_145 = 7'h30 == total_offset_1[6:0] ? phv_data_48 : _GEN_144; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_146 = 7'h31 == total_offset_1[6:0] ? phv_data_49 : _GEN_145; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_147 = 7'h32 == total_offset_1[6:0] ? phv_data_50 : _GEN_146; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_148 = 7'h33 == total_offset_1[6:0] ? phv_data_51 : _GEN_147; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_149 = 7'h34 == total_offset_1[6:0] ? phv_data_52 : _GEN_148; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_150 = 7'h35 == total_offset_1[6:0] ? phv_data_53 : _GEN_149; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_151 = 7'h36 == total_offset_1[6:0] ? phv_data_54 : _GEN_150; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_152 = 7'h37 == total_offset_1[6:0] ? phv_data_55 : _GEN_151; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_153 = 7'h38 == total_offset_1[6:0] ? phv_data_56 : _GEN_152; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_154 = 7'h39 == total_offset_1[6:0] ? phv_data_57 : _GEN_153; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_155 = 7'h3a == total_offset_1[6:0] ? phv_data_58 : _GEN_154; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_156 = 7'h3b == total_offset_1[6:0] ? phv_data_59 : _GEN_155; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_157 = 7'h3c == total_offset_1[6:0] ? phv_data_60 : _GEN_156; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_158 = 7'h3d == total_offset_1[6:0] ? phv_data_61 : _GEN_157; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_159 = 7'h3e == total_offset_1[6:0] ? phv_data_62 : _GEN_158; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_160 = 7'h3f == total_offset_1[6:0] ? phv_data_63 : _GEN_159; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_161 = 7'h40 == total_offset_1[6:0] ? phv_data_64 : _GEN_160; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_162 = 7'h41 == total_offset_1[6:0] ? phv_data_65 : _GEN_161; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_163 = 7'h42 == total_offset_1[6:0] ? phv_data_66 : _GEN_162; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_164 = 7'h43 == total_offset_1[6:0] ? phv_data_67 : _GEN_163; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_165 = 7'h44 == total_offset_1[6:0] ? phv_data_68 : _GEN_164; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_166 = 7'h45 == total_offset_1[6:0] ? phv_data_69 : _GEN_165; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_167 = 7'h46 == total_offset_1[6:0] ? phv_data_70 : _GEN_166; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_168 = 7'h47 == total_offset_1[6:0] ? phv_data_71 : _GEN_167; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_169 = 7'h48 == total_offset_1[6:0] ? phv_data_72 : _GEN_168; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_170 = 7'h49 == total_offset_1[6:0] ? phv_data_73 : _GEN_169; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_171 = 7'h4a == total_offset_1[6:0] ? phv_data_74 : _GEN_170; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_172 = 7'h4b == total_offset_1[6:0] ? phv_data_75 : _GEN_171; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_173 = 7'h4c == total_offset_1[6:0] ? phv_data_76 : _GEN_172; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_174 = 7'h4d == total_offset_1[6:0] ? phv_data_77 : _GEN_173; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_175 = 7'h4e == total_offset_1[6:0] ? phv_data_78 : _GEN_174; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_176 = 7'h4f == total_offset_1[6:0] ? phv_data_79 : _GEN_175; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_177 = 7'h50 == total_offset_1[6:0] ? phv_data_80 : _GEN_176; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_178 = 7'h51 == total_offset_1[6:0] ? phv_data_81 : _GEN_177; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_179 = 7'h52 == total_offset_1[6:0] ? phv_data_82 : _GEN_178; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_180 = 7'h53 == total_offset_1[6:0] ? phv_data_83 : _GEN_179; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_181 = 7'h54 == total_offset_1[6:0] ? phv_data_84 : _GEN_180; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_182 = 7'h55 == total_offset_1[6:0] ? phv_data_85 : _GEN_181; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_183 = 7'h56 == total_offset_1[6:0] ? phv_data_86 : _GEN_182; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_184 = 7'h57 == total_offset_1[6:0] ? phv_data_87 : _GEN_183; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_185 = 7'h58 == total_offset_1[6:0] ? phv_data_88 : _GEN_184; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_186 = 7'h59 == total_offset_1[6:0] ? phv_data_89 : _GEN_185; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_187 = 7'h5a == total_offset_1[6:0] ? phv_data_90 : _GEN_186; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_188 = 7'h5b == total_offset_1[6:0] ? phv_data_91 : _GEN_187; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_189 = 7'h5c == total_offset_1[6:0] ? phv_data_92 : _GEN_188; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_190 = 7'h5d == total_offset_1[6:0] ? phv_data_93 : _GEN_189; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_191 = 7'h5e == total_offset_1[6:0] ? phv_data_94 : _GEN_190; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_192 = 7'h5f == total_offset_1[6:0] ? phv_data_95 : _GEN_191; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__1 = 8'h1 < length_0 ? _GEN_192 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_2 = offset_0 + 8'h2; // @[executor.scala 148:53]
  wire [7:0] _GEN_195 = 7'h1 == total_offset_2[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_196 = 7'h2 == total_offset_2[6:0] ? phv_data_2 : _GEN_195; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_197 = 7'h3 == total_offset_2[6:0] ? phv_data_3 : _GEN_196; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_198 = 7'h4 == total_offset_2[6:0] ? phv_data_4 : _GEN_197; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_199 = 7'h5 == total_offset_2[6:0] ? phv_data_5 : _GEN_198; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_200 = 7'h6 == total_offset_2[6:0] ? phv_data_6 : _GEN_199; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_201 = 7'h7 == total_offset_2[6:0] ? phv_data_7 : _GEN_200; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_202 = 7'h8 == total_offset_2[6:0] ? phv_data_8 : _GEN_201; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_203 = 7'h9 == total_offset_2[6:0] ? phv_data_9 : _GEN_202; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_204 = 7'ha == total_offset_2[6:0] ? phv_data_10 : _GEN_203; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_205 = 7'hb == total_offset_2[6:0] ? phv_data_11 : _GEN_204; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_206 = 7'hc == total_offset_2[6:0] ? phv_data_12 : _GEN_205; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_207 = 7'hd == total_offset_2[6:0] ? phv_data_13 : _GEN_206; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_208 = 7'he == total_offset_2[6:0] ? phv_data_14 : _GEN_207; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_209 = 7'hf == total_offset_2[6:0] ? phv_data_15 : _GEN_208; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_210 = 7'h10 == total_offset_2[6:0] ? phv_data_16 : _GEN_209; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_211 = 7'h11 == total_offset_2[6:0] ? phv_data_17 : _GEN_210; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_212 = 7'h12 == total_offset_2[6:0] ? phv_data_18 : _GEN_211; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_213 = 7'h13 == total_offset_2[6:0] ? phv_data_19 : _GEN_212; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_214 = 7'h14 == total_offset_2[6:0] ? phv_data_20 : _GEN_213; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_215 = 7'h15 == total_offset_2[6:0] ? phv_data_21 : _GEN_214; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_216 = 7'h16 == total_offset_2[6:0] ? phv_data_22 : _GEN_215; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_217 = 7'h17 == total_offset_2[6:0] ? phv_data_23 : _GEN_216; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_218 = 7'h18 == total_offset_2[6:0] ? phv_data_24 : _GEN_217; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_219 = 7'h19 == total_offset_2[6:0] ? phv_data_25 : _GEN_218; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_220 = 7'h1a == total_offset_2[6:0] ? phv_data_26 : _GEN_219; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_221 = 7'h1b == total_offset_2[6:0] ? phv_data_27 : _GEN_220; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_222 = 7'h1c == total_offset_2[6:0] ? phv_data_28 : _GEN_221; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_223 = 7'h1d == total_offset_2[6:0] ? phv_data_29 : _GEN_222; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_224 = 7'h1e == total_offset_2[6:0] ? phv_data_30 : _GEN_223; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_225 = 7'h1f == total_offset_2[6:0] ? phv_data_31 : _GEN_224; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_226 = 7'h20 == total_offset_2[6:0] ? phv_data_32 : _GEN_225; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_227 = 7'h21 == total_offset_2[6:0] ? phv_data_33 : _GEN_226; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_228 = 7'h22 == total_offset_2[6:0] ? phv_data_34 : _GEN_227; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_229 = 7'h23 == total_offset_2[6:0] ? phv_data_35 : _GEN_228; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_230 = 7'h24 == total_offset_2[6:0] ? phv_data_36 : _GEN_229; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_231 = 7'h25 == total_offset_2[6:0] ? phv_data_37 : _GEN_230; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_232 = 7'h26 == total_offset_2[6:0] ? phv_data_38 : _GEN_231; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_233 = 7'h27 == total_offset_2[6:0] ? phv_data_39 : _GEN_232; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_234 = 7'h28 == total_offset_2[6:0] ? phv_data_40 : _GEN_233; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_235 = 7'h29 == total_offset_2[6:0] ? phv_data_41 : _GEN_234; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_236 = 7'h2a == total_offset_2[6:0] ? phv_data_42 : _GEN_235; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_237 = 7'h2b == total_offset_2[6:0] ? phv_data_43 : _GEN_236; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_238 = 7'h2c == total_offset_2[6:0] ? phv_data_44 : _GEN_237; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_239 = 7'h2d == total_offset_2[6:0] ? phv_data_45 : _GEN_238; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_240 = 7'h2e == total_offset_2[6:0] ? phv_data_46 : _GEN_239; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_241 = 7'h2f == total_offset_2[6:0] ? phv_data_47 : _GEN_240; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_242 = 7'h30 == total_offset_2[6:0] ? phv_data_48 : _GEN_241; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_243 = 7'h31 == total_offset_2[6:0] ? phv_data_49 : _GEN_242; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_244 = 7'h32 == total_offset_2[6:0] ? phv_data_50 : _GEN_243; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_245 = 7'h33 == total_offset_2[6:0] ? phv_data_51 : _GEN_244; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_246 = 7'h34 == total_offset_2[6:0] ? phv_data_52 : _GEN_245; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_247 = 7'h35 == total_offset_2[6:0] ? phv_data_53 : _GEN_246; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_248 = 7'h36 == total_offset_2[6:0] ? phv_data_54 : _GEN_247; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_249 = 7'h37 == total_offset_2[6:0] ? phv_data_55 : _GEN_248; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_250 = 7'h38 == total_offset_2[6:0] ? phv_data_56 : _GEN_249; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_251 = 7'h39 == total_offset_2[6:0] ? phv_data_57 : _GEN_250; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_252 = 7'h3a == total_offset_2[6:0] ? phv_data_58 : _GEN_251; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_253 = 7'h3b == total_offset_2[6:0] ? phv_data_59 : _GEN_252; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_254 = 7'h3c == total_offset_2[6:0] ? phv_data_60 : _GEN_253; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_255 = 7'h3d == total_offset_2[6:0] ? phv_data_61 : _GEN_254; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_256 = 7'h3e == total_offset_2[6:0] ? phv_data_62 : _GEN_255; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_257 = 7'h3f == total_offset_2[6:0] ? phv_data_63 : _GEN_256; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_258 = 7'h40 == total_offset_2[6:0] ? phv_data_64 : _GEN_257; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_259 = 7'h41 == total_offset_2[6:0] ? phv_data_65 : _GEN_258; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_260 = 7'h42 == total_offset_2[6:0] ? phv_data_66 : _GEN_259; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_261 = 7'h43 == total_offset_2[6:0] ? phv_data_67 : _GEN_260; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_262 = 7'h44 == total_offset_2[6:0] ? phv_data_68 : _GEN_261; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_263 = 7'h45 == total_offset_2[6:0] ? phv_data_69 : _GEN_262; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_264 = 7'h46 == total_offset_2[6:0] ? phv_data_70 : _GEN_263; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_265 = 7'h47 == total_offset_2[6:0] ? phv_data_71 : _GEN_264; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_266 = 7'h48 == total_offset_2[6:0] ? phv_data_72 : _GEN_265; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_267 = 7'h49 == total_offset_2[6:0] ? phv_data_73 : _GEN_266; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_268 = 7'h4a == total_offset_2[6:0] ? phv_data_74 : _GEN_267; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_269 = 7'h4b == total_offset_2[6:0] ? phv_data_75 : _GEN_268; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_270 = 7'h4c == total_offset_2[6:0] ? phv_data_76 : _GEN_269; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_271 = 7'h4d == total_offset_2[6:0] ? phv_data_77 : _GEN_270; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_272 = 7'h4e == total_offset_2[6:0] ? phv_data_78 : _GEN_271; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_273 = 7'h4f == total_offset_2[6:0] ? phv_data_79 : _GEN_272; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_274 = 7'h50 == total_offset_2[6:0] ? phv_data_80 : _GEN_273; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_275 = 7'h51 == total_offset_2[6:0] ? phv_data_81 : _GEN_274; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_276 = 7'h52 == total_offset_2[6:0] ? phv_data_82 : _GEN_275; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_277 = 7'h53 == total_offset_2[6:0] ? phv_data_83 : _GEN_276; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_278 = 7'h54 == total_offset_2[6:0] ? phv_data_84 : _GEN_277; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_279 = 7'h55 == total_offset_2[6:0] ? phv_data_85 : _GEN_278; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_280 = 7'h56 == total_offset_2[6:0] ? phv_data_86 : _GEN_279; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_281 = 7'h57 == total_offset_2[6:0] ? phv_data_87 : _GEN_280; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_282 = 7'h58 == total_offset_2[6:0] ? phv_data_88 : _GEN_281; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_283 = 7'h59 == total_offset_2[6:0] ? phv_data_89 : _GEN_282; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_284 = 7'h5a == total_offset_2[6:0] ? phv_data_90 : _GEN_283; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_285 = 7'h5b == total_offset_2[6:0] ? phv_data_91 : _GEN_284; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_286 = 7'h5c == total_offset_2[6:0] ? phv_data_92 : _GEN_285; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_287 = 7'h5d == total_offset_2[6:0] ? phv_data_93 : _GEN_286; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_288 = 7'h5e == total_offset_2[6:0] ? phv_data_94 : _GEN_287; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_289 = 7'h5f == total_offset_2[6:0] ? phv_data_95 : _GEN_288; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__2 = 8'h2 < length_0 ? _GEN_289 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_3 = offset_0 + 8'h3; // @[executor.scala 148:53]
  wire [7:0] _GEN_292 = 7'h1 == total_offset_3[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_293 = 7'h2 == total_offset_3[6:0] ? phv_data_2 : _GEN_292; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_294 = 7'h3 == total_offset_3[6:0] ? phv_data_3 : _GEN_293; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_295 = 7'h4 == total_offset_3[6:0] ? phv_data_4 : _GEN_294; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_296 = 7'h5 == total_offset_3[6:0] ? phv_data_5 : _GEN_295; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_297 = 7'h6 == total_offset_3[6:0] ? phv_data_6 : _GEN_296; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_298 = 7'h7 == total_offset_3[6:0] ? phv_data_7 : _GEN_297; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_299 = 7'h8 == total_offset_3[6:0] ? phv_data_8 : _GEN_298; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_300 = 7'h9 == total_offset_3[6:0] ? phv_data_9 : _GEN_299; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_301 = 7'ha == total_offset_3[6:0] ? phv_data_10 : _GEN_300; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_302 = 7'hb == total_offset_3[6:0] ? phv_data_11 : _GEN_301; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_303 = 7'hc == total_offset_3[6:0] ? phv_data_12 : _GEN_302; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_304 = 7'hd == total_offset_3[6:0] ? phv_data_13 : _GEN_303; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_305 = 7'he == total_offset_3[6:0] ? phv_data_14 : _GEN_304; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_306 = 7'hf == total_offset_3[6:0] ? phv_data_15 : _GEN_305; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_307 = 7'h10 == total_offset_3[6:0] ? phv_data_16 : _GEN_306; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_308 = 7'h11 == total_offset_3[6:0] ? phv_data_17 : _GEN_307; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_309 = 7'h12 == total_offset_3[6:0] ? phv_data_18 : _GEN_308; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_310 = 7'h13 == total_offset_3[6:0] ? phv_data_19 : _GEN_309; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_311 = 7'h14 == total_offset_3[6:0] ? phv_data_20 : _GEN_310; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_312 = 7'h15 == total_offset_3[6:0] ? phv_data_21 : _GEN_311; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_313 = 7'h16 == total_offset_3[6:0] ? phv_data_22 : _GEN_312; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_314 = 7'h17 == total_offset_3[6:0] ? phv_data_23 : _GEN_313; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_315 = 7'h18 == total_offset_3[6:0] ? phv_data_24 : _GEN_314; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_316 = 7'h19 == total_offset_3[6:0] ? phv_data_25 : _GEN_315; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_317 = 7'h1a == total_offset_3[6:0] ? phv_data_26 : _GEN_316; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_318 = 7'h1b == total_offset_3[6:0] ? phv_data_27 : _GEN_317; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_319 = 7'h1c == total_offset_3[6:0] ? phv_data_28 : _GEN_318; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_320 = 7'h1d == total_offset_3[6:0] ? phv_data_29 : _GEN_319; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_321 = 7'h1e == total_offset_3[6:0] ? phv_data_30 : _GEN_320; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_322 = 7'h1f == total_offset_3[6:0] ? phv_data_31 : _GEN_321; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_323 = 7'h20 == total_offset_3[6:0] ? phv_data_32 : _GEN_322; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_324 = 7'h21 == total_offset_3[6:0] ? phv_data_33 : _GEN_323; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_325 = 7'h22 == total_offset_3[6:0] ? phv_data_34 : _GEN_324; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_326 = 7'h23 == total_offset_3[6:0] ? phv_data_35 : _GEN_325; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_327 = 7'h24 == total_offset_3[6:0] ? phv_data_36 : _GEN_326; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_328 = 7'h25 == total_offset_3[6:0] ? phv_data_37 : _GEN_327; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_329 = 7'h26 == total_offset_3[6:0] ? phv_data_38 : _GEN_328; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_330 = 7'h27 == total_offset_3[6:0] ? phv_data_39 : _GEN_329; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_331 = 7'h28 == total_offset_3[6:0] ? phv_data_40 : _GEN_330; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_332 = 7'h29 == total_offset_3[6:0] ? phv_data_41 : _GEN_331; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_333 = 7'h2a == total_offset_3[6:0] ? phv_data_42 : _GEN_332; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_334 = 7'h2b == total_offset_3[6:0] ? phv_data_43 : _GEN_333; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_335 = 7'h2c == total_offset_3[6:0] ? phv_data_44 : _GEN_334; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_336 = 7'h2d == total_offset_3[6:0] ? phv_data_45 : _GEN_335; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_337 = 7'h2e == total_offset_3[6:0] ? phv_data_46 : _GEN_336; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_338 = 7'h2f == total_offset_3[6:0] ? phv_data_47 : _GEN_337; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_339 = 7'h30 == total_offset_3[6:0] ? phv_data_48 : _GEN_338; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_340 = 7'h31 == total_offset_3[6:0] ? phv_data_49 : _GEN_339; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_341 = 7'h32 == total_offset_3[6:0] ? phv_data_50 : _GEN_340; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_342 = 7'h33 == total_offset_3[6:0] ? phv_data_51 : _GEN_341; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_343 = 7'h34 == total_offset_3[6:0] ? phv_data_52 : _GEN_342; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_344 = 7'h35 == total_offset_3[6:0] ? phv_data_53 : _GEN_343; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_345 = 7'h36 == total_offset_3[6:0] ? phv_data_54 : _GEN_344; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_346 = 7'h37 == total_offset_3[6:0] ? phv_data_55 : _GEN_345; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_347 = 7'h38 == total_offset_3[6:0] ? phv_data_56 : _GEN_346; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_348 = 7'h39 == total_offset_3[6:0] ? phv_data_57 : _GEN_347; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_349 = 7'h3a == total_offset_3[6:0] ? phv_data_58 : _GEN_348; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_350 = 7'h3b == total_offset_3[6:0] ? phv_data_59 : _GEN_349; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_351 = 7'h3c == total_offset_3[6:0] ? phv_data_60 : _GEN_350; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_352 = 7'h3d == total_offset_3[6:0] ? phv_data_61 : _GEN_351; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_353 = 7'h3e == total_offset_3[6:0] ? phv_data_62 : _GEN_352; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_354 = 7'h3f == total_offset_3[6:0] ? phv_data_63 : _GEN_353; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_355 = 7'h40 == total_offset_3[6:0] ? phv_data_64 : _GEN_354; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_356 = 7'h41 == total_offset_3[6:0] ? phv_data_65 : _GEN_355; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_357 = 7'h42 == total_offset_3[6:0] ? phv_data_66 : _GEN_356; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_358 = 7'h43 == total_offset_3[6:0] ? phv_data_67 : _GEN_357; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_359 = 7'h44 == total_offset_3[6:0] ? phv_data_68 : _GEN_358; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_360 = 7'h45 == total_offset_3[6:0] ? phv_data_69 : _GEN_359; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_361 = 7'h46 == total_offset_3[6:0] ? phv_data_70 : _GEN_360; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_362 = 7'h47 == total_offset_3[6:0] ? phv_data_71 : _GEN_361; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_363 = 7'h48 == total_offset_3[6:0] ? phv_data_72 : _GEN_362; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_364 = 7'h49 == total_offset_3[6:0] ? phv_data_73 : _GEN_363; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_365 = 7'h4a == total_offset_3[6:0] ? phv_data_74 : _GEN_364; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_366 = 7'h4b == total_offset_3[6:0] ? phv_data_75 : _GEN_365; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_367 = 7'h4c == total_offset_3[6:0] ? phv_data_76 : _GEN_366; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_368 = 7'h4d == total_offset_3[6:0] ? phv_data_77 : _GEN_367; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_369 = 7'h4e == total_offset_3[6:0] ? phv_data_78 : _GEN_368; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_370 = 7'h4f == total_offset_3[6:0] ? phv_data_79 : _GEN_369; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_371 = 7'h50 == total_offset_3[6:0] ? phv_data_80 : _GEN_370; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_372 = 7'h51 == total_offset_3[6:0] ? phv_data_81 : _GEN_371; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_373 = 7'h52 == total_offset_3[6:0] ? phv_data_82 : _GEN_372; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_374 = 7'h53 == total_offset_3[6:0] ? phv_data_83 : _GEN_373; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_375 = 7'h54 == total_offset_3[6:0] ? phv_data_84 : _GEN_374; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_376 = 7'h55 == total_offset_3[6:0] ? phv_data_85 : _GEN_375; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_377 = 7'h56 == total_offset_3[6:0] ? phv_data_86 : _GEN_376; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_378 = 7'h57 == total_offset_3[6:0] ? phv_data_87 : _GEN_377; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_379 = 7'h58 == total_offset_3[6:0] ? phv_data_88 : _GEN_378; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_380 = 7'h59 == total_offset_3[6:0] ? phv_data_89 : _GEN_379; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_381 = 7'h5a == total_offset_3[6:0] ? phv_data_90 : _GEN_380; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_382 = 7'h5b == total_offset_3[6:0] ? phv_data_91 : _GEN_381; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_383 = 7'h5c == total_offset_3[6:0] ? phv_data_92 : _GEN_382; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_384 = 7'h5d == total_offset_3[6:0] ? phv_data_93 : _GEN_383; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_385 = 7'h5e == total_offset_3[6:0] ? phv_data_94 : _GEN_384; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_386 = 7'h5f == total_offset_3[6:0] ? phv_data_95 : _GEN_385; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__3 = 8'h3 < length_0 ? _GEN_386 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_4 = offset_0 + 8'h4; // @[executor.scala 148:53]
  wire [7:0] _GEN_389 = 7'h1 == total_offset_4[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_390 = 7'h2 == total_offset_4[6:0] ? phv_data_2 : _GEN_389; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_391 = 7'h3 == total_offset_4[6:0] ? phv_data_3 : _GEN_390; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_392 = 7'h4 == total_offset_4[6:0] ? phv_data_4 : _GEN_391; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_393 = 7'h5 == total_offset_4[6:0] ? phv_data_5 : _GEN_392; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_394 = 7'h6 == total_offset_4[6:0] ? phv_data_6 : _GEN_393; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_395 = 7'h7 == total_offset_4[6:0] ? phv_data_7 : _GEN_394; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_396 = 7'h8 == total_offset_4[6:0] ? phv_data_8 : _GEN_395; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_397 = 7'h9 == total_offset_4[6:0] ? phv_data_9 : _GEN_396; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_398 = 7'ha == total_offset_4[6:0] ? phv_data_10 : _GEN_397; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_399 = 7'hb == total_offset_4[6:0] ? phv_data_11 : _GEN_398; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_400 = 7'hc == total_offset_4[6:0] ? phv_data_12 : _GEN_399; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_401 = 7'hd == total_offset_4[6:0] ? phv_data_13 : _GEN_400; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_402 = 7'he == total_offset_4[6:0] ? phv_data_14 : _GEN_401; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_403 = 7'hf == total_offset_4[6:0] ? phv_data_15 : _GEN_402; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_404 = 7'h10 == total_offset_4[6:0] ? phv_data_16 : _GEN_403; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_405 = 7'h11 == total_offset_4[6:0] ? phv_data_17 : _GEN_404; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_406 = 7'h12 == total_offset_4[6:0] ? phv_data_18 : _GEN_405; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_407 = 7'h13 == total_offset_4[6:0] ? phv_data_19 : _GEN_406; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_408 = 7'h14 == total_offset_4[6:0] ? phv_data_20 : _GEN_407; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_409 = 7'h15 == total_offset_4[6:0] ? phv_data_21 : _GEN_408; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_410 = 7'h16 == total_offset_4[6:0] ? phv_data_22 : _GEN_409; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_411 = 7'h17 == total_offset_4[6:0] ? phv_data_23 : _GEN_410; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_412 = 7'h18 == total_offset_4[6:0] ? phv_data_24 : _GEN_411; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_413 = 7'h19 == total_offset_4[6:0] ? phv_data_25 : _GEN_412; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_414 = 7'h1a == total_offset_4[6:0] ? phv_data_26 : _GEN_413; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_415 = 7'h1b == total_offset_4[6:0] ? phv_data_27 : _GEN_414; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_416 = 7'h1c == total_offset_4[6:0] ? phv_data_28 : _GEN_415; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_417 = 7'h1d == total_offset_4[6:0] ? phv_data_29 : _GEN_416; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_418 = 7'h1e == total_offset_4[6:0] ? phv_data_30 : _GEN_417; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_419 = 7'h1f == total_offset_4[6:0] ? phv_data_31 : _GEN_418; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_420 = 7'h20 == total_offset_4[6:0] ? phv_data_32 : _GEN_419; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_421 = 7'h21 == total_offset_4[6:0] ? phv_data_33 : _GEN_420; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_422 = 7'h22 == total_offset_4[6:0] ? phv_data_34 : _GEN_421; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_423 = 7'h23 == total_offset_4[6:0] ? phv_data_35 : _GEN_422; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_424 = 7'h24 == total_offset_4[6:0] ? phv_data_36 : _GEN_423; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_425 = 7'h25 == total_offset_4[6:0] ? phv_data_37 : _GEN_424; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_426 = 7'h26 == total_offset_4[6:0] ? phv_data_38 : _GEN_425; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_427 = 7'h27 == total_offset_4[6:0] ? phv_data_39 : _GEN_426; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_428 = 7'h28 == total_offset_4[6:0] ? phv_data_40 : _GEN_427; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_429 = 7'h29 == total_offset_4[6:0] ? phv_data_41 : _GEN_428; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_430 = 7'h2a == total_offset_4[6:0] ? phv_data_42 : _GEN_429; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_431 = 7'h2b == total_offset_4[6:0] ? phv_data_43 : _GEN_430; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_432 = 7'h2c == total_offset_4[6:0] ? phv_data_44 : _GEN_431; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_433 = 7'h2d == total_offset_4[6:0] ? phv_data_45 : _GEN_432; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_434 = 7'h2e == total_offset_4[6:0] ? phv_data_46 : _GEN_433; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_435 = 7'h2f == total_offset_4[6:0] ? phv_data_47 : _GEN_434; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_436 = 7'h30 == total_offset_4[6:0] ? phv_data_48 : _GEN_435; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_437 = 7'h31 == total_offset_4[6:0] ? phv_data_49 : _GEN_436; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_438 = 7'h32 == total_offset_4[6:0] ? phv_data_50 : _GEN_437; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_439 = 7'h33 == total_offset_4[6:0] ? phv_data_51 : _GEN_438; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_440 = 7'h34 == total_offset_4[6:0] ? phv_data_52 : _GEN_439; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_441 = 7'h35 == total_offset_4[6:0] ? phv_data_53 : _GEN_440; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_442 = 7'h36 == total_offset_4[6:0] ? phv_data_54 : _GEN_441; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_443 = 7'h37 == total_offset_4[6:0] ? phv_data_55 : _GEN_442; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_444 = 7'h38 == total_offset_4[6:0] ? phv_data_56 : _GEN_443; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_445 = 7'h39 == total_offset_4[6:0] ? phv_data_57 : _GEN_444; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_446 = 7'h3a == total_offset_4[6:0] ? phv_data_58 : _GEN_445; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_447 = 7'h3b == total_offset_4[6:0] ? phv_data_59 : _GEN_446; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_448 = 7'h3c == total_offset_4[6:0] ? phv_data_60 : _GEN_447; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_449 = 7'h3d == total_offset_4[6:0] ? phv_data_61 : _GEN_448; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_450 = 7'h3e == total_offset_4[6:0] ? phv_data_62 : _GEN_449; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_451 = 7'h3f == total_offset_4[6:0] ? phv_data_63 : _GEN_450; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_452 = 7'h40 == total_offset_4[6:0] ? phv_data_64 : _GEN_451; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_453 = 7'h41 == total_offset_4[6:0] ? phv_data_65 : _GEN_452; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_454 = 7'h42 == total_offset_4[6:0] ? phv_data_66 : _GEN_453; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_455 = 7'h43 == total_offset_4[6:0] ? phv_data_67 : _GEN_454; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_456 = 7'h44 == total_offset_4[6:0] ? phv_data_68 : _GEN_455; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_457 = 7'h45 == total_offset_4[6:0] ? phv_data_69 : _GEN_456; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_458 = 7'h46 == total_offset_4[6:0] ? phv_data_70 : _GEN_457; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_459 = 7'h47 == total_offset_4[6:0] ? phv_data_71 : _GEN_458; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_460 = 7'h48 == total_offset_4[6:0] ? phv_data_72 : _GEN_459; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_461 = 7'h49 == total_offset_4[6:0] ? phv_data_73 : _GEN_460; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_462 = 7'h4a == total_offset_4[6:0] ? phv_data_74 : _GEN_461; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_463 = 7'h4b == total_offset_4[6:0] ? phv_data_75 : _GEN_462; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_464 = 7'h4c == total_offset_4[6:0] ? phv_data_76 : _GEN_463; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_465 = 7'h4d == total_offset_4[6:0] ? phv_data_77 : _GEN_464; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_466 = 7'h4e == total_offset_4[6:0] ? phv_data_78 : _GEN_465; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_467 = 7'h4f == total_offset_4[6:0] ? phv_data_79 : _GEN_466; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_468 = 7'h50 == total_offset_4[6:0] ? phv_data_80 : _GEN_467; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_469 = 7'h51 == total_offset_4[6:0] ? phv_data_81 : _GEN_468; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_470 = 7'h52 == total_offset_4[6:0] ? phv_data_82 : _GEN_469; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_471 = 7'h53 == total_offset_4[6:0] ? phv_data_83 : _GEN_470; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_472 = 7'h54 == total_offset_4[6:0] ? phv_data_84 : _GEN_471; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_473 = 7'h55 == total_offset_4[6:0] ? phv_data_85 : _GEN_472; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_474 = 7'h56 == total_offset_4[6:0] ? phv_data_86 : _GEN_473; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_475 = 7'h57 == total_offset_4[6:0] ? phv_data_87 : _GEN_474; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_476 = 7'h58 == total_offset_4[6:0] ? phv_data_88 : _GEN_475; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_477 = 7'h59 == total_offset_4[6:0] ? phv_data_89 : _GEN_476; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_478 = 7'h5a == total_offset_4[6:0] ? phv_data_90 : _GEN_477; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_479 = 7'h5b == total_offset_4[6:0] ? phv_data_91 : _GEN_478; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_480 = 7'h5c == total_offset_4[6:0] ? phv_data_92 : _GEN_479; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_481 = 7'h5d == total_offset_4[6:0] ? phv_data_93 : _GEN_480; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_482 = 7'h5e == total_offset_4[6:0] ? phv_data_94 : _GEN_481; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_483 = 7'h5f == total_offset_4[6:0] ? phv_data_95 : _GEN_482; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__4 = 8'h4 < length_0 ? _GEN_483 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_5 = offset_0 + 8'h5; // @[executor.scala 148:53]
  wire [7:0] _GEN_486 = 7'h1 == total_offset_5[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_487 = 7'h2 == total_offset_5[6:0] ? phv_data_2 : _GEN_486; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_488 = 7'h3 == total_offset_5[6:0] ? phv_data_3 : _GEN_487; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_489 = 7'h4 == total_offset_5[6:0] ? phv_data_4 : _GEN_488; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_490 = 7'h5 == total_offset_5[6:0] ? phv_data_5 : _GEN_489; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_491 = 7'h6 == total_offset_5[6:0] ? phv_data_6 : _GEN_490; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_492 = 7'h7 == total_offset_5[6:0] ? phv_data_7 : _GEN_491; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_493 = 7'h8 == total_offset_5[6:0] ? phv_data_8 : _GEN_492; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_494 = 7'h9 == total_offset_5[6:0] ? phv_data_9 : _GEN_493; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_495 = 7'ha == total_offset_5[6:0] ? phv_data_10 : _GEN_494; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_496 = 7'hb == total_offset_5[6:0] ? phv_data_11 : _GEN_495; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_497 = 7'hc == total_offset_5[6:0] ? phv_data_12 : _GEN_496; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_498 = 7'hd == total_offset_5[6:0] ? phv_data_13 : _GEN_497; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_499 = 7'he == total_offset_5[6:0] ? phv_data_14 : _GEN_498; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_500 = 7'hf == total_offset_5[6:0] ? phv_data_15 : _GEN_499; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_501 = 7'h10 == total_offset_5[6:0] ? phv_data_16 : _GEN_500; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_502 = 7'h11 == total_offset_5[6:0] ? phv_data_17 : _GEN_501; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_503 = 7'h12 == total_offset_5[6:0] ? phv_data_18 : _GEN_502; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_504 = 7'h13 == total_offset_5[6:0] ? phv_data_19 : _GEN_503; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_505 = 7'h14 == total_offset_5[6:0] ? phv_data_20 : _GEN_504; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_506 = 7'h15 == total_offset_5[6:0] ? phv_data_21 : _GEN_505; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_507 = 7'h16 == total_offset_5[6:0] ? phv_data_22 : _GEN_506; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_508 = 7'h17 == total_offset_5[6:0] ? phv_data_23 : _GEN_507; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_509 = 7'h18 == total_offset_5[6:0] ? phv_data_24 : _GEN_508; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_510 = 7'h19 == total_offset_5[6:0] ? phv_data_25 : _GEN_509; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_511 = 7'h1a == total_offset_5[6:0] ? phv_data_26 : _GEN_510; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_512 = 7'h1b == total_offset_5[6:0] ? phv_data_27 : _GEN_511; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_513 = 7'h1c == total_offset_5[6:0] ? phv_data_28 : _GEN_512; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_514 = 7'h1d == total_offset_5[6:0] ? phv_data_29 : _GEN_513; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_515 = 7'h1e == total_offset_5[6:0] ? phv_data_30 : _GEN_514; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_516 = 7'h1f == total_offset_5[6:0] ? phv_data_31 : _GEN_515; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_517 = 7'h20 == total_offset_5[6:0] ? phv_data_32 : _GEN_516; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_518 = 7'h21 == total_offset_5[6:0] ? phv_data_33 : _GEN_517; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_519 = 7'h22 == total_offset_5[6:0] ? phv_data_34 : _GEN_518; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_520 = 7'h23 == total_offset_5[6:0] ? phv_data_35 : _GEN_519; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_521 = 7'h24 == total_offset_5[6:0] ? phv_data_36 : _GEN_520; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_522 = 7'h25 == total_offset_5[6:0] ? phv_data_37 : _GEN_521; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_523 = 7'h26 == total_offset_5[6:0] ? phv_data_38 : _GEN_522; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_524 = 7'h27 == total_offset_5[6:0] ? phv_data_39 : _GEN_523; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_525 = 7'h28 == total_offset_5[6:0] ? phv_data_40 : _GEN_524; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_526 = 7'h29 == total_offset_5[6:0] ? phv_data_41 : _GEN_525; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_527 = 7'h2a == total_offset_5[6:0] ? phv_data_42 : _GEN_526; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_528 = 7'h2b == total_offset_5[6:0] ? phv_data_43 : _GEN_527; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_529 = 7'h2c == total_offset_5[6:0] ? phv_data_44 : _GEN_528; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_530 = 7'h2d == total_offset_5[6:0] ? phv_data_45 : _GEN_529; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_531 = 7'h2e == total_offset_5[6:0] ? phv_data_46 : _GEN_530; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_532 = 7'h2f == total_offset_5[6:0] ? phv_data_47 : _GEN_531; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_533 = 7'h30 == total_offset_5[6:0] ? phv_data_48 : _GEN_532; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_534 = 7'h31 == total_offset_5[6:0] ? phv_data_49 : _GEN_533; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_535 = 7'h32 == total_offset_5[6:0] ? phv_data_50 : _GEN_534; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_536 = 7'h33 == total_offset_5[6:0] ? phv_data_51 : _GEN_535; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_537 = 7'h34 == total_offset_5[6:0] ? phv_data_52 : _GEN_536; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_538 = 7'h35 == total_offset_5[6:0] ? phv_data_53 : _GEN_537; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_539 = 7'h36 == total_offset_5[6:0] ? phv_data_54 : _GEN_538; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_540 = 7'h37 == total_offset_5[6:0] ? phv_data_55 : _GEN_539; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_541 = 7'h38 == total_offset_5[6:0] ? phv_data_56 : _GEN_540; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_542 = 7'h39 == total_offset_5[6:0] ? phv_data_57 : _GEN_541; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_543 = 7'h3a == total_offset_5[6:0] ? phv_data_58 : _GEN_542; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_544 = 7'h3b == total_offset_5[6:0] ? phv_data_59 : _GEN_543; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_545 = 7'h3c == total_offset_5[6:0] ? phv_data_60 : _GEN_544; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_546 = 7'h3d == total_offset_5[6:0] ? phv_data_61 : _GEN_545; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_547 = 7'h3e == total_offset_5[6:0] ? phv_data_62 : _GEN_546; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_548 = 7'h3f == total_offset_5[6:0] ? phv_data_63 : _GEN_547; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_549 = 7'h40 == total_offset_5[6:0] ? phv_data_64 : _GEN_548; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_550 = 7'h41 == total_offset_5[6:0] ? phv_data_65 : _GEN_549; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_551 = 7'h42 == total_offset_5[6:0] ? phv_data_66 : _GEN_550; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_552 = 7'h43 == total_offset_5[6:0] ? phv_data_67 : _GEN_551; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_553 = 7'h44 == total_offset_5[6:0] ? phv_data_68 : _GEN_552; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_554 = 7'h45 == total_offset_5[6:0] ? phv_data_69 : _GEN_553; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_555 = 7'h46 == total_offset_5[6:0] ? phv_data_70 : _GEN_554; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_556 = 7'h47 == total_offset_5[6:0] ? phv_data_71 : _GEN_555; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_557 = 7'h48 == total_offset_5[6:0] ? phv_data_72 : _GEN_556; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_558 = 7'h49 == total_offset_5[6:0] ? phv_data_73 : _GEN_557; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_559 = 7'h4a == total_offset_5[6:0] ? phv_data_74 : _GEN_558; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_560 = 7'h4b == total_offset_5[6:0] ? phv_data_75 : _GEN_559; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_561 = 7'h4c == total_offset_5[6:0] ? phv_data_76 : _GEN_560; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_562 = 7'h4d == total_offset_5[6:0] ? phv_data_77 : _GEN_561; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_563 = 7'h4e == total_offset_5[6:0] ? phv_data_78 : _GEN_562; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_564 = 7'h4f == total_offset_5[6:0] ? phv_data_79 : _GEN_563; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_565 = 7'h50 == total_offset_5[6:0] ? phv_data_80 : _GEN_564; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_566 = 7'h51 == total_offset_5[6:0] ? phv_data_81 : _GEN_565; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_567 = 7'h52 == total_offset_5[6:0] ? phv_data_82 : _GEN_566; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_568 = 7'h53 == total_offset_5[6:0] ? phv_data_83 : _GEN_567; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_569 = 7'h54 == total_offset_5[6:0] ? phv_data_84 : _GEN_568; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_570 = 7'h55 == total_offset_5[6:0] ? phv_data_85 : _GEN_569; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_571 = 7'h56 == total_offset_5[6:0] ? phv_data_86 : _GEN_570; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_572 = 7'h57 == total_offset_5[6:0] ? phv_data_87 : _GEN_571; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_573 = 7'h58 == total_offset_5[6:0] ? phv_data_88 : _GEN_572; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_574 = 7'h59 == total_offset_5[6:0] ? phv_data_89 : _GEN_573; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_575 = 7'h5a == total_offset_5[6:0] ? phv_data_90 : _GEN_574; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_576 = 7'h5b == total_offset_5[6:0] ? phv_data_91 : _GEN_575; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_577 = 7'h5c == total_offset_5[6:0] ? phv_data_92 : _GEN_576; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_578 = 7'h5d == total_offset_5[6:0] ? phv_data_93 : _GEN_577; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_579 = 7'h5e == total_offset_5[6:0] ? phv_data_94 : _GEN_578; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_580 = 7'h5f == total_offset_5[6:0] ? phv_data_95 : _GEN_579; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__5 = 8'h5 < length_0 ? _GEN_580 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_6 = offset_0 + 8'h6; // @[executor.scala 148:53]
  wire [7:0] _GEN_583 = 7'h1 == total_offset_6[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_584 = 7'h2 == total_offset_6[6:0] ? phv_data_2 : _GEN_583; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_585 = 7'h3 == total_offset_6[6:0] ? phv_data_3 : _GEN_584; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_586 = 7'h4 == total_offset_6[6:0] ? phv_data_4 : _GEN_585; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_587 = 7'h5 == total_offset_6[6:0] ? phv_data_5 : _GEN_586; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_588 = 7'h6 == total_offset_6[6:0] ? phv_data_6 : _GEN_587; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_589 = 7'h7 == total_offset_6[6:0] ? phv_data_7 : _GEN_588; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_590 = 7'h8 == total_offset_6[6:0] ? phv_data_8 : _GEN_589; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_591 = 7'h9 == total_offset_6[6:0] ? phv_data_9 : _GEN_590; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_592 = 7'ha == total_offset_6[6:0] ? phv_data_10 : _GEN_591; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_593 = 7'hb == total_offset_6[6:0] ? phv_data_11 : _GEN_592; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_594 = 7'hc == total_offset_6[6:0] ? phv_data_12 : _GEN_593; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_595 = 7'hd == total_offset_6[6:0] ? phv_data_13 : _GEN_594; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_596 = 7'he == total_offset_6[6:0] ? phv_data_14 : _GEN_595; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_597 = 7'hf == total_offset_6[6:0] ? phv_data_15 : _GEN_596; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_598 = 7'h10 == total_offset_6[6:0] ? phv_data_16 : _GEN_597; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_599 = 7'h11 == total_offset_6[6:0] ? phv_data_17 : _GEN_598; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_600 = 7'h12 == total_offset_6[6:0] ? phv_data_18 : _GEN_599; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_601 = 7'h13 == total_offset_6[6:0] ? phv_data_19 : _GEN_600; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_602 = 7'h14 == total_offset_6[6:0] ? phv_data_20 : _GEN_601; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_603 = 7'h15 == total_offset_6[6:0] ? phv_data_21 : _GEN_602; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_604 = 7'h16 == total_offset_6[6:0] ? phv_data_22 : _GEN_603; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_605 = 7'h17 == total_offset_6[6:0] ? phv_data_23 : _GEN_604; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_606 = 7'h18 == total_offset_6[6:0] ? phv_data_24 : _GEN_605; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_607 = 7'h19 == total_offset_6[6:0] ? phv_data_25 : _GEN_606; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_608 = 7'h1a == total_offset_6[6:0] ? phv_data_26 : _GEN_607; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_609 = 7'h1b == total_offset_6[6:0] ? phv_data_27 : _GEN_608; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_610 = 7'h1c == total_offset_6[6:0] ? phv_data_28 : _GEN_609; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_611 = 7'h1d == total_offset_6[6:0] ? phv_data_29 : _GEN_610; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_612 = 7'h1e == total_offset_6[6:0] ? phv_data_30 : _GEN_611; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_613 = 7'h1f == total_offset_6[6:0] ? phv_data_31 : _GEN_612; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_614 = 7'h20 == total_offset_6[6:0] ? phv_data_32 : _GEN_613; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_615 = 7'h21 == total_offset_6[6:0] ? phv_data_33 : _GEN_614; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_616 = 7'h22 == total_offset_6[6:0] ? phv_data_34 : _GEN_615; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_617 = 7'h23 == total_offset_6[6:0] ? phv_data_35 : _GEN_616; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_618 = 7'h24 == total_offset_6[6:0] ? phv_data_36 : _GEN_617; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_619 = 7'h25 == total_offset_6[6:0] ? phv_data_37 : _GEN_618; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_620 = 7'h26 == total_offset_6[6:0] ? phv_data_38 : _GEN_619; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_621 = 7'h27 == total_offset_6[6:0] ? phv_data_39 : _GEN_620; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_622 = 7'h28 == total_offset_6[6:0] ? phv_data_40 : _GEN_621; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_623 = 7'h29 == total_offset_6[6:0] ? phv_data_41 : _GEN_622; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_624 = 7'h2a == total_offset_6[6:0] ? phv_data_42 : _GEN_623; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_625 = 7'h2b == total_offset_6[6:0] ? phv_data_43 : _GEN_624; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_626 = 7'h2c == total_offset_6[6:0] ? phv_data_44 : _GEN_625; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_627 = 7'h2d == total_offset_6[6:0] ? phv_data_45 : _GEN_626; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_628 = 7'h2e == total_offset_6[6:0] ? phv_data_46 : _GEN_627; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_629 = 7'h2f == total_offset_6[6:0] ? phv_data_47 : _GEN_628; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_630 = 7'h30 == total_offset_6[6:0] ? phv_data_48 : _GEN_629; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_631 = 7'h31 == total_offset_6[6:0] ? phv_data_49 : _GEN_630; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_632 = 7'h32 == total_offset_6[6:0] ? phv_data_50 : _GEN_631; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_633 = 7'h33 == total_offset_6[6:0] ? phv_data_51 : _GEN_632; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_634 = 7'h34 == total_offset_6[6:0] ? phv_data_52 : _GEN_633; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_635 = 7'h35 == total_offset_6[6:0] ? phv_data_53 : _GEN_634; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_636 = 7'h36 == total_offset_6[6:0] ? phv_data_54 : _GEN_635; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_637 = 7'h37 == total_offset_6[6:0] ? phv_data_55 : _GEN_636; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_638 = 7'h38 == total_offset_6[6:0] ? phv_data_56 : _GEN_637; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_639 = 7'h39 == total_offset_6[6:0] ? phv_data_57 : _GEN_638; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_640 = 7'h3a == total_offset_6[6:0] ? phv_data_58 : _GEN_639; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_641 = 7'h3b == total_offset_6[6:0] ? phv_data_59 : _GEN_640; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_642 = 7'h3c == total_offset_6[6:0] ? phv_data_60 : _GEN_641; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_643 = 7'h3d == total_offset_6[6:0] ? phv_data_61 : _GEN_642; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_644 = 7'h3e == total_offset_6[6:0] ? phv_data_62 : _GEN_643; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_645 = 7'h3f == total_offset_6[6:0] ? phv_data_63 : _GEN_644; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_646 = 7'h40 == total_offset_6[6:0] ? phv_data_64 : _GEN_645; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_647 = 7'h41 == total_offset_6[6:0] ? phv_data_65 : _GEN_646; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_648 = 7'h42 == total_offset_6[6:0] ? phv_data_66 : _GEN_647; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_649 = 7'h43 == total_offset_6[6:0] ? phv_data_67 : _GEN_648; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_650 = 7'h44 == total_offset_6[6:0] ? phv_data_68 : _GEN_649; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_651 = 7'h45 == total_offset_6[6:0] ? phv_data_69 : _GEN_650; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_652 = 7'h46 == total_offset_6[6:0] ? phv_data_70 : _GEN_651; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_653 = 7'h47 == total_offset_6[6:0] ? phv_data_71 : _GEN_652; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_654 = 7'h48 == total_offset_6[6:0] ? phv_data_72 : _GEN_653; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_655 = 7'h49 == total_offset_6[6:0] ? phv_data_73 : _GEN_654; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_656 = 7'h4a == total_offset_6[6:0] ? phv_data_74 : _GEN_655; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_657 = 7'h4b == total_offset_6[6:0] ? phv_data_75 : _GEN_656; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_658 = 7'h4c == total_offset_6[6:0] ? phv_data_76 : _GEN_657; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_659 = 7'h4d == total_offset_6[6:0] ? phv_data_77 : _GEN_658; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_660 = 7'h4e == total_offset_6[6:0] ? phv_data_78 : _GEN_659; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_661 = 7'h4f == total_offset_6[6:0] ? phv_data_79 : _GEN_660; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_662 = 7'h50 == total_offset_6[6:0] ? phv_data_80 : _GEN_661; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_663 = 7'h51 == total_offset_6[6:0] ? phv_data_81 : _GEN_662; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_664 = 7'h52 == total_offset_6[6:0] ? phv_data_82 : _GEN_663; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_665 = 7'h53 == total_offset_6[6:0] ? phv_data_83 : _GEN_664; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_666 = 7'h54 == total_offset_6[6:0] ? phv_data_84 : _GEN_665; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_667 = 7'h55 == total_offset_6[6:0] ? phv_data_85 : _GEN_666; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_668 = 7'h56 == total_offset_6[6:0] ? phv_data_86 : _GEN_667; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_669 = 7'h57 == total_offset_6[6:0] ? phv_data_87 : _GEN_668; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_670 = 7'h58 == total_offset_6[6:0] ? phv_data_88 : _GEN_669; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_671 = 7'h59 == total_offset_6[6:0] ? phv_data_89 : _GEN_670; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_672 = 7'h5a == total_offset_6[6:0] ? phv_data_90 : _GEN_671; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_673 = 7'h5b == total_offset_6[6:0] ? phv_data_91 : _GEN_672; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_674 = 7'h5c == total_offset_6[6:0] ? phv_data_92 : _GEN_673; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_675 = 7'h5d == total_offset_6[6:0] ? phv_data_93 : _GEN_674; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_676 = 7'h5e == total_offset_6[6:0] ? phv_data_94 : _GEN_675; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_677 = 7'h5f == total_offset_6[6:0] ? phv_data_95 : _GEN_676; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__6 = 8'h6 < length_0 ? _GEN_677 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_7 = offset_0 + 8'h7; // @[executor.scala 148:53]
  wire [7:0] _GEN_680 = 7'h1 == total_offset_7[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_681 = 7'h2 == total_offset_7[6:0] ? phv_data_2 : _GEN_680; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_682 = 7'h3 == total_offset_7[6:0] ? phv_data_3 : _GEN_681; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_683 = 7'h4 == total_offset_7[6:0] ? phv_data_4 : _GEN_682; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_684 = 7'h5 == total_offset_7[6:0] ? phv_data_5 : _GEN_683; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_685 = 7'h6 == total_offset_7[6:0] ? phv_data_6 : _GEN_684; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_686 = 7'h7 == total_offset_7[6:0] ? phv_data_7 : _GEN_685; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_687 = 7'h8 == total_offset_7[6:0] ? phv_data_8 : _GEN_686; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_688 = 7'h9 == total_offset_7[6:0] ? phv_data_9 : _GEN_687; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_689 = 7'ha == total_offset_7[6:0] ? phv_data_10 : _GEN_688; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_690 = 7'hb == total_offset_7[6:0] ? phv_data_11 : _GEN_689; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_691 = 7'hc == total_offset_7[6:0] ? phv_data_12 : _GEN_690; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_692 = 7'hd == total_offset_7[6:0] ? phv_data_13 : _GEN_691; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_693 = 7'he == total_offset_7[6:0] ? phv_data_14 : _GEN_692; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_694 = 7'hf == total_offset_7[6:0] ? phv_data_15 : _GEN_693; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_695 = 7'h10 == total_offset_7[6:0] ? phv_data_16 : _GEN_694; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_696 = 7'h11 == total_offset_7[6:0] ? phv_data_17 : _GEN_695; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_697 = 7'h12 == total_offset_7[6:0] ? phv_data_18 : _GEN_696; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_698 = 7'h13 == total_offset_7[6:0] ? phv_data_19 : _GEN_697; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_699 = 7'h14 == total_offset_7[6:0] ? phv_data_20 : _GEN_698; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_700 = 7'h15 == total_offset_7[6:0] ? phv_data_21 : _GEN_699; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_701 = 7'h16 == total_offset_7[6:0] ? phv_data_22 : _GEN_700; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_702 = 7'h17 == total_offset_7[6:0] ? phv_data_23 : _GEN_701; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_703 = 7'h18 == total_offset_7[6:0] ? phv_data_24 : _GEN_702; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_704 = 7'h19 == total_offset_7[6:0] ? phv_data_25 : _GEN_703; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_705 = 7'h1a == total_offset_7[6:0] ? phv_data_26 : _GEN_704; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_706 = 7'h1b == total_offset_7[6:0] ? phv_data_27 : _GEN_705; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_707 = 7'h1c == total_offset_7[6:0] ? phv_data_28 : _GEN_706; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_708 = 7'h1d == total_offset_7[6:0] ? phv_data_29 : _GEN_707; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_709 = 7'h1e == total_offset_7[6:0] ? phv_data_30 : _GEN_708; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_710 = 7'h1f == total_offset_7[6:0] ? phv_data_31 : _GEN_709; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_711 = 7'h20 == total_offset_7[6:0] ? phv_data_32 : _GEN_710; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_712 = 7'h21 == total_offset_7[6:0] ? phv_data_33 : _GEN_711; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_713 = 7'h22 == total_offset_7[6:0] ? phv_data_34 : _GEN_712; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_714 = 7'h23 == total_offset_7[6:0] ? phv_data_35 : _GEN_713; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_715 = 7'h24 == total_offset_7[6:0] ? phv_data_36 : _GEN_714; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_716 = 7'h25 == total_offset_7[6:0] ? phv_data_37 : _GEN_715; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_717 = 7'h26 == total_offset_7[6:0] ? phv_data_38 : _GEN_716; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_718 = 7'h27 == total_offset_7[6:0] ? phv_data_39 : _GEN_717; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_719 = 7'h28 == total_offset_7[6:0] ? phv_data_40 : _GEN_718; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_720 = 7'h29 == total_offset_7[6:0] ? phv_data_41 : _GEN_719; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_721 = 7'h2a == total_offset_7[6:0] ? phv_data_42 : _GEN_720; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_722 = 7'h2b == total_offset_7[6:0] ? phv_data_43 : _GEN_721; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_723 = 7'h2c == total_offset_7[6:0] ? phv_data_44 : _GEN_722; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_724 = 7'h2d == total_offset_7[6:0] ? phv_data_45 : _GEN_723; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_725 = 7'h2e == total_offset_7[6:0] ? phv_data_46 : _GEN_724; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_726 = 7'h2f == total_offset_7[6:0] ? phv_data_47 : _GEN_725; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_727 = 7'h30 == total_offset_7[6:0] ? phv_data_48 : _GEN_726; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_728 = 7'h31 == total_offset_7[6:0] ? phv_data_49 : _GEN_727; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_729 = 7'h32 == total_offset_7[6:0] ? phv_data_50 : _GEN_728; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_730 = 7'h33 == total_offset_7[6:0] ? phv_data_51 : _GEN_729; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_731 = 7'h34 == total_offset_7[6:0] ? phv_data_52 : _GEN_730; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_732 = 7'h35 == total_offset_7[6:0] ? phv_data_53 : _GEN_731; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_733 = 7'h36 == total_offset_7[6:0] ? phv_data_54 : _GEN_732; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_734 = 7'h37 == total_offset_7[6:0] ? phv_data_55 : _GEN_733; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_735 = 7'h38 == total_offset_7[6:0] ? phv_data_56 : _GEN_734; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_736 = 7'h39 == total_offset_7[6:0] ? phv_data_57 : _GEN_735; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_737 = 7'h3a == total_offset_7[6:0] ? phv_data_58 : _GEN_736; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_738 = 7'h3b == total_offset_7[6:0] ? phv_data_59 : _GEN_737; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_739 = 7'h3c == total_offset_7[6:0] ? phv_data_60 : _GEN_738; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_740 = 7'h3d == total_offset_7[6:0] ? phv_data_61 : _GEN_739; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_741 = 7'h3e == total_offset_7[6:0] ? phv_data_62 : _GEN_740; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_742 = 7'h3f == total_offset_7[6:0] ? phv_data_63 : _GEN_741; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_743 = 7'h40 == total_offset_7[6:0] ? phv_data_64 : _GEN_742; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_744 = 7'h41 == total_offset_7[6:0] ? phv_data_65 : _GEN_743; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_745 = 7'h42 == total_offset_7[6:0] ? phv_data_66 : _GEN_744; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_746 = 7'h43 == total_offset_7[6:0] ? phv_data_67 : _GEN_745; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_747 = 7'h44 == total_offset_7[6:0] ? phv_data_68 : _GEN_746; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_748 = 7'h45 == total_offset_7[6:0] ? phv_data_69 : _GEN_747; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_749 = 7'h46 == total_offset_7[6:0] ? phv_data_70 : _GEN_748; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_750 = 7'h47 == total_offset_7[6:0] ? phv_data_71 : _GEN_749; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_751 = 7'h48 == total_offset_7[6:0] ? phv_data_72 : _GEN_750; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_752 = 7'h49 == total_offset_7[6:0] ? phv_data_73 : _GEN_751; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_753 = 7'h4a == total_offset_7[6:0] ? phv_data_74 : _GEN_752; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_754 = 7'h4b == total_offset_7[6:0] ? phv_data_75 : _GEN_753; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_755 = 7'h4c == total_offset_7[6:0] ? phv_data_76 : _GEN_754; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_756 = 7'h4d == total_offset_7[6:0] ? phv_data_77 : _GEN_755; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_757 = 7'h4e == total_offset_7[6:0] ? phv_data_78 : _GEN_756; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_758 = 7'h4f == total_offset_7[6:0] ? phv_data_79 : _GEN_757; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_759 = 7'h50 == total_offset_7[6:0] ? phv_data_80 : _GEN_758; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_760 = 7'h51 == total_offset_7[6:0] ? phv_data_81 : _GEN_759; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_761 = 7'h52 == total_offset_7[6:0] ? phv_data_82 : _GEN_760; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_762 = 7'h53 == total_offset_7[6:0] ? phv_data_83 : _GEN_761; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_763 = 7'h54 == total_offset_7[6:0] ? phv_data_84 : _GEN_762; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_764 = 7'h55 == total_offset_7[6:0] ? phv_data_85 : _GEN_763; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_765 = 7'h56 == total_offset_7[6:0] ? phv_data_86 : _GEN_764; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_766 = 7'h57 == total_offset_7[6:0] ? phv_data_87 : _GEN_765; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_767 = 7'h58 == total_offset_7[6:0] ? phv_data_88 : _GEN_766; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_768 = 7'h59 == total_offset_7[6:0] ? phv_data_89 : _GEN_767; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_769 = 7'h5a == total_offset_7[6:0] ? phv_data_90 : _GEN_768; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_770 = 7'h5b == total_offset_7[6:0] ? phv_data_91 : _GEN_769; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_771 = 7'h5c == total_offset_7[6:0] ? phv_data_92 : _GEN_770; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_772 = 7'h5d == total_offset_7[6:0] ? phv_data_93 : _GEN_771; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_773 = 7'h5e == total_offset_7[6:0] ? phv_data_94 : _GEN_772; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_774 = 7'h5f == total_offset_7[6:0] ? phv_data_95 : _GEN_773; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes__7 = 8'h7 < length_0 ? _GEN_774 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [63:0] _io_field_out_0_T = {bytes__0,bytes__1,bytes__2,bytes__3,bytes__4,bytes__5,bytes__6,bytes__7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset = io_field_out_0_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length = io_field_out_0_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_8 = {{6'd0}, args_offset}; // @[executor.scala 163:56]
  wire [7:0] total_offset_8 = _total_offset_T_8[7:0]; // @[executor.scala 163:56]
  wire [7:0] _GEN_3368 = {{5'd0}, args_length}; // @[executor.scala 164:44]
  wire [7:0] _GEN_777 = 3'h1 == total_offset_8[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_778 = 3'h2 == total_offset_8[2:0] ? args_2 : _GEN_777; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_779 = 3'h3 == total_offset_8[2:0] ? args_3 : _GEN_778; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_780 = 3'h4 == total_offset_8[2:0] ? args_4 : _GEN_779; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_781 = 3'h5 == total_offset_8[2:0] ? args_5 : _GEN_780; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_782 = 3'h6 == total_offset_8[2:0] ? args_6 : _GEN_781; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_1_0 = 8'h0 < _GEN_3368 ? _GEN_782 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] _GEN_3369 = {{5'd0}, args_offset}; // @[executor.scala 163:56]
  wire [7:0] total_offset_9 = _GEN_3369 + 8'h1; // @[executor.scala 163:56]
  wire [7:0] _GEN_785 = 3'h1 == total_offset_9[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_786 = 3'h2 == total_offset_9[2:0] ? args_2 : _GEN_785; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_787 = 3'h3 == total_offset_9[2:0] ? args_3 : _GEN_786; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_788 = 3'h4 == total_offset_9[2:0] ? args_4 : _GEN_787; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_789 = 3'h5 == total_offset_9[2:0] ? args_5 : _GEN_788; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_790 = 3'h6 == total_offset_9[2:0] ? args_6 : _GEN_789; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_1_1 = 8'h1 < _GEN_3368 ? _GEN_790 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_10 = _GEN_3369 + 8'h2; // @[executor.scala 163:56]
  wire [7:0] _GEN_793 = 3'h1 == total_offset_10[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_794 = 3'h2 == total_offset_10[2:0] ? args_2 : _GEN_793; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_795 = 3'h3 == total_offset_10[2:0] ? args_3 : _GEN_794; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_796 = 3'h4 == total_offset_10[2:0] ? args_4 : _GEN_795; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_797 = 3'h5 == total_offset_10[2:0] ? args_5 : _GEN_796; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_798 = 3'h6 == total_offset_10[2:0] ? args_6 : _GEN_797; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_1_2 = 8'h2 < _GEN_3368 ? _GEN_798 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_11 = _GEN_3369 + 8'h3; // @[executor.scala 163:56]
  wire [7:0] _GEN_801 = 3'h1 == total_offset_11[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_802 = 3'h2 == total_offset_11[2:0] ? args_2 : _GEN_801; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_803 = 3'h3 == total_offset_11[2:0] ? args_3 : _GEN_802; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_804 = 3'h4 == total_offset_11[2:0] ? args_4 : _GEN_803; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_805 = 3'h5 == total_offset_11[2:0] ? args_5 : _GEN_804; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_806 = 3'h6 == total_offset_11[2:0] ? args_6 : _GEN_805; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_1_3 = 8'h3 < _GEN_3368 ? _GEN_806 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_12 = _GEN_3369 + 8'h4; // @[executor.scala 163:56]
  wire [7:0] _GEN_809 = 3'h1 == total_offset_12[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_810 = 3'h2 == total_offset_12[2:0] ? args_2 : _GEN_809; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_811 = 3'h3 == total_offset_12[2:0] ? args_3 : _GEN_810; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_812 = 3'h4 == total_offset_12[2:0] ? args_4 : _GEN_811; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_813 = 3'h5 == total_offset_12[2:0] ? args_5 : _GEN_812; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_814 = 3'h6 == total_offset_12[2:0] ? args_6 : _GEN_813; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_1_4 = 8'h4 < _GEN_3368 ? _GEN_814 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_13 = _GEN_3369 + 8'h5; // @[executor.scala 163:56]
  wire [7:0] _GEN_817 = 3'h1 == total_offset_13[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_818 = 3'h2 == total_offset_13[2:0] ? args_2 : _GEN_817; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_819 = 3'h3 == total_offset_13[2:0] ? args_3 : _GEN_818; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_820 = 3'h4 == total_offset_13[2:0] ? args_4 : _GEN_819; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_821 = 3'h5 == total_offset_13[2:0] ? args_5 : _GEN_820; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_822 = 3'h6 == total_offset_13[2:0] ? args_6 : _GEN_821; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_1_5 = 8'h5 < _GEN_3368 ? _GEN_822 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_14 = _GEN_3369 + 8'h6; // @[executor.scala 163:56]
  wire [7:0] _GEN_825 = 3'h1 == total_offset_14[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_826 = 3'h2 == total_offset_14[2:0] ? args_2 : _GEN_825; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_827 = 3'h3 == total_offset_14[2:0] ? args_3 : _GEN_826; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_828 = 3'h4 == total_offset_14[2:0] ? args_4 : _GEN_827; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_829 = 3'h5 == total_offset_14[2:0] ? args_5 : _GEN_828; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_830 = 3'h6 == total_offset_14[2:0] ? args_6 : _GEN_829; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_1_6 = 8'h6 < _GEN_3368 ? _GEN_830 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [63:0] _io_field_out_0_T_1 = {bytes_1_0,bytes_1_1,bytes_1_2,bytes_1_3,bytes_1_4,bytes_1_5,bytes_1_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_0_hi_12 = io_field_out_0_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_0_T_4 = {io_field_out_0_hi_12,io_field_out_0_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_840 = 4'ha == opcode ? _io_field_out_0_T_1 : _io_field_out_0_T_4; // @[executor.scala 157:51 executor.scala 170:37 executor.scala 173:37]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_1_lo = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire  from_header_1 = length_1 != 8'h0; // @[executor.scala 141:41]
  wire [8:0] _total_offset_T_16 = {{1'd0}, offset_1}; // @[executor.scala 148:53]
  wire [7:0] total_offset_16 = _total_offset_T_16[7:0]; // @[executor.scala 148:53]
  wire [7:0] _GEN_843 = 7'h1 == total_offset_16[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_844 = 7'h2 == total_offset_16[6:0] ? phv_data_2 : _GEN_843; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_845 = 7'h3 == total_offset_16[6:0] ? phv_data_3 : _GEN_844; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_846 = 7'h4 == total_offset_16[6:0] ? phv_data_4 : _GEN_845; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_847 = 7'h5 == total_offset_16[6:0] ? phv_data_5 : _GEN_846; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_848 = 7'h6 == total_offset_16[6:0] ? phv_data_6 : _GEN_847; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_849 = 7'h7 == total_offset_16[6:0] ? phv_data_7 : _GEN_848; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_850 = 7'h8 == total_offset_16[6:0] ? phv_data_8 : _GEN_849; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_851 = 7'h9 == total_offset_16[6:0] ? phv_data_9 : _GEN_850; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_852 = 7'ha == total_offset_16[6:0] ? phv_data_10 : _GEN_851; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_853 = 7'hb == total_offset_16[6:0] ? phv_data_11 : _GEN_852; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_854 = 7'hc == total_offset_16[6:0] ? phv_data_12 : _GEN_853; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_855 = 7'hd == total_offset_16[6:0] ? phv_data_13 : _GEN_854; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_856 = 7'he == total_offset_16[6:0] ? phv_data_14 : _GEN_855; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_857 = 7'hf == total_offset_16[6:0] ? phv_data_15 : _GEN_856; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_858 = 7'h10 == total_offset_16[6:0] ? phv_data_16 : _GEN_857; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_859 = 7'h11 == total_offset_16[6:0] ? phv_data_17 : _GEN_858; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_860 = 7'h12 == total_offset_16[6:0] ? phv_data_18 : _GEN_859; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_861 = 7'h13 == total_offset_16[6:0] ? phv_data_19 : _GEN_860; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_862 = 7'h14 == total_offset_16[6:0] ? phv_data_20 : _GEN_861; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_863 = 7'h15 == total_offset_16[6:0] ? phv_data_21 : _GEN_862; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_864 = 7'h16 == total_offset_16[6:0] ? phv_data_22 : _GEN_863; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_865 = 7'h17 == total_offset_16[6:0] ? phv_data_23 : _GEN_864; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_866 = 7'h18 == total_offset_16[6:0] ? phv_data_24 : _GEN_865; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_867 = 7'h19 == total_offset_16[6:0] ? phv_data_25 : _GEN_866; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_868 = 7'h1a == total_offset_16[6:0] ? phv_data_26 : _GEN_867; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_869 = 7'h1b == total_offset_16[6:0] ? phv_data_27 : _GEN_868; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_870 = 7'h1c == total_offset_16[6:0] ? phv_data_28 : _GEN_869; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_871 = 7'h1d == total_offset_16[6:0] ? phv_data_29 : _GEN_870; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_872 = 7'h1e == total_offset_16[6:0] ? phv_data_30 : _GEN_871; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_873 = 7'h1f == total_offset_16[6:0] ? phv_data_31 : _GEN_872; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_874 = 7'h20 == total_offset_16[6:0] ? phv_data_32 : _GEN_873; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_875 = 7'h21 == total_offset_16[6:0] ? phv_data_33 : _GEN_874; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_876 = 7'h22 == total_offset_16[6:0] ? phv_data_34 : _GEN_875; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_877 = 7'h23 == total_offset_16[6:0] ? phv_data_35 : _GEN_876; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_878 = 7'h24 == total_offset_16[6:0] ? phv_data_36 : _GEN_877; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_879 = 7'h25 == total_offset_16[6:0] ? phv_data_37 : _GEN_878; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_880 = 7'h26 == total_offset_16[6:0] ? phv_data_38 : _GEN_879; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_881 = 7'h27 == total_offset_16[6:0] ? phv_data_39 : _GEN_880; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_882 = 7'h28 == total_offset_16[6:0] ? phv_data_40 : _GEN_881; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_883 = 7'h29 == total_offset_16[6:0] ? phv_data_41 : _GEN_882; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_884 = 7'h2a == total_offset_16[6:0] ? phv_data_42 : _GEN_883; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_885 = 7'h2b == total_offset_16[6:0] ? phv_data_43 : _GEN_884; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_886 = 7'h2c == total_offset_16[6:0] ? phv_data_44 : _GEN_885; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_887 = 7'h2d == total_offset_16[6:0] ? phv_data_45 : _GEN_886; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_888 = 7'h2e == total_offset_16[6:0] ? phv_data_46 : _GEN_887; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_889 = 7'h2f == total_offset_16[6:0] ? phv_data_47 : _GEN_888; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_890 = 7'h30 == total_offset_16[6:0] ? phv_data_48 : _GEN_889; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_891 = 7'h31 == total_offset_16[6:0] ? phv_data_49 : _GEN_890; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_892 = 7'h32 == total_offset_16[6:0] ? phv_data_50 : _GEN_891; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_893 = 7'h33 == total_offset_16[6:0] ? phv_data_51 : _GEN_892; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_894 = 7'h34 == total_offset_16[6:0] ? phv_data_52 : _GEN_893; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_895 = 7'h35 == total_offset_16[6:0] ? phv_data_53 : _GEN_894; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_896 = 7'h36 == total_offset_16[6:0] ? phv_data_54 : _GEN_895; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_897 = 7'h37 == total_offset_16[6:0] ? phv_data_55 : _GEN_896; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_898 = 7'h38 == total_offset_16[6:0] ? phv_data_56 : _GEN_897; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_899 = 7'h39 == total_offset_16[6:0] ? phv_data_57 : _GEN_898; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_900 = 7'h3a == total_offset_16[6:0] ? phv_data_58 : _GEN_899; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_901 = 7'h3b == total_offset_16[6:0] ? phv_data_59 : _GEN_900; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_902 = 7'h3c == total_offset_16[6:0] ? phv_data_60 : _GEN_901; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_903 = 7'h3d == total_offset_16[6:0] ? phv_data_61 : _GEN_902; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_904 = 7'h3e == total_offset_16[6:0] ? phv_data_62 : _GEN_903; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_905 = 7'h3f == total_offset_16[6:0] ? phv_data_63 : _GEN_904; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_906 = 7'h40 == total_offset_16[6:0] ? phv_data_64 : _GEN_905; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_907 = 7'h41 == total_offset_16[6:0] ? phv_data_65 : _GEN_906; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_908 = 7'h42 == total_offset_16[6:0] ? phv_data_66 : _GEN_907; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_909 = 7'h43 == total_offset_16[6:0] ? phv_data_67 : _GEN_908; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_910 = 7'h44 == total_offset_16[6:0] ? phv_data_68 : _GEN_909; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_911 = 7'h45 == total_offset_16[6:0] ? phv_data_69 : _GEN_910; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_912 = 7'h46 == total_offset_16[6:0] ? phv_data_70 : _GEN_911; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_913 = 7'h47 == total_offset_16[6:0] ? phv_data_71 : _GEN_912; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_914 = 7'h48 == total_offset_16[6:0] ? phv_data_72 : _GEN_913; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_915 = 7'h49 == total_offset_16[6:0] ? phv_data_73 : _GEN_914; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_916 = 7'h4a == total_offset_16[6:0] ? phv_data_74 : _GEN_915; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_917 = 7'h4b == total_offset_16[6:0] ? phv_data_75 : _GEN_916; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_918 = 7'h4c == total_offset_16[6:0] ? phv_data_76 : _GEN_917; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_919 = 7'h4d == total_offset_16[6:0] ? phv_data_77 : _GEN_918; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_920 = 7'h4e == total_offset_16[6:0] ? phv_data_78 : _GEN_919; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_921 = 7'h4f == total_offset_16[6:0] ? phv_data_79 : _GEN_920; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_922 = 7'h50 == total_offset_16[6:0] ? phv_data_80 : _GEN_921; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_923 = 7'h51 == total_offset_16[6:0] ? phv_data_81 : _GEN_922; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_924 = 7'h52 == total_offset_16[6:0] ? phv_data_82 : _GEN_923; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_925 = 7'h53 == total_offset_16[6:0] ? phv_data_83 : _GEN_924; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_926 = 7'h54 == total_offset_16[6:0] ? phv_data_84 : _GEN_925; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_927 = 7'h55 == total_offset_16[6:0] ? phv_data_85 : _GEN_926; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_928 = 7'h56 == total_offset_16[6:0] ? phv_data_86 : _GEN_927; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_929 = 7'h57 == total_offset_16[6:0] ? phv_data_87 : _GEN_928; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_930 = 7'h58 == total_offset_16[6:0] ? phv_data_88 : _GEN_929; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_931 = 7'h59 == total_offset_16[6:0] ? phv_data_89 : _GEN_930; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_932 = 7'h5a == total_offset_16[6:0] ? phv_data_90 : _GEN_931; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_933 = 7'h5b == total_offset_16[6:0] ? phv_data_91 : _GEN_932; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_934 = 7'h5c == total_offset_16[6:0] ? phv_data_92 : _GEN_933; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_935 = 7'h5d == total_offset_16[6:0] ? phv_data_93 : _GEN_934; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_936 = 7'h5e == total_offset_16[6:0] ? phv_data_94 : _GEN_935; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_937 = 7'h5f == total_offset_16[6:0] ? phv_data_95 : _GEN_936; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_0 = 8'h0 < length_1 ? _GEN_937 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_17 = offset_1 + 8'h1; // @[executor.scala 148:53]
  wire [7:0] _GEN_940 = 7'h1 == total_offset_17[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_941 = 7'h2 == total_offset_17[6:0] ? phv_data_2 : _GEN_940; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_942 = 7'h3 == total_offset_17[6:0] ? phv_data_3 : _GEN_941; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_943 = 7'h4 == total_offset_17[6:0] ? phv_data_4 : _GEN_942; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_944 = 7'h5 == total_offset_17[6:0] ? phv_data_5 : _GEN_943; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_945 = 7'h6 == total_offset_17[6:0] ? phv_data_6 : _GEN_944; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_946 = 7'h7 == total_offset_17[6:0] ? phv_data_7 : _GEN_945; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_947 = 7'h8 == total_offset_17[6:0] ? phv_data_8 : _GEN_946; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_948 = 7'h9 == total_offset_17[6:0] ? phv_data_9 : _GEN_947; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_949 = 7'ha == total_offset_17[6:0] ? phv_data_10 : _GEN_948; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_950 = 7'hb == total_offset_17[6:0] ? phv_data_11 : _GEN_949; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_951 = 7'hc == total_offset_17[6:0] ? phv_data_12 : _GEN_950; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_952 = 7'hd == total_offset_17[6:0] ? phv_data_13 : _GEN_951; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_953 = 7'he == total_offset_17[6:0] ? phv_data_14 : _GEN_952; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_954 = 7'hf == total_offset_17[6:0] ? phv_data_15 : _GEN_953; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_955 = 7'h10 == total_offset_17[6:0] ? phv_data_16 : _GEN_954; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_956 = 7'h11 == total_offset_17[6:0] ? phv_data_17 : _GEN_955; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_957 = 7'h12 == total_offset_17[6:0] ? phv_data_18 : _GEN_956; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_958 = 7'h13 == total_offset_17[6:0] ? phv_data_19 : _GEN_957; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_959 = 7'h14 == total_offset_17[6:0] ? phv_data_20 : _GEN_958; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_960 = 7'h15 == total_offset_17[6:0] ? phv_data_21 : _GEN_959; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_961 = 7'h16 == total_offset_17[6:0] ? phv_data_22 : _GEN_960; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_962 = 7'h17 == total_offset_17[6:0] ? phv_data_23 : _GEN_961; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_963 = 7'h18 == total_offset_17[6:0] ? phv_data_24 : _GEN_962; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_964 = 7'h19 == total_offset_17[6:0] ? phv_data_25 : _GEN_963; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_965 = 7'h1a == total_offset_17[6:0] ? phv_data_26 : _GEN_964; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_966 = 7'h1b == total_offset_17[6:0] ? phv_data_27 : _GEN_965; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_967 = 7'h1c == total_offset_17[6:0] ? phv_data_28 : _GEN_966; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_968 = 7'h1d == total_offset_17[6:0] ? phv_data_29 : _GEN_967; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_969 = 7'h1e == total_offset_17[6:0] ? phv_data_30 : _GEN_968; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_970 = 7'h1f == total_offset_17[6:0] ? phv_data_31 : _GEN_969; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_971 = 7'h20 == total_offset_17[6:0] ? phv_data_32 : _GEN_970; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_972 = 7'h21 == total_offset_17[6:0] ? phv_data_33 : _GEN_971; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_973 = 7'h22 == total_offset_17[6:0] ? phv_data_34 : _GEN_972; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_974 = 7'h23 == total_offset_17[6:0] ? phv_data_35 : _GEN_973; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_975 = 7'h24 == total_offset_17[6:0] ? phv_data_36 : _GEN_974; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_976 = 7'h25 == total_offset_17[6:0] ? phv_data_37 : _GEN_975; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_977 = 7'h26 == total_offset_17[6:0] ? phv_data_38 : _GEN_976; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_978 = 7'h27 == total_offset_17[6:0] ? phv_data_39 : _GEN_977; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_979 = 7'h28 == total_offset_17[6:0] ? phv_data_40 : _GEN_978; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_980 = 7'h29 == total_offset_17[6:0] ? phv_data_41 : _GEN_979; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_981 = 7'h2a == total_offset_17[6:0] ? phv_data_42 : _GEN_980; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_982 = 7'h2b == total_offset_17[6:0] ? phv_data_43 : _GEN_981; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_983 = 7'h2c == total_offset_17[6:0] ? phv_data_44 : _GEN_982; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_984 = 7'h2d == total_offset_17[6:0] ? phv_data_45 : _GEN_983; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_985 = 7'h2e == total_offset_17[6:0] ? phv_data_46 : _GEN_984; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_986 = 7'h2f == total_offset_17[6:0] ? phv_data_47 : _GEN_985; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_987 = 7'h30 == total_offset_17[6:0] ? phv_data_48 : _GEN_986; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_988 = 7'h31 == total_offset_17[6:0] ? phv_data_49 : _GEN_987; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_989 = 7'h32 == total_offset_17[6:0] ? phv_data_50 : _GEN_988; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_990 = 7'h33 == total_offset_17[6:0] ? phv_data_51 : _GEN_989; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_991 = 7'h34 == total_offset_17[6:0] ? phv_data_52 : _GEN_990; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_992 = 7'h35 == total_offset_17[6:0] ? phv_data_53 : _GEN_991; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_993 = 7'h36 == total_offset_17[6:0] ? phv_data_54 : _GEN_992; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_994 = 7'h37 == total_offset_17[6:0] ? phv_data_55 : _GEN_993; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_995 = 7'h38 == total_offset_17[6:0] ? phv_data_56 : _GEN_994; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_996 = 7'h39 == total_offset_17[6:0] ? phv_data_57 : _GEN_995; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_997 = 7'h3a == total_offset_17[6:0] ? phv_data_58 : _GEN_996; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_998 = 7'h3b == total_offset_17[6:0] ? phv_data_59 : _GEN_997; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_999 = 7'h3c == total_offset_17[6:0] ? phv_data_60 : _GEN_998; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1000 = 7'h3d == total_offset_17[6:0] ? phv_data_61 : _GEN_999; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1001 = 7'h3e == total_offset_17[6:0] ? phv_data_62 : _GEN_1000; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1002 = 7'h3f == total_offset_17[6:0] ? phv_data_63 : _GEN_1001; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1003 = 7'h40 == total_offset_17[6:0] ? phv_data_64 : _GEN_1002; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1004 = 7'h41 == total_offset_17[6:0] ? phv_data_65 : _GEN_1003; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1005 = 7'h42 == total_offset_17[6:0] ? phv_data_66 : _GEN_1004; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1006 = 7'h43 == total_offset_17[6:0] ? phv_data_67 : _GEN_1005; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1007 = 7'h44 == total_offset_17[6:0] ? phv_data_68 : _GEN_1006; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1008 = 7'h45 == total_offset_17[6:0] ? phv_data_69 : _GEN_1007; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1009 = 7'h46 == total_offset_17[6:0] ? phv_data_70 : _GEN_1008; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1010 = 7'h47 == total_offset_17[6:0] ? phv_data_71 : _GEN_1009; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1011 = 7'h48 == total_offset_17[6:0] ? phv_data_72 : _GEN_1010; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1012 = 7'h49 == total_offset_17[6:0] ? phv_data_73 : _GEN_1011; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1013 = 7'h4a == total_offset_17[6:0] ? phv_data_74 : _GEN_1012; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1014 = 7'h4b == total_offset_17[6:0] ? phv_data_75 : _GEN_1013; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1015 = 7'h4c == total_offset_17[6:0] ? phv_data_76 : _GEN_1014; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1016 = 7'h4d == total_offset_17[6:0] ? phv_data_77 : _GEN_1015; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1017 = 7'h4e == total_offset_17[6:0] ? phv_data_78 : _GEN_1016; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1018 = 7'h4f == total_offset_17[6:0] ? phv_data_79 : _GEN_1017; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1019 = 7'h50 == total_offset_17[6:0] ? phv_data_80 : _GEN_1018; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1020 = 7'h51 == total_offset_17[6:0] ? phv_data_81 : _GEN_1019; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1021 = 7'h52 == total_offset_17[6:0] ? phv_data_82 : _GEN_1020; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1022 = 7'h53 == total_offset_17[6:0] ? phv_data_83 : _GEN_1021; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1023 = 7'h54 == total_offset_17[6:0] ? phv_data_84 : _GEN_1022; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1024 = 7'h55 == total_offset_17[6:0] ? phv_data_85 : _GEN_1023; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1025 = 7'h56 == total_offset_17[6:0] ? phv_data_86 : _GEN_1024; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1026 = 7'h57 == total_offset_17[6:0] ? phv_data_87 : _GEN_1025; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1027 = 7'h58 == total_offset_17[6:0] ? phv_data_88 : _GEN_1026; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1028 = 7'h59 == total_offset_17[6:0] ? phv_data_89 : _GEN_1027; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1029 = 7'h5a == total_offset_17[6:0] ? phv_data_90 : _GEN_1028; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1030 = 7'h5b == total_offset_17[6:0] ? phv_data_91 : _GEN_1029; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1031 = 7'h5c == total_offset_17[6:0] ? phv_data_92 : _GEN_1030; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1032 = 7'h5d == total_offset_17[6:0] ? phv_data_93 : _GEN_1031; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1033 = 7'h5e == total_offset_17[6:0] ? phv_data_94 : _GEN_1032; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1034 = 7'h5f == total_offset_17[6:0] ? phv_data_95 : _GEN_1033; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_1 = 8'h1 < length_1 ? _GEN_1034 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_18 = offset_1 + 8'h2; // @[executor.scala 148:53]
  wire [7:0] _GEN_1037 = 7'h1 == total_offset_18[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1038 = 7'h2 == total_offset_18[6:0] ? phv_data_2 : _GEN_1037; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1039 = 7'h3 == total_offset_18[6:0] ? phv_data_3 : _GEN_1038; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1040 = 7'h4 == total_offset_18[6:0] ? phv_data_4 : _GEN_1039; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1041 = 7'h5 == total_offset_18[6:0] ? phv_data_5 : _GEN_1040; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1042 = 7'h6 == total_offset_18[6:0] ? phv_data_6 : _GEN_1041; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1043 = 7'h7 == total_offset_18[6:0] ? phv_data_7 : _GEN_1042; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1044 = 7'h8 == total_offset_18[6:0] ? phv_data_8 : _GEN_1043; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1045 = 7'h9 == total_offset_18[6:0] ? phv_data_9 : _GEN_1044; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1046 = 7'ha == total_offset_18[6:0] ? phv_data_10 : _GEN_1045; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1047 = 7'hb == total_offset_18[6:0] ? phv_data_11 : _GEN_1046; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1048 = 7'hc == total_offset_18[6:0] ? phv_data_12 : _GEN_1047; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1049 = 7'hd == total_offset_18[6:0] ? phv_data_13 : _GEN_1048; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1050 = 7'he == total_offset_18[6:0] ? phv_data_14 : _GEN_1049; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1051 = 7'hf == total_offset_18[6:0] ? phv_data_15 : _GEN_1050; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1052 = 7'h10 == total_offset_18[6:0] ? phv_data_16 : _GEN_1051; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1053 = 7'h11 == total_offset_18[6:0] ? phv_data_17 : _GEN_1052; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1054 = 7'h12 == total_offset_18[6:0] ? phv_data_18 : _GEN_1053; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1055 = 7'h13 == total_offset_18[6:0] ? phv_data_19 : _GEN_1054; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1056 = 7'h14 == total_offset_18[6:0] ? phv_data_20 : _GEN_1055; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1057 = 7'h15 == total_offset_18[6:0] ? phv_data_21 : _GEN_1056; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1058 = 7'h16 == total_offset_18[6:0] ? phv_data_22 : _GEN_1057; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1059 = 7'h17 == total_offset_18[6:0] ? phv_data_23 : _GEN_1058; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1060 = 7'h18 == total_offset_18[6:0] ? phv_data_24 : _GEN_1059; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1061 = 7'h19 == total_offset_18[6:0] ? phv_data_25 : _GEN_1060; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1062 = 7'h1a == total_offset_18[6:0] ? phv_data_26 : _GEN_1061; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1063 = 7'h1b == total_offset_18[6:0] ? phv_data_27 : _GEN_1062; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1064 = 7'h1c == total_offset_18[6:0] ? phv_data_28 : _GEN_1063; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1065 = 7'h1d == total_offset_18[6:0] ? phv_data_29 : _GEN_1064; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1066 = 7'h1e == total_offset_18[6:0] ? phv_data_30 : _GEN_1065; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1067 = 7'h1f == total_offset_18[6:0] ? phv_data_31 : _GEN_1066; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1068 = 7'h20 == total_offset_18[6:0] ? phv_data_32 : _GEN_1067; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1069 = 7'h21 == total_offset_18[6:0] ? phv_data_33 : _GEN_1068; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1070 = 7'h22 == total_offset_18[6:0] ? phv_data_34 : _GEN_1069; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1071 = 7'h23 == total_offset_18[6:0] ? phv_data_35 : _GEN_1070; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1072 = 7'h24 == total_offset_18[6:0] ? phv_data_36 : _GEN_1071; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1073 = 7'h25 == total_offset_18[6:0] ? phv_data_37 : _GEN_1072; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1074 = 7'h26 == total_offset_18[6:0] ? phv_data_38 : _GEN_1073; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1075 = 7'h27 == total_offset_18[6:0] ? phv_data_39 : _GEN_1074; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1076 = 7'h28 == total_offset_18[6:0] ? phv_data_40 : _GEN_1075; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1077 = 7'h29 == total_offset_18[6:0] ? phv_data_41 : _GEN_1076; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1078 = 7'h2a == total_offset_18[6:0] ? phv_data_42 : _GEN_1077; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1079 = 7'h2b == total_offset_18[6:0] ? phv_data_43 : _GEN_1078; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1080 = 7'h2c == total_offset_18[6:0] ? phv_data_44 : _GEN_1079; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1081 = 7'h2d == total_offset_18[6:0] ? phv_data_45 : _GEN_1080; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1082 = 7'h2e == total_offset_18[6:0] ? phv_data_46 : _GEN_1081; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1083 = 7'h2f == total_offset_18[6:0] ? phv_data_47 : _GEN_1082; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1084 = 7'h30 == total_offset_18[6:0] ? phv_data_48 : _GEN_1083; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1085 = 7'h31 == total_offset_18[6:0] ? phv_data_49 : _GEN_1084; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1086 = 7'h32 == total_offset_18[6:0] ? phv_data_50 : _GEN_1085; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1087 = 7'h33 == total_offset_18[6:0] ? phv_data_51 : _GEN_1086; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1088 = 7'h34 == total_offset_18[6:0] ? phv_data_52 : _GEN_1087; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1089 = 7'h35 == total_offset_18[6:0] ? phv_data_53 : _GEN_1088; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1090 = 7'h36 == total_offset_18[6:0] ? phv_data_54 : _GEN_1089; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1091 = 7'h37 == total_offset_18[6:0] ? phv_data_55 : _GEN_1090; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1092 = 7'h38 == total_offset_18[6:0] ? phv_data_56 : _GEN_1091; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1093 = 7'h39 == total_offset_18[6:0] ? phv_data_57 : _GEN_1092; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1094 = 7'h3a == total_offset_18[6:0] ? phv_data_58 : _GEN_1093; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1095 = 7'h3b == total_offset_18[6:0] ? phv_data_59 : _GEN_1094; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1096 = 7'h3c == total_offset_18[6:0] ? phv_data_60 : _GEN_1095; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1097 = 7'h3d == total_offset_18[6:0] ? phv_data_61 : _GEN_1096; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1098 = 7'h3e == total_offset_18[6:0] ? phv_data_62 : _GEN_1097; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1099 = 7'h3f == total_offset_18[6:0] ? phv_data_63 : _GEN_1098; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1100 = 7'h40 == total_offset_18[6:0] ? phv_data_64 : _GEN_1099; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1101 = 7'h41 == total_offset_18[6:0] ? phv_data_65 : _GEN_1100; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1102 = 7'h42 == total_offset_18[6:0] ? phv_data_66 : _GEN_1101; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1103 = 7'h43 == total_offset_18[6:0] ? phv_data_67 : _GEN_1102; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1104 = 7'h44 == total_offset_18[6:0] ? phv_data_68 : _GEN_1103; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1105 = 7'h45 == total_offset_18[6:0] ? phv_data_69 : _GEN_1104; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1106 = 7'h46 == total_offset_18[6:0] ? phv_data_70 : _GEN_1105; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1107 = 7'h47 == total_offset_18[6:0] ? phv_data_71 : _GEN_1106; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1108 = 7'h48 == total_offset_18[6:0] ? phv_data_72 : _GEN_1107; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1109 = 7'h49 == total_offset_18[6:0] ? phv_data_73 : _GEN_1108; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1110 = 7'h4a == total_offset_18[6:0] ? phv_data_74 : _GEN_1109; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1111 = 7'h4b == total_offset_18[6:0] ? phv_data_75 : _GEN_1110; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1112 = 7'h4c == total_offset_18[6:0] ? phv_data_76 : _GEN_1111; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1113 = 7'h4d == total_offset_18[6:0] ? phv_data_77 : _GEN_1112; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1114 = 7'h4e == total_offset_18[6:0] ? phv_data_78 : _GEN_1113; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1115 = 7'h4f == total_offset_18[6:0] ? phv_data_79 : _GEN_1114; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1116 = 7'h50 == total_offset_18[6:0] ? phv_data_80 : _GEN_1115; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1117 = 7'h51 == total_offset_18[6:0] ? phv_data_81 : _GEN_1116; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1118 = 7'h52 == total_offset_18[6:0] ? phv_data_82 : _GEN_1117; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1119 = 7'h53 == total_offset_18[6:0] ? phv_data_83 : _GEN_1118; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1120 = 7'h54 == total_offset_18[6:0] ? phv_data_84 : _GEN_1119; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1121 = 7'h55 == total_offset_18[6:0] ? phv_data_85 : _GEN_1120; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1122 = 7'h56 == total_offset_18[6:0] ? phv_data_86 : _GEN_1121; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1123 = 7'h57 == total_offset_18[6:0] ? phv_data_87 : _GEN_1122; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1124 = 7'h58 == total_offset_18[6:0] ? phv_data_88 : _GEN_1123; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1125 = 7'h59 == total_offset_18[6:0] ? phv_data_89 : _GEN_1124; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1126 = 7'h5a == total_offset_18[6:0] ? phv_data_90 : _GEN_1125; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1127 = 7'h5b == total_offset_18[6:0] ? phv_data_91 : _GEN_1126; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1128 = 7'h5c == total_offset_18[6:0] ? phv_data_92 : _GEN_1127; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1129 = 7'h5d == total_offset_18[6:0] ? phv_data_93 : _GEN_1128; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1130 = 7'h5e == total_offset_18[6:0] ? phv_data_94 : _GEN_1129; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1131 = 7'h5f == total_offset_18[6:0] ? phv_data_95 : _GEN_1130; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_2 = 8'h2 < length_1 ? _GEN_1131 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_19 = offset_1 + 8'h3; // @[executor.scala 148:53]
  wire [7:0] _GEN_1134 = 7'h1 == total_offset_19[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1135 = 7'h2 == total_offset_19[6:0] ? phv_data_2 : _GEN_1134; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1136 = 7'h3 == total_offset_19[6:0] ? phv_data_3 : _GEN_1135; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1137 = 7'h4 == total_offset_19[6:0] ? phv_data_4 : _GEN_1136; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1138 = 7'h5 == total_offset_19[6:0] ? phv_data_5 : _GEN_1137; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1139 = 7'h6 == total_offset_19[6:0] ? phv_data_6 : _GEN_1138; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1140 = 7'h7 == total_offset_19[6:0] ? phv_data_7 : _GEN_1139; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1141 = 7'h8 == total_offset_19[6:0] ? phv_data_8 : _GEN_1140; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1142 = 7'h9 == total_offset_19[6:0] ? phv_data_9 : _GEN_1141; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1143 = 7'ha == total_offset_19[6:0] ? phv_data_10 : _GEN_1142; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1144 = 7'hb == total_offset_19[6:0] ? phv_data_11 : _GEN_1143; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1145 = 7'hc == total_offset_19[6:0] ? phv_data_12 : _GEN_1144; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1146 = 7'hd == total_offset_19[6:0] ? phv_data_13 : _GEN_1145; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1147 = 7'he == total_offset_19[6:0] ? phv_data_14 : _GEN_1146; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1148 = 7'hf == total_offset_19[6:0] ? phv_data_15 : _GEN_1147; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1149 = 7'h10 == total_offset_19[6:0] ? phv_data_16 : _GEN_1148; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1150 = 7'h11 == total_offset_19[6:0] ? phv_data_17 : _GEN_1149; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1151 = 7'h12 == total_offset_19[6:0] ? phv_data_18 : _GEN_1150; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1152 = 7'h13 == total_offset_19[6:0] ? phv_data_19 : _GEN_1151; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1153 = 7'h14 == total_offset_19[6:0] ? phv_data_20 : _GEN_1152; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1154 = 7'h15 == total_offset_19[6:0] ? phv_data_21 : _GEN_1153; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1155 = 7'h16 == total_offset_19[6:0] ? phv_data_22 : _GEN_1154; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1156 = 7'h17 == total_offset_19[6:0] ? phv_data_23 : _GEN_1155; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1157 = 7'h18 == total_offset_19[6:0] ? phv_data_24 : _GEN_1156; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1158 = 7'h19 == total_offset_19[6:0] ? phv_data_25 : _GEN_1157; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1159 = 7'h1a == total_offset_19[6:0] ? phv_data_26 : _GEN_1158; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1160 = 7'h1b == total_offset_19[6:0] ? phv_data_27 : _GEN_1159; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1161 = 7'h1c == total_offset_19[6:0] ? phv_data_28 : _GEN_1160; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1162 = 7'h1d == total_offset_19[6:0] ? phv_data_29 : _GEN_1161; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1163 = 7'h1e == total_offset_19[6:0] ? phv_data_30 : _GEN_1162; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1164 = 7'h1f == total_offset_19[6:0] ? phv_data_31 : _GEN_1163; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1165 = 7'h20 == total_offset_19[6:0] ? phv_data_32 : _GEN_1164; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1166 = 7'h21 == total_offset_19[6:0] ? phv_data_33 : _GEN_1165; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1167 = 7'h22 == total_offset_19[6:0] ? phv_data_34 : _GEN_1166; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1168 = 7'h23 == total_offset_19[6:0] ? phv_data_35 : _GEN_1167; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1169 = 7'h24 == total_offset_19[6:0] ? phv_data_36 : _GEN_1168; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1170 = 7'h25 == total_offset_19[6:0] ? phv_data_37 : _GEN_1169; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1171 = 7'h26 == total_offset_19[6:0] ? phv_data_38 : _GEN_1170; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1172 = 7'h27 == total_offset_19[6:0] ? phv_data_39 : _GEN_1171; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1173 = 7'h28 == total_offset_19[6:0] ? phv_data_40 : _GEN_1172; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1174 = 7'h29 == total_offset_19[6:0] ? phv_data_41 : _GEN_1173; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1175 = 7'h2a == total_offset_19[6:0] ? phv_data_42 : _GEN_1174; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1176 = 7'h2b == total_offset_19[6:0] ? phv_data_43 : _GEN_1175; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1177 = 7'h2c == total_offset_19[6:0] ? phv_data_44 : _GEN_1176; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1178 = 7'h2d == total_offset_19[6:0] ? phv_data_45 : _GEN_1177; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1179 = 7'h2e == total_offset_19[6:0] ? phv_data_46 : _GEN_1178; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1180 = 7'h2f == total_offset_19[6:0] ? phv_data_47 : _GEN_1179; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1181 = 7'h30 == total_offset_19[6:0] ? phv_data_48 : _GEN_1180; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1182 = 7'h31 == total_offset_19[6:0] ? phv_data_49 : _GEN_1181; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1183 = 7'h32 == total_offset_19[6:0] ? phv_data_50 : _GEN_1182; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1184 = 7'h33 == total_offset_19[6:0] ? phv_data_51 : _GEN_1183; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1185 = 7'h34 == total_offset_19[6:0] ? phv_data_52 : _GEN_1184; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1186 = 7'h35 == total_offset_19[6:0] ? phv_data_53 : _GEN_1185; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1187 = 7'h36 == total_offset_19[6:0] ? phv_data_54 : _GEN_1186; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1188 = 7'h37 == total_offset_19[6:0] ? phv_data_55 : _GEN_1187; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1189 = 7'h38 == total_offset_19[6:0] ? phv_data_56 : _GEN_1188; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1190 = 7'h39 == total_offset_19[6:0] ? phv_data_57 : _GEN_1189; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1191 = 7'h3a == total_offset_19[6:0] ? phv_data_58 : _GEN_1190; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1192 = 7'h3b == total_offset_19[6:0] ? phv_data_59 : _GEN_1191; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1193 = 7'h3c == total_offset_19[6:0] ? phv_data_60 : _GEN_1192; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1194 = 7'h3d == total_offset_19[6:0] ? phv_data_61 : _GEN_1193; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1195 = 7'h3e == total_offset_19[6:0] ? phv_data_62 : _GEN_1194; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1196 = 7'h3f == total_offset_19[6:0] ? phv_data_63 : _GEN_1195; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1197 = 7'h40 == total_offset_19[6:0] ? phv_data_64 : _GEN_1196; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1198 = 7'h41 == total_offset_19[6:0] ? phv_data_65 : _GEN_1197; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1199 = 7'h42 == total_offset_19[6:0] ? phv_data_66 : _GEN_1198; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1200 = 7'h43 == total_offset_19[6:0] ? phv_data_67 : _GEN_1199; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1201 = 7'h44 == total_offset_19[6:0] ? phv_data_68 : _GEN_1200; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1202 = 7'h45 == total_offset_19[6:0] ? phv_data_69 : _GEN_1201; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1203 = 7'h46 == total_offset_19[6:0] ? phv_data_70 : _GEN_1202; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1204 = 7'h47 == total_offset_19[6:0] ? phv_data_71 : _GEN_1203; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1205 = 7'h48 == total_offset_19[6:0] ? phv_data_72 : _GEN_1204; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1206 = 7'h49 == total_offset_19[6:0] ? phv_data_73 : _GEN_1205; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1207 = 7'h4a == total_offset_19[6:0] ? phv_data_74 : _GEN_1206; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1208 = 7'h4b == total_offset_19[6:0] ? phv_data_75 : _GEN_1207; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1209 = 7'h4c == total_offset_19[6:0] ? phv_data_76 : _GEN_1208; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1210 = 7'h4d == total_offset_19[6:0] ? phv_data_77 : _GEN_1209; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1211 = 7'h4e == total_offset_19[6:0] ? phv_data_78 : _GEN_1210; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1212 = 7'h4f == total_offset_19[6:0] ? phv_data_79 : _GEN_1211; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1213 = 7'h50 == total_offset_19[6:0] ? phv_data_80 : _GEN_1212; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1214 = 7'h51 == total_offset_19[6:0] ? phv_data_81 : _GEN_1213; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1215 = 7'h52 == total_offset_19[6:0] ? phv_data_82 : _GEN_1214; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1216 = 7'h53 == total_offset_19[6:0] ? phv_data_83 : _GEN_1215; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1217 = 7'h54 == total_offset_19[6:0] ? phv_data_84 : _GEN_1216; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1218 = 7'h55 == total_offset_19[6:0] ? phv_data_85 : _GEN_1217; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1219 = 7'h56 == total_offset_19[6:0] ? phv_data_86 : _GEN_1218; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1220 = 7'h57 == total_offset_19[6:0] ? phv_data_87 : _GEN_1219; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1221 = 7'h58 == total_offset_19[6:0] ? phv_data_88 : _GEN_1220; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1222 = 7'h59 == total_offset_19[6:0] ? phv_data_89 : _GEN_1221; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1223 = 7'h5a == total_offset_19[6:0] ? phv_data_90 : _GEN_1222; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1224 = 7'h5b == total_offset_19[6:0] ? phv_data_91 : _GEN_1223; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1225 = 7'h5c == total_offset_19[6:0] ? phv_data_92 : _GEN_1224; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1226 = 7'h5d == total_offset_19[6:0] ? phv_data_93 : _GEN_1225; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1227 = 7'h5e == total_offset_19[6:0] ? phv_data_94 : _GEN_1226; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1228 = 7'h5f == total_offset_19[6:0] ? phv_data_95 : _GEN_1227; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_3 = 8'h3 < length_1 ? _GEN_1228 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_20 = offset_1 + 8'h4; // @[executor.scala 148:53]
  wire [7:0] _GEN_1231 = 7'h1 == total_offset_20[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1232 = 7'h2 == total_offset_20[6:0] ? phv_data_2 : _GEN_1231; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1233 = 7'h3 == total_offset_20[6:0] ? phv_data_3 : _GEN_1232; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1234 = 7'h4 == total_offset_20[6:0] ? phv_data_4 : _GEN_1233; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1235 = 7'h5 == total_offset_20[6:0] ? phv_data_5 : _GEN_1234; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1236 = 7'h6 == total_offset_20[6:0] ? phv_data_6 : _GEN_1235; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1237 = 7'h7 == total_offset_20[6:0] ? phv_data_7 : _GEN_1236; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1238 = 7'h8 == total_offset_20[6:0] ? phv_data_8 : _GEN_1237; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1239 = 7'h9 == total_offset_20[6:0] ? phv_data_9 : _GEN_1238; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1240 = 7'ha == total_offset_20[6:0] ? phv_data_10 : _GEN_1239; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1241 = 7'hb == total_offset_20[6:0] ? phv_data_11 : _GEN_1240; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1242 = 7'hc == total_offset_20[6:0] ? phv_data_12 : _GEN_1241; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1243 = 7'hd == total_offset_20[6:0] ? phv_data_13 : _GEN_1242; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1244 = 7'he == total_offset_20[6:0] ? phv_data_14 : _GEN_1243; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1245 = 7'hf == total_offset_20[6:0] ? phv_data_15 : _GEN_1244; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1246 = 7'h10 == total_offset_20[6:0] ? phv_data_16 : _GEN_1245; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1247 = 7'h11 == total_offset_20[6:0] ? phv_data_17 : _GEN_1246; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1248 = 7'h12 == total_offset_20[6:0] ? phv_data_18 : _GEN_1247; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1249 = 7'h13 == total_offset_20[6:0] ? phv_data_19 : _GEN_1248; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1250 = 7'h14 == total_offset_20[6:0] ? phv_data_20 : _GEN_1249; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1251 = 7'h15 == total_offset_20[6:0] ? phv_data_21 : _GEN_1250; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1252 = 7'h16 == total_offset_20[6:0] ? phv_data_22 : _GEN_1251; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1253 = 7'h17 == total_offset_20[6:0] ? phv_data_23 : _GEN_1252; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1254 = 7'h18 == total_offset_20[6:0] ? phv_data_24 : _GEN_1253; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1255 = 7'h19 == total_offset_20[6:0] ? phv_data_25 : _GEN_1254; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1256 = 7'h1a == total_offset_20[6:0] ? phv_data_26 : _GEN_1255; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1257 = 7'h1b == total_offset_20[6:0] ? phv_data_27 : _GEN_1256; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1258 = 7'h1c == total_offset_20[6:0] ? phv_data_28 : _GEN_1257; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1259 = 7'h1d == total_offset_20[6:0] ? phv_data_29 : _GEN_1258; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1260 = 7'h1e == total_offset_20[6:0] ? phv_data_30 : _GEN_1259; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1261 = 7'h1f == total_offset_20[6:0] ? phv_data_31 : _GEN_1260; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1262 = 7'h20 == total_offset_20[6:0] ? phv_data_32 : _GEN_1261; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1263 = 7'h21 == total_offset_20[6:0] ? phv_data_33 : _GEN_1262; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1264 = 7'h22 == total_offset_20[6:0] ? phv_data_34 : _GEN_1263; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1265 = 7'h23 == total_offset_20[6:0] ? phv_data_35 : _GEN_1264; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1266 = 7'h24 == total_offset_20[6:0] ? phv_data_36 : _GEN_1265; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1267 = 7'h25 == total_offset_20[6:0] ? phv_data_37 : _GEN_1266; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1268 = 7'h26 == total_offset_20[6:0] ? phv_data_38 : _GEN_1267; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1269 = 7'h27 == total_offset_20[6:0] ? phv_data_39 : _GEN_1268; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1270 = 7'h28 == total_offset_20[6:0] ? phv_data_40 : _GEN_1269; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1271 = 7'h29 == total_offset_20[6:0] ? phv_data_41 : _GEN_1270; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1272 = 7'h2a == total_offset_20[6:0] ? phv_data_42 : _GEN_1271; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1273 = 7'h2b == total_offset_20[6:0] ? phv_data_43 : _GEN_1272; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1274 = 7'h2c == total_offset_20[6:0] ? phv_data_44 : _GEN_1273; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1275 = 7'h2d == total_offset_20[6:0] ? phv_data_45 : _GEN_1274; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1276 = 7'h2e == total_offset_20[6:0] ? phv_data_46 : _GEN_1275; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1277 = 7'h2f == total_offset_20[6:0] ? phv_data_47 : _GEN_1276; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1278 = 7'h30 == total_offset_20[6:0] ? phv_data_48 : _GEN_1277; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1279 = 7'h31 == total_offset_20[6:0] ? phv_data_49 : _GEN_1278; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1280 = 7'h32 == total_offset_20[6:0] ? phv_data_50 : _GEN_1279; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1281 = 7'h33 == total_offset_20[6:0] ? phv_data_51 : _GEN_1280; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1282 = 7'h34 == total_offset_20[6:0] ? phv_data_52 : _GEN_1281; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1283 = 7'h35 == total_offset_20[6:0] ? phv_data_53 : _GEN_1282; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1284 = 7'h36 == total_offset_20[6:0] ? phv_data_54 : _GEN_1283; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1285 = 7'h37 == total_offset_20[6:0] ? phv_data_55 : _GEN_1284; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1286 = 7'h38 == total_offset_20[6:0] ? phv_data_56 : _GEN_1285; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1287 = 7'h39 == total_offset_20[6:0] ? phv_data_57 : _GEN_1286; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1288 = 7'h3a == total_offset_20[6:0] ? phv_data_58 : _GEN_1287; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1289 = 7'h3b == total_offset_20[6:0] ? phv_data_59 : _GEN_1288; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1290 = 7'h3c == total_offset_20[6:0] ? phv_data_60 : _GEN_1289; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1291 = 7'h3d == total_offset_20[6:0] ? phv_data_61 : _GEN_1290; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1292 = 7'h3e == total_offset_20[6:0] ? phv_data_62 : _GEN_1291; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1293 = 7'h3f == total_offset_20[6:0] ? phv_data_63 : _GEN_1292; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1294 = 7'h40 == total_offset_20[6:0] ? phv_data_64 : _GEN_1293; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1295 = 7'h41 == total_offset_20[6:0] ? phv_data_65 : _GEN_1294; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1296 = 7'h42 == total_offset_20[6:0] ? phv_data_66 : _GEN_1295; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1297 = 7'h43 == total_offset_20[6:0] ? phv_data_67 : _GEN_1296; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1298 = 7'h44 == total_offset_20[6:0] ? phv_data_68 : _GEN_1297; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1299 = 7'h45 == total_offset_20[6:0] ? phv_data_69 : _GEN_1298; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1300 = 7'h46 == total_offset_20[6:0] ? phv_data_70 : _GEN_1299; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1301 = 7'h47 == total_offset_20[6:0] ? phv_data_71 : _GEN_1300; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1302 = 7'h48 == total_offset_20[6:0] ? phv_data_72 : _GEN_1301; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1303 = 7'h49 == total_offset_20[6:0] ? phv_data_73 : _GEN_1302; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1304 = 7'h4a == total_offset_20[6:0] ? phv_data_74 : _GEN_1303; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1305 = 7'h4b == total_offset_20[6:0] ? phv_data_75 : _GEN_1304; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1306 = 7'h4c == total_offset_20[6:0] ? phv_data_76 : _GEN_1305; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1307 = 7'h4d == total_offset_20[6:0] ? phv_data_77 : _GEN_1306; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1308 = 7'h4e == total_offset_20[6:0] ? phv_data_78 : _GEN_1307; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1309 = 7'h4f == total_offset_20[6:0] ? phv_data_79 : _GEN_1308; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1310 = 7'h50 == total_offset_20[6:0] ? phv_data_80 : _GEN_1309; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1311 = 7'h51 == total_offset_20[6:0] ? phv_data_81 : _GEN_1310; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1312 = 7'h52 == total_offset_20[6:0] ? phv_data_82 : _GEN_1311; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1313 = 7'h53 == total_offset_20[6:0] ? phv_data_83 : _GEN_1312; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1314 = 7'h54 == total_offset_20[6:0] ? phv_data_84 : _GEN_1313; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1315 = 7'h55 == total_offset_20[6:0] ? phv_data_85 : _GEN_1314; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1316 = 7'h56 == total_offset_20[6:0] ? phv_data_86 : _GEN_1315; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1317 = 7'h57 == total_offset_20[6:0] ? phv_data_87 : _GEN_1316; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1318 = 7'h58 == total_offset_20[6:0] ? phv_data_88 : _GEN_1317; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1319 = 7'h59 == total_offset_20[6:0] ? phv_data_89 : _GEN_1318; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1320 = 7'h5a == total_offset_20[6:0] ? phv_data_90 : _GEN_1319; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1321 = 7'h5b == total_offset_20[6:0] ? phv_data_91 : _GEN_1320; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1322 = 7'h5c == total_offset_20[6:0] ? phv_data_92 : _GEN_1321; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1323 = 7'h5d == total_offset_20[6:0] ? phv_data_93 : _GEN_1322; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1324 = 7'h5e == total_offset_20[6:0] ? phv_data_94 : _GEN_1323; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1325 = 7'h5f == total_offset_20[6:0] ? phv_data_95 : _GEN_1324; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_4 = 8'h4 < length_1 ? _GEN_1325 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_21 = offset_1 + 8'h5; // @[executor.scala 148:53]
  wire [7:0] _GEN_1328 = 7'h1 == total_offset_21[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1329 = 7'h2 == total_offset_21[6:0] ? phv_data_2 : _GEN_1328; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1330 = 7'h3 == total_offset_21[6:0] ? phv_data_3 : _GEN_1329; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1331 = 7'h4 == total_offset_21[6:0] ? phv_data_4 : _GEN_1330; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1332 = 7'h5 == total_offset_21[6:0] ? phv_data_5 : _GEN_1331; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1333 = 7'h6 == total_offset_21[6:0] ? phv_data_6 : _GEN_1332; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1334 = 7'h7 == total_offset_21[6:0] ? phv_data_7 : _GEN_1333; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1335 = 7'h8 == total_offset_21[6:0] ? phv_data_8 : _GEN_1334; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1336 = 7'h9 == total_offset_21[6:0] ? phv_data_9 : _GEN_1335; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1337 = 7'ha == total_offset_21[6:0] ? phv_data_10 : _GEN_1336; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1338 = 7'hb == total_offset_21[6:0] ? phv_data_11 : _GEN_1337; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1339 = 7'hc == total_offset_21[6:0] ? phv_data_12 : _GEN_1338; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1340 = 7'hd == total_offset_21[6:0] ? phv_data_13 : _GEN_1339; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1341 = 7'he == total_offset_21[6:0] ? phv_data_14 : _GEN_1340; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1342 = 7'hf == total_offset_21[6:0] ? phv_data_15 : _GEN_1341; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1343 = 7'h10 == total_offset_21[6:0] ? phv_data_16 : _GEN_1342; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1344 = 7'h11 == total_offset_21[6:0] ? phv_data_17 : _GEN_1343; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1345 = 7'h12 == total_offset_21[6:0] ? phv_data_18 : _GEN_1344; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1346 = 7'h13 == total_offset_21[6:0] ? phv_data_19 : _GEN_1345; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1347 = 7'h14 == total_offset_21[6:0] ? phv_data_20 : _GEN_1346; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1348 = 7'h15 == total_offset_21[6:0] ? phv_data_21 : _GEN_1347; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1349 = 7'h16 == total_offset_21[6:0] ? phv_data_22 : _GEN_1348; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1350 = 7'h17 == total_offset_21[6:0] ? phv_data_23 : _GEN_1349; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1351 = 7'h18 == total_offset_21[6:0] ? phv_data_24 : _GEN_1350; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1352 = 7'h19 == total_offset_21[6:0] ? phv_data_25 : _GEN_1351; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1353 = 7'h1a == total_offset_21[6:0] ? phv_data_26 : _GEN_1352; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1354 = 7'h1b == total_offset_21[6:0] ? phv_data_27 : _GEN_1353; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1355 = 7'h1c == total_offset_21[6:0] ? phv_data_28 : _GEN_1354; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1356 = 7'h1d == total_offset_21[6:0] ? phv_data_29 : _GEN_1355; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1357 = 7'h1e == total_offset_21[6:0] ? phv_data_30 : _GEN_1356; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1358 = 7'h1f == total_offset_21[6:0] ? phv_data_31 : _GEN_1357; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1359 = 7'h20 == total_offset_21[6:0] ? phv_data_32 : _GEN_1358; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1360 = 7'h21 == total_offset_21[6:0] ? phv_data_33 : _GEN_1359; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1361 = 7'h22 == total_offset_21[6:0] ? phv_data_34 : _GEN_1360; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1362 = 7'h23 == total_offset_21[6:0] ? phv_data_35 : _GEN_1361; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1363 = 7'h24 == total_offset_21[6:0] ? phv_data_36 : _GEN_1362; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1364 = 7'h25 == total_offset_21[6:0] ? phv_data_37 : _GEN_1363; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1365 = 7'h26 == total_offset_21[6:0] ? phv_data_38 : _GEN_1364; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1366 = 7'h27 == total_offset_21[6:0] ? phv_data_39 : _GEN_1365; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1367 = 7'h28 == total_offset_21[6:0] ? phv_data_40 : _GEN_1366; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1368 = 7'h29 == total_offset_21[6:0] ? phv_data_41 : _GEN_1367; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1369 = 7'h2a == total_offset_21[6:0] ? phv_data_42 : _GEN_1368; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1370 = 7'h2b == total_offset_21[6:0] ? phv_data_43 : _GEN_1369; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1371 = 7'h2c == total_offset_21[6:0] ? phv_data_44 : _GEN_1370; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1372 = 7'h2d == total_offset_21[6:0] ? phv_data_45 : _GEN_1371; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1373 = 7'h2e == total_offset_21[6:0] ? phv_data_46 : _GEN_1372; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1374 = 7'h2f == total_offset_21[6:0] ? phv_data_47 : _GEN_1373; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1375 = 7'h30 == total_offset_21[6:0] ? phv_data_48 : _GEN_1374; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1376 = 7'h31 == total_offset_21[6:0] ? phv_data_49 : _GEN_1375; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1377 = 7'h32 == total_offset_21[6:0] ? phv_data_50 : _GEN_1376; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1378 = 7'h33 == total_offset_21[6:0] ? phv_data_51 : _GEN_1377; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1379 = 7'h34 == total_offset_21[6:0] ? phv_data_52 : _GEN_1378; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1380 = 7'h35 == total_offset_21[6:0] ? phv_data_53 : _GEN_1379; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1381 = 7'h36 == total_offset_21[6:0] ? phv_data_54 : _GEN_1380; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1382 = 7'h37 == total_offset_21[6:0] ? phv_data_55 : _GEN_1381; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1383 = 7'h38 == total_offset_21[6:0] ? phv_data_56 : _GEN_1382; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1384 = 7'h39 == total_offset_21[6:0] ? phv_data_57 : _GEN_1383; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1385 = 7'h3a == total_offset_21[6:0] ? phv_data_58 : _GEN_1384; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1386 = 7'h3b == total_offset_21[6:0] ? phv_data_59 : _GEN_1385; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1387 = 7'h3c == total_offset_21[6:0] ? phv_data_60 : _GEN_1386; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1388 = 7'h3d == total_offset_21[6:0] ? phv_data_61 : _GEN_1387; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1389 = 7'h3e == total_offset_21[6:0] ? phv_data_62 : _GEN_1388; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1390 = 7'h3f == total_offset_21[6:0] ? phv_data_63 : _GEN_1389; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1391 = 7'h40 == total_offset_21[6:0] ? phv_data_64 : _GEN_1390; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1392 = 7'h41 == total_offset_21[6:0] ? phv_data_65 : _GEN_1391; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1393 = 7'h42 == total_offset_21[6:0] ? phv_data_66 : _GEN_1392; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1394 = 7'h43 == total_offset_21[6:0] ? phv_data_67 : _GEN_1393; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1395 = 7'h44 == total_offset_21[6:0] ? phv_data_68 : _GEN_1394; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1396 = 7'h45 == total_offset_21[6:0] ? phv_data_69 : _GEN_1395; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1397 = 7'h46 == total_offset_21[6:0] ? phv_data_70 : _GEN_1396; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1398 = 7'h47 == total_offset_21[6:0] ? phv_data_71 : _GEN_1397; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1399 = 7'h48 == total_offset_21[6:0] ? phv_data_72 : _GEN_1398; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1400 = 7'h49 == total_offset_21[6:0] ? phv_data_73 : _GEN_1399; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1401 = 7'h4a == total_offset_21[6:0] ? phv_data_74 : _GEN_1400; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1402 = 7'h4b == total_offset_21[6:0] ? phv_data_75 : _GEN_1401; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1403 = 7'h4c == total_offset_21[6:0] ? phv_data_76 : _GEN_1402; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1404 = 7'h4d == total_offset_21[6:0] ? phv_data_77 : _GEN_1403; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1405 = 7'h4e == total_offset_21[6:0] ? phv_data_78 : _GEN_1404; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1406 = 7'h4f == total_offset_21[6:0] ? phv_data_79 : _GEN_1405; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1407 = 7'h50 == total_offset_21[6:0] ? phv_data_80 : _GEN_1406; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1408 = 7'h51 == total_offset_21[6:0] ? phv_data_81 : _GEN_1407; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1409 = 7'h52 == total_offset_21[6:0] ? phv_data_82 : _GEN_1408; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1410 = 7'h53 == total_offset_21[6:0] ? phv_data_83 : _GEN_1409; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1411 = 7'h54 == total_offset_21[6:0] ? phv_data_84 : _GEN_1410; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1412 = 7'h55 == total_offset_21[6:0] ? phv_data_85 : _GEN_1411; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1413 = 7'h56 == total_offset_21[6:0] ? phv_data_86 : _GEN_1412; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1414 = 7'h57 == total_offset_21[6:0] ? phv_data_87 : _GEN_1413; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1415 = 7'h58 == total_offset_21[6:0] ? phv_data_88 : _GEN_1414; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1416 = 7'h59 == total_offset_21[6:0] ? phv_data_89 : _GEN_1415; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1417 = 7'h5a == total_offset_21[6:0] ? phv_data_90 : _GEN_1416; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1418 = 7'h5b == total_offset_21[6:0] ? phv_data_91 : _GEN_1417; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1419 = 7'h5c == total_offset_21[6:0] ? phv_data_92 : _GEN_1418; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1420 = 7'h5d == total_offset_21[6:0] ? phv_data_93 : _GEN_1419; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1421 = 7'h5e == total_offset_21[6:0] ? phv_data_94 : _GEN_1420; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1422 = 7'h5f == total_offset_21[6:0] ? phv_data_95 : _GEN_1421; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_5 = 8'h5 < length_1 ? _GEN_1422 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_22 = offset_1 + 8'h6; // @[executor.scala 148:53]
  wire [7:0] _GEN_1425 = 7'h1 == total_offset_22[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1426 = 7'h2 == total_offset_22[6:0] ? phv_data_2 : _GEN_1425; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1427 = 7'h3 == total_offset_22[6:0] ? phv_data_3 : _GEN_1426; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1428 = 7'h4 == total_offset_22[6:0] ? phv_data_4 : _GEN_1427; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1429 = 7'h5 == total_offset_22[6:0] ? phv_data_5 : _GEN_1428; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1430 = 7'h6 == total_offset_22[6:0] ? phv_data_6 : _GEN_1429; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1431 = 7'h7 == total_offset_22[6:0] ? phv_data_7 : _GEN_1430; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1432 = 7'h8 == total_offset_22[6:0] ? phv_data_8 : _GEN_1431; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1433 = 7'h9 == total_offset_22[6:0] ? phv_data_9 : _GEN_1432; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1434 = 7'ha == total_offset_22[6:0] ? phv_data_10 : _GEN_1433; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1435 = 7'hb == total_offset_22[6:0] ? phv_data_11 : _GEN_1434; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1436 = 7'hc == total_offset_22[6:0] ? phv_data_12 : _GEN_1435; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1437 = 7'hd == total_offset_22[6:0] ? phv_data_13 : _GEN_1436; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1438 = 7'he == total_offset_22[6:0] ? phv_data_14 : _GEN_1437; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1439 = 7'hf == total_offset_22[6:0] ? phv_data_15 : _GEN_1438; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1440 = 7'h10 == total_offset_22[6:0] ? phv_data_16 : _GEN_1439; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1441 = 7'h11 == total_offset_22[6:0] ? phv_data_17 : _GEN_1440; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1442 = 7'h12 == total_offset_22[6:0] ? phv_data_18 : _GEN_1441; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1443 = 7'h13 == total_offset_22[6:0] ? phv_data_19 : _GEN_1442; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1444 = 7'h14 == total_offset_22[6:0] ? phv_data_20 : _GEN_1443; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1445 = 7'h15 == total_offset_22[6:0] ? phv_data_21 : _GEN_1444; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1446 = 7'h16 == total_offset_22[6:0] ? phv_data_22 : _GEN_1445; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1447 = 7'h17 == total_offset_22[6:0] ? phv_data_23 : _GEN_1446; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1448 = 7'h18 == total_offset_22[6:0] ? phv_data_24 : _GEN_1447; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1449 = 7'h19 == total_offset_22[6:0] ? phv_data_25 : _GEN_1448; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1450 = 7'h1a == total_offset_22[6:0] ? phv_data_26 : _GEN_1449; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1451 = 7'h1b == total_offset_22[6:0] ? phv_data_27 : _GEN_1450; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1452 = 7'h1c == total_offset_22[6:0] ? phv_data_28 : _GEN_1451; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1453 = 7'h1d == total_offset_22[6:0] ? phv_data_29 : _GEN_1452; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1454 = 7'h1e == total_offset_22[6:0] ? phv_data_30 : _GEN_1453; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1455 = 7'h1f == total_offset_22[6:0] ? phv_data_31 : _GEN_1454; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1456 = 7'h20 == total_offset_22[6:0] ? phv_data_32 : _GEN_1455; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1457 = 7'h21 == total_offset_22[6:0] ? phv_data_33 : _GEN_1456; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1458 = 7'h22 == total_offset_22[6:0] ? phv_data_34 : _GEN_1457; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1459 = 7'h23 == total_offset_22[6:0] ? phv_data_35 : _GEN_1458; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1460 = 7'h24 == total_offset_22[6:0] ? phv_data_36 : _GEN_1459; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1461 = 7'h25 == total_offset_22[6:0] ? phv_data_37 : _GEN_1460; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1462 = 7'h26 == total_offset_22[6:0] ? phv_data_38 : _GEN_1461; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1463 = 7'h27 == total_offset_22[6:0] ? phv_data_39 : _GEN_1462; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1464 = 7'h28 == total_offset_22[6:0] ? phv_data_40 : _GEN_1463; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1465 = 7'h29 == total_offset_22[6:0] ? phv_data_41 : _GEN_1464; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1466 = 7'h2a == total_offset_22[6:0] ? phv_data_42 : _GEN_1465; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1467 = 7'h2b == total_offset_22[6:0] ? phv_data_43 : _GEN_1466; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1468 = 7'h2c == total_offset_22[6:0] ? phv_data_44 : _GEN_1467; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1469 = 7'h2d == total_offset_22[6:0] ? phv_data_45 : _GEN_1468; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1470 = 7'h2e == total_offset_22[6:0] ? phv_data_46 : _GEN_1469; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1471 = 7'h2f == total_offset_22[6:0] ? phv_data_47 : _GEN_1470; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1472 = 7'h30 == total_offset_22[6:0] ? phv_data_48 : _GEN_1471; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1473 = 7'h31 == total_offset_22[6:0] ? phv_data_49 : _GEN_1472; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1474 = 7'h32 == total_offset_22[6:0] ? phv_data_50 : _GEN_1473; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1475 = 7'h33 == total_offset_22[6:0] ? phv_data_51 : _GEN_1474; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1476 = 7'h34 == total_offset_22[6:0] ? phv_data_52 : _GEN_1475; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1477 = 7'h35 == total_offset_22[6:0] ? phv_data_53 : _GEN_1476; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1478 = 7'h36 == total_offset_22[6:0] ? phv_data_54 : _GEN_1477; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1479 = 7'h37 == total_offset_22[6:0] ? phv_data_55 : _GEN_1478; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1480 = 7'h38 == total_offset_22[6:0] ? phv_data_56 : _GEN_1479; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1481 = 7'h39 == total_offset_22[6:0] ? phv_data_57 : _GEN_1480; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1482 = 7'h3a == total_offset_22[6:0] ? phv_data_58 : _GEN_1481; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1483 = 7'h3b == total_offset_22[6:0] ? phv_data_59 : _GEN_1482; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1484 = 7'h3c == total_offset_22[6:0] ? phv_data_60 : _GEN_1483; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1485 = 7'h3d == total_offset_22[6:0] ? phv_data_61 : _GEN_1484; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1486 = 7'h3e == total_offset_22[6:0] ? phv_data_62 : _GEN_1485; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1487 = 7'h3f == total_offset_22[6:0] ? phv_data_63 : _GEN_1486; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1488 = 7'h40 == total_offset_22[6:0] ? phv_data_64 : _GEN_1487; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1489 = 7'h41 == total_offset_22[6:0] ? phv_data_65 : _GEN_1488; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1490 = 7'h42 == total_offset_22[6:0] ? phv_data_66 : _GEN_1489; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1491 = 7'h43 == total_offset_22[6:0] ? phv_data_67 : _GEN_1490; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1492 = 7'h44 == total_offset_22[6:0] ? phv_data_68 : _GEN_1491; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1493 = 7'h45 == total_offset_22[6:0] ? phv_data_69 : _GEN_1492; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1494 = 7'h46 == total_offset_22[6:0] ? phv_data_70 : _GEN_1493; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1495 = 7'h47 == total_offset_22[6:0] ? phv_data_71 : _GEN_1494; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1496 = 7'h48 == total_offset_22[6:0] ? phv_data_72 : _GEN_1495; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1497 = 7'h49 == total_offset_22[6:0] ? phv_data_73 : _GEN_1496; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1498 = 7'h4a == total_offset_22[6:0] ? phv_data_74 : _GEN_1497; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1499 = 7'h4b == total_offset_22[6:0] ? phv_data_75 : _GEN_1498; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1500 = 7'h4c == total_offset_22[6:0] ? phv_data_76 : _GEN_1499; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1501 = 7'h4d == total_offset_22[6:0] ? phv_data_77 : _GEN_1500; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1502 = 7'h4e == total_offset_22[6:0] ? phv_data_78 : _GEN_1501; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1503 = 7'h4f == total_offset_22[6:0] ? phv_data_79 : _GEN_1502; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1504 = 7'h50 == total_offset_22[6:0] ? phv_data_80 : _GEN_1503; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1505 = 7'h51 == total_offset_22[6:0] ? phv_data_81 : _GEN_1504; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1506 = 7'h52 == total_offset_22[6:0] ? phv_data_82 : _GEN_1505; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1507 = 7'h53 == total_offset_22[6:0] ? phv_data_83 : _GEN_1506; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1508 = 7'h54 == total_offset_22[6:0] ? phv_data_84 : _GEN_1507; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1509 = 7'h55 == total_offset_22[6:0] ? phv_data_85 : _GEN_1508; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1510 = 7'h56 == total_offset_22[6:0] ? phv_data_86 : _GEN_1509; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1511 = 7'h57 == total_offset_22[6:0] ? phv_data_87 : _GEN_1510; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1512 = 7'h58 == total_offset_22[6:0] ? phv_data_88 : _GEN_1511; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1513 = 7'h59 == total_offset_22[6:0] ? phv_data_89 : _GEN_1512; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1514 = 7'h5a == total_offset_22[6:0] ? phv_data_90 : _GEN_1513; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1515 = 7'h5b == total_offset_22[6:0] ? phv_data_91 : _GEN_1514; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1516 = 7'h5c == total_offset_22[6:0] ? phv_data_92 : _GEN_1515; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1517 = 7'h5d == total_offset_22[6:0] ? phv_data_93 : _GEN_1516; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1518 = 7'h5e == total_offset_22[6:0] ? phv_data_94 : _GEN_1517; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1519 = 7'h5f == total_offset_22[6:0] ? phv_data_95 : _GEN_1518; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_6 = 8'h6 < length_1 ? _GEN_1519 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_23 = offset_1 + 8'h7; // @[executor.scala 148:53]
  wire [7:0] _GEN_1522 = 7'h1 == total_offset_23[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1523 = 7'h2 == total_offset_23[6:0] ? phv_data_2 : _GEN_1522; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1524 = 7'h3 == total_offset_23[6:0] ? phv_data_3 : _GEN_1523; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1525 = 7'h4 == total_offset_23[6:0] ? phv_data_4 : _GEN_1524; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1526 = 7'h5 == total_offset_23[6:0] ? phv_data_5 : _GEN_1525; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1527 = 7'h6 == total_offset_23[6:0] ? phv_data_6 : _GEN_1526; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1528 = 7'h7 == total_offset_23[6:0] ? phv_data_7 : _GEN_1527; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1529 = 7'h8 == total_offset_23[6:0] ? phv_data_8 : _GEN_1528; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1530 = 7'h9 == total_offset_23[6:0] ? phv_data_9 : _GEN_1529; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1531 = 7'ha == total_offset_23[6:0] ? phv_data_10 : _GEN_1530; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1532 = 7'hb == total_offset_23[6:0] ? phv_data_11 : _GEN_1531; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1533 = 7'hc == total_offset_23[6:0] ? phv_data_12 : _GEN_1532; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1534 = 7'hd == total_offset_23[6:0] ? phv_data_13 : _GEN_1533; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1535 = 7'he == total_offset_23[6:0] ? phv_data_14 : _GEN_1534; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1536 = 7'hf == total_offset_23[6:0] ? phv_data_15 : _GEN_1535; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1537 = 7'h10 == total_offset_23[6:0] ? phv_data_16 : _GEN_1536; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1538 = 7'h11 == total_offset_23[6:0] ? phv_data_17 : _GEN_1537; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1539 = 7'h12 == total_offset_23[6:0] ? phv_data_18 : _GEN_1538; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1540 = 7'h13 == total_offset_23[6:0] ? phv_data_19 : _GEN_1539; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1541 = 7'h14 == total_offset_23[6:0] ? phv_data_20 : _GEN_1540; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1542 = 7'h15 == total_offset_23[6:0] ? phv_data_21 : _GEN_1541; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1543 = 7'h16 == total_offset_23[6:0] ? phv_data_22 : _GEN_1542; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1544 = 7'h17 == total_offset_23[6:0] ? phv_data_23 : _GEN_1543; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1545 = 7'h18 == total_offset_23[6:0] ? phv_data_24 : _GEN_1544; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1546 = 7'h19 == total_offset_23[6:0] ? phv_data_25 : _GEN_1545; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1547 = 7'h1a == total_offset_23[6:0] ? phv_data_26 : _GEN_1546; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1548 = 7'h1b == total_offset_23[6:0] ? phv_data_27 : _GEN_1547; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1549 = 7'h1c == total_offset_23[6:0] ? phv_data_28 : _GEN_1548; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1550 = 7'h1d == total_offset_23[6:0] ? phv_data_29 : _GEN_1549; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1551 = 7'h1e == total_offset_23[6:0] ? phv_data_30 : _GEN_1550; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1552 = 7'h1f == total_offset_23[6:0] ? phv_data_31 : _GEN_1551; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1553 = 7'h20 == total_offset_23[6:0] ? phv_data_32 : _GEN_1552; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1554 = 7'h21 == total_offset_23[6:0] ? phv_data_33 : _GEN_1553; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1555 = 7'h22 == total_offset_23[6:0] ? phv_data_34 : _GEN_1554; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1556 = 7'h23 == total_offset_23[6:0] ? phv_data_35 : _GEN_1555; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1557 = 7'h24 == total_offset_23[6:0] ? phv_data_36 : _GEN_1556; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1558 = 7'h25 == total_offset_23[6:0] ? phv_data_37 : _GEN_1557; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1559 = 7'h26 == total_offset_23[6:0] ? phv_data_38 : _GEN_1558; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1560 = 7'h27 == total_offset_23[6:0] ? phv_data_39 : _GEN_1559; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1561 = 7'h28 == total_offset_23[6:0] ? phv_data_40 : _GEN_1560; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1562 = 7'h29 == total_offset_23[6:0] ? phv_data_41 : _GEN_1561; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1563 = 7'h2a == total_offset_23[6:0] ? phv_data_42 : _GEN_1562; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1564 = 7'h2b == total_offset_23[6:0] ? phv_data_43 : _GEN_1563; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1565 = 7'h2c == total_offset_23[6:0] ? phv_data_44 : _GEN_1564; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1566 = 7'h2d == total_offset_23[6:0] ? phv_data_45 : _GEN_1565; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1567 = 7'h2e == total_offset_23[6:0] ? phv_data_46 : _GEN_1566; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1568 = 7'h2f == total_offset_23[6:0] ? phv_data_47 : _GEN_1567; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1569 = 7'h30 == total_offset_23[6:0] ? phv_data_48 : _GEN_1568; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1570 = 7'h31 == total_offset_23[6:0] ? phv_data_49 : _GEN_1569; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1571 = 7'h32 == total_offset_23[6:0] ? phv_data_50 : _GEN_1570; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1572 = 7'h33 == total_offset_23[6:0] ? phv_data_51 : _GEN_1571; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1573 = 7'h34 == total_offset_23[6:0] ? phv_data_52 : _GEN_1572; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1574 = 7'h35 == total_offset_23[6:0] ? phv_data_53 : _GEN_1573; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1575 = 7'h36 == total_offset_23[6:0] ? phv_data_54 : _GEN_1574; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1576 = 7'h37 == total_offset_23[6:0] ? phv_data_55 : _GEN_1575; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1577 = 7'h38 == total_offset_23[6:0] ? phv_data_56 : _GEN_1576; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1578 = 7'h39 == total_offset_23[6:0] ? phv_data_57 : _GEN_1577; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1579 = 7'h3a == total_offset_23[6:0] ? phv_data_58 : _GEN_1578; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1580 = 7'h3b == total_offset_23[6:0] ? phv_data_59 : _GEN_1579; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1581 = 7'h3c == total_offset_23[6:0] ? phv_data_60 : _GEN_1580; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1582 = 7'h3d == total_offset_23[6:0] ? phv_data_61 : _GEN_1581; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1583 = 7'h3e == total_offset_23[6:0] ? phv_data_62 : _GEN_1582; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1584 = 7'h3f == total_offset_23[6:0] ? phv_data_63 : _GEN_1583; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1585 = 7'h40 == total_offset_23[6:0] ? phv_data_64 : _GEN_1584; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1586 = 7'h41 == total_offset_23[6:0] ? phv_data_65 : _GEN_1585; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1587 = 7'h42 == total_offset_23[6:0] ? phv_data_66 : _GEN_1586; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1588 = 7'h43 == total_offset_23[6:0] ? phv_data_67 : _GEN_1587; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1589 = 7'h44 == total_offset_23[6:0] ? phv_data_68 : _GEN_1588; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1590 = 7'h45 == total_offset_23[6:0] ? phv_data_69 : _GEN_1589; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1591 = 7'h46 == total_offset_23[6:0] ? phv_data_70 : _GEN_1590; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1592 = 7'h47 == total_offset_23[6:0] ? phv_data_71 : _GEN_1591; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1593 = 7'h48 == total_offset_23[6:0] ? phv_data_72 : _GEN_1592; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1594 = 7'h49 == total_offset_23[6:0] ? phv_data_73 : _GEN_1593; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1595 = 7'h4a == total_offset_23[6:0] ? phv_data_74 : _GEN_1594; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1596 = 7'h4b == total_offset_23[6:0] ? phv_data_75 : _GEN_1595; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1597 = 7'h4c == total_offset_23[6:0] ? phv_data_76 : _GEN_1596; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1598 = 7'h4d == total_offset_23[6:0] ? phv_data_77 : _GEN_1597; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1599 = 7'h4e == total_offset_23[6:0] ? phv_data_78 : _GEN_1598; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1600 = 7'h4f == total_offset_23[6:0] ? phv_data_79 : _GEN_1599; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1601 = 7'h50 == total_offset_23[6:0] ? phv_data_80 : _GEN_1600; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1602 = 7'h51 == total_offset_23[6:0] ? phv_data_81 : _GEN_1601; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1603 = 7'h52 == total_offset_23[6:0] ? phv_data_82 : _GEN_1602; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1604 = 7'h53 == total_offset_23[6:0] ? phv_data_83 : _GEN_1603; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1605 = 7'h54 == total_offset_23[6:0] ? phv_data_84 : _GEN_1604; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1606 = 7'h55 == total_offset_23[6:0] ? phv_data_85 : _GEN_1605; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1607 = 7'h56 == total_offset_23[6:0] ? phv_data_86 : _GEN_1606; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1608 = 7'h57 == total_offset_23[6:0] ? phv_data_87 : _GEN_1607; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1609 = 7'h58 == total_offset_23[6:0] ? phv_data_88 : _GEN_1608; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1610 = 7'h59 == total_offset_23[6:0] ? phv_data_89 : _GEN_1609; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1611 = 7'h5a == total_offset_23[6:0] ? phv_data_90 : _GEN_1610; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1612 = 7'h5b == total_offset_23[6:0] ? phv_data_91 : _GEN_1611; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1613 = 7'h5c == total_offset_23[6:0] ? phv_data_92 : _GEN_1612; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1614 = 7'h5d == total_offset_23[6:0] ? phv_data_93 : _GEN_1613; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1615 = 7'h5e == total_offset_23[6:0] ? phv_data_94 : _GEN_1614; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1616 = 7'h5f == total_offset_23[6:0] ? phv_data_95 : _GEN_1615; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_2_7 = 8'h7 < length_1 ? _GEN_1616 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [63:0] _io_field_out_1_T = {bytes_2_0,bytes_2_1,bytes_2_2,bytes_2_3,bytes_2_4,bytes_2_5,bytes_2_6,bytes_2_7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_1 = io_field_out_1_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length_1 = io_field_out_1_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_24 = {{6'd0}, args_offset_1}; // @[executor.scala 163:56]
  wire [7:0] total_offset_24 = _total_offset_T_24[7:0]; // @[executor.scala 163:56]
  wire [7:0] _GEN_3382 = {{5'd0}, args_length_1}; // @[executor.scala 164:44]
  wire [7:0] _GEN_1619 = 3'h1 == total_offset_24[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1620 = 3'h2 == total_offset_24[2:0] ? args_2 : _GEN_1619; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1621 = 3'h3 == total_offset_24[2:0] ? args_3 : _GEN_1620; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1622 = 3'h4 == total_offset_24[2:0] ? args_4 : _GEN_1621; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1623 = 3'h5 == total_offset_24[2:0] ? args_5 : _GEN_1622; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1624 = 3'h6 == total_offset_24[2:0] ? args_6 : _GEN_1623; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_3_0 = 8'h0 < _GEN_3382 ? _GEN_1624 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] _GEN_3383 = {{5'd0}, args_offset_1}; // @[executor.scala 163:56]
  wire [7:0] total_offset_25 = _GEN_3383 + 8'h1; // @[executor.scala 163:56]
  wire [7:0] _GEN_1627 = 3'h1 == total_offset_25[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1628 = 3'h2 == total_offset_25[2:0] ? args_2 : _GEN_1627; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1629 = 3'h3 == total_offset_25[2:0] ? args_3 : _GEN_1628; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1630 = 3'h4 == total_offset_25[2:0] ? args_4 : _GEN_1629; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1631 = 3'h5 == total_offset_25[2:0] ? args_5 : _GEN_1630; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1632 = 3'h6 == total_offset_25[2:0] ? args_6 : _GEN_1631; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_3_1 = 8'h1 < _GEN_3382 ? _GEN_1632 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_26 = _GEN_3383 + 8'h2; // @[executor.scala 163:56]
  wire [7:0] _GEN_1635 = 3'h1 == total_offset_26[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1636 = 3'h2 == total_offset_26[2:0] ? args_2 : _GEN_1635; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1637 = 3'h3 == total_offset_26[2:0] ? args_3 : _GEN_1636; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1638 = 3'h4 == total_offset_26[2:0] ? args_4 : _GEN_1637; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1639 = 3'h5 == total_offset_26[2:0] ? args_5 : _GEN_1638; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1640 = 3'h6 == total_offset_26[2:0] ? args_6 : _GEN_1639; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_3_2 = 8'h2 < _GEN_3382 ? _GEN_1640 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_27 = _GEN_3383 + 8'h3; // @[executor.scala 163:56]
  wire [7:0] _GEN_1643 = 3'h1 == total_offset_27[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1644 = 3'h2 == total_offset_27[2:0] ? args_2 : _GEN_1643; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1645 = 3'h3 == total_offset_27[2:0] ? args_3 : _GEN_1644; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1646 = 3'h4 == total_offset_27[2:0] ? args_4 : _GEN_1645; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1647 = 3'h5 == total_offset_27[2:0] ? args_5 : _GEN_1646; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1648 = 3'h6 == total_offset_27[2:0] ? args_6 : _GEN_1647; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_3_3 = 8'h3 < _GEN_3382 ? _GEN_1648 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_28 = _GEN_3383 + 8'h4; // @[executor.scala 163:56]
  wire [7:0] _GEN_1651 = 3'h1 == total_offset_28[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1652 = 3'h2 == total_offset_28[2:0] ? args_2 : _GEN_1651; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1653 = 3'h3 == total_offset_28[2:0] ? args_3 : _GEN_1652; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1654 = 3'h4 == total_offset_28[2:0] ? args_4 : _GEN_1653; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1655 = 3'h5 == total_offset_28[2:0] ? args_5 : _GEN_1654; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1656 = 3'h6 == total_offset_28[2:0] ? args_6 : _GEN_1655; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_3_4 = 8'h4 < _GEN_3382 ? _GEN_1656 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_29 = _GEN_3383 + 8'h5; // @[executor.scala 163:56]
  wire [7:0] _GEN_1659 = 3'h1 == total_offset_29[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1660 = 3'h2 == total_offset_29[2:0] ? args_2 : _GEN_1659; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1661 = 3'h3 == total_offset_29[2:0] ? args_3 : _GEN_1660; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1662 = 3'h4 == total_offset_29[2:0] ? args_4 : _GEN_1661; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1663 = 3'h5 == total_offset_29[2:0] ? args_5 : _GEN_1662; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1664 = 3'h6 == total_offset_29[2:0] ? args_6 : _GEN_1663; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_3_5 = 8'h5 < _GEN_3382 ? _GEN_1664 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_30 = _GEN_3383 + 8'h6; // @[executor.scala 163:56]
  wire [7:0] _GEN_1667 = 3'h1 == total_offset_30[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1668 = 3'h2 == total_offset_30[2:0] ? args_2 : _GEN_1667; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1669 = 3'h3 == total_offset_30[2:0] ? args_3 : _GEN_1668; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1670 = 3'h4 == total_offset_30[2:0] ? args_4 : _GEN_1669; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1671 = 3'h5 == total_offset_30[2:0] ? args_5 : _GEN_1670; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_1672 = 3'h6 == total_offset_30[2:0] ? args_6 : _GEN_1671; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_3_6 = 8'h6 < _GEN_3382 ? _GEN_1672 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [63:0] _io_field_out_1_T_1 = {bytes_3_0,bytes_3_1,bytes_3_2,bytes_3_3,bytes_3_4,bytes_3_5,bytes_3_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_1_hi_12 = io_field_out_1_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_1_T_4 = {io_field_out_1_hi_12,io_field_out_1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_1682 = 4'ha == opcode_1 ? _io_field_out_1_T_1 : _io_field_out_1_T_4; // @[executor.scala 157:51 executor.scala 170:37 executor.scala 173:37]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_2_lo = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire  from_header_2 = length_2 != 8'h0; // @[executor.scala 141:41]
  wire [8:0] _total_offset_T_32 = {{1'd0}, offset_2}; // @[executor.scala 148:53]
  wire [7:0] total_offset_32 = _total_offset_T_32[7:0]; // @[executor.scala 148:53]
  wire [7:0] _GEN_1685 = 7'h1 == total_offset_32[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1686 = 7'h2 == total_offset_32[6:0] ? phv_data_2 : _GEN_1685; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1687 = 7'h3 == total_offset_32[6:0] ? phv_data_3 : _GEN_1686; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1688 = 7'h4 == total_offset_32[6:0] ? phv_data_4 : _GEN_1687; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1689 = 7'h5 == total_offset_32[6:0] ? phv_data_5 : _GEN_1688; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1690 = 7'h6 == total_offset_32[6:0] ? phv_data_6 : _GEN_1689; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1691 = 7'h7 == total_offset_32[6:0] ? phv_data_7 : _GEN_1690; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1692 = 7'h8 == total_offset_32[6:0] ? phv_data_8 : _GEN_1691; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1693 = 7'h9 == total_offset_32[6:0] ? phv_data_9 : _GEN_1692; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1694 = 7'ha == total_offset_32[6:0] ? phv_data_10 : _GEN_1693; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1695 = 7'hb == total_offset_32[6:0] ? phv_data_11 : _GEN_1694; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1696 = 7'hc == total_offset_32[6:0] ? phv_data_12 : _GEN_1695; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1697 = 7'hd == total_offset_32[6:0] ? phv_data_13 : _GEN_1696; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1698 = 7'he == total_offset_32[6:0] ? phv_data_14 : _GEN_1697; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1699 = 7'hf == total_offset_32[6:0] ? phv_data_15 : _GEN_1698; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1700 = 7'h10 == total_offset_32[6:0] ? phv_data_16 : _GEN_1699; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1701 = 7'h11 == total_offset_32[6:0] ? phv_data_17 : _GEN_1700; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1702 = 7'h12 == total_offset_32[6:0] ? phv_data_18 : _GEN_1701; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1703 = 7'h13 == total_offset_32[6:0] ? phv_data_19 : _GEN_1702; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1704 = 7'h14 == total_offset_32[6:0] ? phv_data_20 : _GEN_1703; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1705 = 7'h15 == total_offset_32[6:0] ? phv_data_21 : _GEN_1704; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1706 = 7'h16 == total_offset_32[6:0] ? phv_data_22 : _GEN_1705; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1707 = 7'h17 == total_offset_32[6:0] ? phv_data_23 : _GEN_1706; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1708 = 7'h18 == total_offset_32[6:0] ? phv_data_24 : _GEN_1707; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1709 = 7'h19 == total_offset_32[6:0] ? phv_data_25 : _GEN_1708; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1710 = 7'h1a == total_offset_32[6:0] ? phv_data_26 : _GEN_1709; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1711 = 7'h1b == total_offset_32[6:0] ? phv_data_27 : _GEN_1710; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1712 = 7'h1c == total_offset_32[6:0] ? phv_data_28 : _GEN_1711; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1713 = 7'h1d == total_offset_32[6:0] ? phv_data_29 : _GEN_1712; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1714 = 7'h1e == total_offset_32[6:0] ? phv_data_30 : _GEN_1713; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1715 = 7'h1f == total_offset_32[6:0] ? phv_data_31 : _GEN_1714; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1716 = 7'h20 == total_offset_32[6:0] ? phv_data_32 : _GEN_1715; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1717 = 7'h21 == total_offset_32[6:0] ? phv_data_33 : _GEN_1716; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1718 = 7'h22 == total_offset_32[6:0] ? phv_data_34 : _GEN_1717; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1719 = 7'h23 == total_offset_32[6:0] ? phv_data_35 : _GEN_1718; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1720 = 7'h24 == total_offset_32[6:0] ? phv_data_36 : _GEN_1719; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1721 = 7'h25 == total_offset_32[6:0] ? phv_data_37 : _GEN_1720; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1722 = 7'h26 == total_offset_32[6:0] ? phv_data_38 : _GEN_1721; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1723 = 7'h27 == total_offset_32[6:0] ? phv_data_39 : _GEN_1722; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1724 = 7'h28 == total_offset_32[6:0] ? phv_data_40 : _GEN_1723; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1725 = 7'h29 == total_offset_32[6:0] ? phv_data_41 : _GEN_1724; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1726 = 7'h2a == total_offset_32[6:0] ? phv_data_42 : _GEN_1725; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1727 = 7'h2b == total_offset_32[6:0] ? phv_data_43 : _GEN_1726; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1728 = 7'h2c == total_offset_32[6:0] ? phv_data_44 : _GEN_1727; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1729 = 7'h2d == total_offset_32[6:0] ? phv_data_45 : _GEN_1728; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1730 = 7'h2e == total_offset_32[6:0] ? phv_data_46 : _GEN_1729; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1731 = 7'h2f == total_offset_32[6:0] ? phv_data_47 : _GEN_1730; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1732 = 7'h30 == total_offset_32[6:0] ? phv_data_48 : _GEN_1731; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1733 = 7'h31 == total_offset_32[6:0] ? phv_data_49 : _GEN_1732; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1734 = 7'h32 == total_offset_32[6:0] ? phv_data_50 : _GEN_1733; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1735 = 7'h33 == total_offset_32[6:0] ? phv_data_51 : _GEN_1734; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1736 = 7'h34 == total_offset_32[6:0] ? phv_data_52 : _GEN_1735; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1737 = 7'h35 == total_offset_32[6:0] ? phv_data_53 : _GEN_1736; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1738 = 7'h36 == total_offset_32[6:0] ? phv_data_54 : _GEN_1737; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1739 = 7'h37 == total_offset_32[6:0] ? phv_data_55 : _GEN_1738; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1740 = 7'h38 == total_offset_32[6:0] ? phv_data_56 : _GEN_1739; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1741 = 7'h39 == total_offset_32[6:0] ? phv_data_57 : _GEN_1740; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1742 = 7'h3a == total_offset_32[6:0] ? phv_data_58 : _GEN_1741; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1743 = 7'h3b == total_offset_32[6:0] ? phv_data_59 : _GEN_1742; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1744 = 7'h3c == total_offset_32[6:0] ? phv_data_60 : _GEN_1743; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1745 = 7'h3d == total_offset_32[6:0] ? phv_data_61 : _GEN_1744; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1746 = 7'h3e == total_offset_32[6:0] ? phv_data_62 : _GEN_1745; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1747 = 7'h3f == total_offset_32[6:0] ? phv_data_63 : _GEN_1746; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1748 = 7'h40 == total_offset_32[6:0] ? phv_data_64 : _GEN_1747; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1749 = 7'h41 == total_offset_32[6:0] ? phv_data_65 : _GEN_1748; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1750 = 7'h42 == total_offset_32[6:0] ? phv_data_66 : _GEN_1749; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1751 = 7'h43 == total_offset_32[6:0] ? phv_data_67 : _GEN_1750; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1752 = 7'h44 == total_offset_32[6:0] ? phv_data_68 : _GEN_1751; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1753 = 7'h45 == total_offset_32[6:0] ? phv_data_69 : _GEN_1752; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1754 = 7'h46 == total_offset_32[6:0] ? phv_data_70 : _GEN_1753; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1755 = 7'h47 == total_offset_32[6:0] ? phv_data_71 : _GEN_1754; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1756 = 7'h48 == total_offset_32[6:0] ? phv_data_72 : _GEN_1755; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1757 = 7'h49 == total_offset_32[6:0] ? phv_data_73 : _GEN_1756; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1758 = 7'h4a == total_offset_32[6:0] ? phv_data_74 : _GEN_1757; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1759 = 7'h4b == total_offset_32[6:0] ? phv_data_75 : _GEN_1758; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1760 = 7'h4c == total_offset_32[6:0] ? phv_data_76 : _GEN_1759; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1761 = 7'h4d == total_offset_32[6:0] ? phv_data_77 : _GEN_1760; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1762 = 7'h4e == total_offset_32[6:0] ? phv_data_78 : _GEN_1761; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1763 = 7'h4f == total_offset_32[6:0] ? phv_data_79 : _GEN_1762; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1764 = 7'h50 == total_offset_32[6:0] ? phv_data_80 : _GEN_1763; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1765 = 7'h51 == total_offset_32[6:0] ? phv_data_81 : _GEN_1764; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1766 = 7'h52 == total_offset_32[6:0] ? phv_data_82 : _GEN_1765; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1767 = 7'h53 == total_offset_32[6:0] ? phv_data_83 : _GEN_1766; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1768 = 7'h54 == total_offset_32[6:0] ? phv_data_84 : _GEN_1767; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1769 = 7'h55 == total_offset_32[6:0] ? phv_data_85 : _GEN_1768; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1770 = 7'h56 == total_offset_32[6:0] ? phv_data_86 : _GEN_1769; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1771 = 7'h57 == total_offset_32[6:0] ? phv_data_87 : _GEN_1770; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1772 = 7'h58 == total_offset_32[6:0] ? phv_data_88 : _GEN_1771; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1773 = 7'h59 == total_offset_32[6:0] ? phv_data_89 : _GEN_1772; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1774 = 7'h5a == total_offset_32[6:0] ? phv_data_90 : _GEN_1773; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1775 = 7'h5b == total_offset_32[6:0] ? phv_data_91 : _GEN_1774; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1776 = 7'h5c == total_offset_32[6:0] ? phv_data_92 : _GEN_1775; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1777 = 7'h5d == total_offset_32[6:0] ? phv_data_93 : _GEN_1776; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1778 = 7'h5e == total_offset_32[6:0] ? phv_data_94 : _GEN_1777; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1779 = 7'h5f == total_offset_32[6:0] ? phv_data_95 : _GEN_1778; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_0 = 8'h0 < length_2 ? _GEN_1779 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_33 = offset_2 + 8'h1; // @[executor.scala 148:53]
  wire [7:0] _GEN_1782 = 7'h1 == total_offset_33[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1783 = 7'h2 == total_offset_33[6:0] ? phv_data_2 : _GEN_1782; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1784 = 7'h3 == total_offset_33[6:0] ? phv_data_3 : _GEN_1783; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1785 = 7'h4 == total_offset_33[6:0] ? phv_data_4 : _GEN_1784; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1786 = 7'h5 == total_offset_33[6:0] ? phv_data_5 : _GEN_1785; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1787 = 7'h6 == total_offset_33[6:0] ? phv_data_6 : _GEN_1786; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1788 = 7'h7 == total_offset_33[6:0] ? phv_data_7 : _GEN_1787; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1789 = 7'h8 == total_offset_33[6:0] ? phv_data_8 : _GEN_1788; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1790 = 7'h9 == total_offset_33[6:0] ? phv_data_9 : _GEN_1789; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1791 = 7'ha == total_offset_33[6:0] ? phv_data_10 : _GEN_1790; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1792 = 7'hb == total_offset_33[6:0] ? phv_data_11 : _GEN_1791; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1793 = 7'hc == total_offset_33[6:0] ? phv_data_12 : _GEN_1792; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1794 = 7'hd == total_offset_33[6:0] ? phv_data_13 : _GEN_1793; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1795 = 7'he == total_offset_33[6:0] ? phv_data_14 : _GEN_1794; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1796 = 7'hf == total_offset_33[6:0] ? phv_data_15 : _GEN_1795; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1797 = 7'h10 == total_offset_33[6:0] ? phv_data_16 : _GEN_1796; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1798 = 7'h11 == total_offset_33[6:0] ? phv_data_17 : _GEN_1797; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1799 = 7'h12 == total_offset_33[6:0] ? phv_data_18 : _GEN_1798; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1800 = 7'h13 == total_offset_33[6:0] ? phv_data_19 : _GEN_1799; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1801 = 7'h14 == total_offset_33[6:0] ? phv_data_20 : _GEN_1800; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1802 = 7'h15 == total_offset_33[6:0] ? phv_data_21 : _GEN_1801; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1803 = 7'h16 == total_offset_33[6:0] ? phv_data_22 : _GEN_1802; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1804 = 7'h17 == total_offset_33[6:0] ? phv_data_23 : _GEN_1803; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1805 = 7'h18 == total_offset_33[6:0] ? phv_data_24 : _GEN_1804; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1806 = 7'h19 == total_offset_33[6:0] ? phv_data_25 : _GEN_1805; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1807 = 7'h1a == total_offset_33[6:0] ? phv_data_26 : _GEN_1806; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1808 = 7'h1b == total_offset_33[6:0] ? phv_data_27 : _GEN_1807; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1809 = 7'h1c == total_offset_33[6:0] ? phv_data_28 : _GEN_1808; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1810 = 7'h1d == total_offset_33[6:0] ? phv_data_29 : _GEN_1809; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1811 = 7'h1e == total_offset_33[6:0] ? phv_data_30 : _GEN_1810; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1812 = 7'h1f == total_offset_33[6:0] ? phv_data_31 : _GEN_1811; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1813 = 7'h20 == total_offset_33[6:0] ? phv_data_32 : _GEN_1812; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1814 = 7'h21 == total_offset_33[6:0] ? phv_data_33 : _GEN_1813; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1815 = 7'h22 == total_offset_33[6:0] ? phv_data_34 : _GEN_1814; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1816 = 7'h23 == total_offset_33[6:0] ? phv_data_35 : _GEN_1815; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1817 = 7'h24 == total_offset_33[6:0] ? phv_data_36 : _GEN_1816; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1818 = 7'h25 == total_offset_33[6:0] ? phv_data_37 : _GEN_1817; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1819 = 7'h26 == total_offset_33[6:0] ? phv_data_38 : _GEN_1818; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1820 = 7'h27 == total_offset_33[6:0] ? phv_data_39 : _GEN_1819; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1821 = 7'h28 == total_offset_33[6:0] ? phv_data_40 : _GEN_1820; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1822 = 7'h29 == total_offset_33[6:0] ? phv_data_41 : _GEN_1821; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1823 = 7'h2a == total_offset_33[6:0] ? phv_data_42 : _GEN_1822; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1824 = 7'h2b == total_offset_33[6:0] ? phv_data_43 : _GEN_1823; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1825 = 7'h2c == total_offset_33[6:0] ? phv_data_44 : _GEN_1824; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1826 = 7'h2d == total_offset_33[6:0] ? phv_data_45 : _GEN_1825; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1827 = 7'h2e == total_offset_33[6:0] ? phv_data_46 : _GEN_1826; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1828 = 7'h2f == total_offset_33[6:0] ? phv_data_47 : _GEN_1827; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1829 = 7'h30 == total_offset_33[6:0] ? phv_data_48 : _GEN_1828; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1830 = 7'h31 == total_offset_33[6:0] ? phv_data_49 : _GEN_1829; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1831 = 7'h32 == total_offset_33[6:0] ? phv_data_50 : _GEN_1830; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1832 = 7'h33 == total_offset_33[6:0] ? phv_data_51 : _GEN_1831; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1833 = 7'h34 == total_offset_33[6:0] ? phv_data_52 : _GEN_1832; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1834 = 7'h35 == total_offset_33[6:0] ? phv_data_53 : _GEN_1833; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1835 = 7'h36 == total_offset_33[6:0] ? phv_data_54 : _GEN_1834; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1836 = 7'h37 == total_offset_33[6:0] ? phv_data_55 : _GEN_1835; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1837 = 7'h38 == total_offset_33[6:0] ? phv_data_56 : _GEN_1836; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1838 = 7'h39 == total_offset_33[6:0] ? phv_data_57 : _GEN_1837; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1839 = 7'h3a == total_offset_33[6:0] ? phv_data_58 : _GEN_1838; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1840 = 7'h3b == total_offset_33[6:0] ? phv_data_59 : _GEN_1839; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1841 = 7'h3c == total_offset_33[6:0] ? phv_data_60 : _GEN_1840; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1842 = 7'h3d == total_offset_33[6:0] ? phv_data_61 : _GEN_1841; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1843 = 7'h3e == total_offset_33[6:0] ? phv_data_62 : _GEN_1842; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1844 = 7'h3f == total_offset_33[6:0] ? phv_data_63 : _GEN_1843; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1845 = 7'h40 == total_offset_33[6:0] ? phv_data_64 : _GEN_1844; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1846 = 7'h41 == total_offset_33[6:0] ? phv_data_65 : _GEN_1845; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1847 = 7'h42 == total_offset_33[6:0] ? phv_data_66 : _GEN_1846; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1848 = 7'h43 == total_offset_33[6:0] ? phv_data_67 : _GEN_1847; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1849 = 7'h44 == total_offset_33[6:0] ? phv_data_68 : _GEN_1848; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1850 = 7'h45 == total_offset_33[6:0] ? phv_data_69 : _GEN_1849; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1851 = 7'h46 == total_offset_33[6:0] ? phv_data_70 : _GEN_1850; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1852 = 7'h47 == total_offset_33[6:0] ? phv_data_71 : _GEN_1851; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1853 = 7'h48 == total_offset_33[6:0] ? phv_data_72 : _GEN_1852; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1854 = 7'h49 == total_offset_33[6:0] ? phv_data_73 : _GEN_1853; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1855 = 7'h4a == total_offset_33[6:0] ? phv_data_74 : _GEN_1854; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1856 = 7'h4b == total_offset_33[6:0] ? phv_data_75 : _GEN_1855; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1857 = 7'h4c == total_offset_33[6:0] ? phv_data_76 : _GEN_1856; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1858 = 7'h4d == total_offset_33[6:0] ? phv_data_77 : _GEN_1857; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1859 = 7'h4e == total_offset_33[6:0] ? phv_data_78 : _GEN_1858; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1860 = 7'h4f == total_offset_33[6:0] ? phv_data_79 : _GEN_1859; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1861 = 7'h50 == total_offset_33[6:0] ? phv_data_80 : _GEN_1860; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1862 = 7'h51 == total_offset_33[6:0] ? phv_data_81 : _GEN_1861; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1863 = 7'h52 == total_offset_33[6:0] ? phv_data_82 : _GEN_1862; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1864 = 7'h53 == total_offset_33[6:0] ? phv_data_83 : _GEN_1863; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1865 = 7'h54 == total_offset_33[6:0] ? phv_data_84 : _GEN_1864; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1866 = 7'h55 == total_offset_33[6:0] ? phv_data_85 : _GEN_1865; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1867 = 7'h56 == total_offset_33[6:0] ? phv_data_86 : _GEN_1866; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1868 = 7'h57 == total_offset_33[6:0] ? phv_data_87 : _GEN_1867; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1869 = 7'h58 == total_offset_33[6:0] ? phv_data_88 : _GEN_1868; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1870 = 7'h59 == total_offset_33[6:0] ? phv_data_89 : _GEN_1869; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1871 = 7'h5a == total_offset_33[6:0] ? phv_data_90 : _GEN_1870; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1872 = 7'h5b == total_offset_33[6:0] ? phv_data_91 : _GEN_1871; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1873 = 7'h5c == total_offset_33[6:0] ? phv_data_92 : _GEN_1872; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1874 = 7'h5d == total_offset_33[6:0] ? phv_data_93 : _GEN_1873; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1875 = 7'h5e == total_offset_33[6:0] ? phv_data_94 : _GEN_1874; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1876 = 7'h5f == total_offset_33[6:0] ? phv_data_95 : _GEN_1875; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_1 = 8'h1 < length_2 ? _GEN_1876 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_34 = offset_2 + 8'h2; // @[executor.scala 148:53]
  wire [7:0] _GEN_1879 = 7'h1 == total_offset_34[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1880 = 7'h2 == total_offset_34[6:0] ? phv_data_2 : _GEN_1879; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1881 = 7'h3 == total_offset_34[6:0] ? phv_data_3 : _GEN_1880; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1882 = 7'h4 == total_offset_34[6:0] ? phv_data_4 : _GEN_1881; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1883 = 7'h5 == total_offset_34[6:0] ? phv_data_5 : _GEN_1882; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1884 = 7'h6 == total_offset_34[6:0] ? phv_data_6 : _GEN_1883; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1885 = 7'h7 == total_offset_34[6:0] ? phv_data_7 : _GEN_1884; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1886 = 7'h8 == total_offset_34[6:0] ? phv_data_8 : _GEN_1885; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1887 = 7'h9 == total_offset_34[6:0] ? phv_data_9 : _GEN_1886; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1888 = 7'ha == total_offset_34[6:0] ? phv_data_10 : _GEN_1887; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1889 = 7'hb == total_offset_34[6:0] ? phv_data_11 : _GEN_1888; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1890 = 7'hc == total_offset_34[6:0] ? phv_data_12 : _GEN_1889; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1891 = 7'hd == total_offset_34[6:0] ? phv_data_13 : _GEN_1890; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1892 = 7'he == total_offset_34[6:0] ? phv_data_14 : _GEN_1891; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1893 = 7'hf == total_offset_34[6:0] ? phv_data_15 : _GEN_1892; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1894 = 7'h10 == total_offset_34[6:0] ? phv_data_16 : _GEN_1893; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1895 = 7'h11 == total_offset_34[6:0] ? phv_data_17 : _GEN_1894; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1896 = 7'h12 == total_offset_34[6:0] ? phv_data_18 : _GEN_1895; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1897 = 7'h13 == total_offset_34[6:0] ? phv_data_19 : _GEN_1896; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1898 = 7'h14 == total_offset_34[6:0] ? phv_data_20 : _GEN_1897; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1899 = 7'h15 == total_offset_34[6:0] ? phv_data_21 : _GEN_1898; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1900 = 7'h16 == total_offset_34[6:0] ? phv_data_22 : _GEN_1899; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1901 = 7'h17 == total_offset_34[6:0] ? phv_data_23 : _GEN_1900; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1902 = 7'h18 == total_offset_34[6:0] ? phv_data_24 : _GEN_1901; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1903 = 7'h19 == total_offset_34[6:0] ? phv_data_25 : _GEN_1902; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1904 = 7'h1a == total_offset_34[6:0] ? phv_data_26 : _GEN_1903; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1905 = 7'h1b == total_offset_34[6:0] ? phv_data_27 : _GEN_1904; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1906 = 7'h1c == total_offset_34[6:0] ? phv_data_28 : _GEN_1905; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1907 = 7'h1d == total_offset_34[6:0] ? phv_data_29 : _GEN_1906; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1908 = 7'h1e == total_offset_34[6:0] ? phv_data_30 : _GEN_1907; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1909 = 7'h1f == total_offset_34[6:0] ? phv_data_31 : _GEN_1908; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1910 = 7'h20 == total_offset_34[6:0] ? phv_data_32 : _GEN_1909; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1911 = 7'h21 == total_offset_34[6:0] ? phv_data_33 : _GEN_1910; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1912 = 7'h22 == total_offset_34[6:0] ? phv_data_34 : _GEN_1911; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1913 = 7'h23 == total_offset_34[6:0] ? phv_data_35 : _GEN_1912; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1914 = 7'h24 == total_offset_34[6:0] ? phv_data_36 : _GEN_1913; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1915 = 7'h25 == total_offset_34[6:0] ? phv_data_37 : _GEN_1914; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1916 = 7'h26 == total_offset_34[6:0] ? phv_data_38 : _GEN_1915; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1917 = 7'h27 == total_offset_34[6:0] ? phv_data_39 : _GEN_1916; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1918 = 7'h28 == total_offset_34[6:0] ? phv_data_40 : _GEN_1917; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1919 = 7'h29 == total_offset_34[6:0] ? phv_data_41 : _GEN_1918; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1920 = 7'h2a == total_offset_34[6:0] ? phv_data_42 : _GEN_1919; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1921 = 7'h2b == total_offset_34[6:0] ? phv_data_43 : _GEN_1920; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1922 = 7'h2c == total_offset_34[6:0] ? phv_data_44 : _GEN_1921; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1923 = 7'h2d == total_offset_34[6:0] ? phv_data_45 : _GEN_1922; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1924 = 7'h2e == total_offset_34[6:0] ? phv_data_46 : _GEN_1923; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1925 = 7'h2f == total_offset_34[6:0] ? phv_data_47 : _GEN_1924; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1926 = 7'h30 == total_offset_34[6:0] ? phv_data_48 : _GEN_1925; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1927 = 7'h31 == total_offset_34[6:0] ? phv_data_49 : _GEN_1926; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1928 = 7'h32 == total_offset_34[6:0] ? phv_data_50 : _GEN_1927; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1929 = 7'h33 == total_offset_34[6:0] ? phv_data_51 : _GEN_1928; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1930 = 7'h34 == total_offset_34[6:0] ? phv_data_52 : _GEN_1929; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1931 = 7'h35 == total_offset_34[6:0] ? phv_data_53 : _GEN_1930; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1932 = 7'h36 == total_offset_34[6:0] ? phv_data_54 : _GEN_1931; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1933 = 7'h37 == total_offset_34[6:0] ? phv_data_55 : _GEN_1932; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1934 = 7'h38 == total_offset_34[6:0] ? phv_data_56 : _GEN_1933; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1935 = 7'h39 == total_offset_34[6:0] ? phv_data_57 : _GEN_1934; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1936 = 7'h3a == total_offset_34[6:0] ? phv_data_58 : _GEN_1935; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1937 = 7'h3b == total_offset_34[6:0] ? phv_data_59 : _GEN_1936; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1938 = 7'h3c == total_offset_34[6:0] ? phv_data_60 : _GEN_1937; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1939 = 7'h3d == total_offset_34[6:0] ? phv_data_61 : _GEN_1938; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1940 = 7'h3e == total_offset_34[6:0] ? phv_data_62 : _GEN_1939; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1941 = 7'h3f == total_offset_34[6:0] ? phv_data_63 : _GEN_1940; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1942 = 7'h40 == total_offset_34[6:0] ? phv_data_64 : _GEN_1941; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1943 = 7'h41 == total_offset_34[6:0] ? phv_data_65 : _GEN_1942; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1944 = 7'h42 == total_offset_34[6:0] ? phv_data_66 : _GEN_1943; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1945 = 7'h43 == total_offset_34[6:0] ? phv_data_67 : _GEN_1944; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1946 = 7'h44 == total_offset_34[6:0] ? phv_data_68 : _GEN_1945; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1947 = 7'h45 == total_offset_34[6:0] ? phv_data_69 : _GEN_1946; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1948 = 7'h46 == total_offset_34[6:0] ? phv_data_70 : _GEN_1947; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1949 = 7'h47 == total_offset_34[6:0] ? phv_data_71 : _GEN_1948; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1950 = 7'h48 == total_offset_34[6:0] ? phv_data_72 : _GEN_1949; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1951 = 7'h49 == total_offset_34[6:0] ? phv_data_73 : _GEN_1950; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1952 = 7'h4a == total_offset_34[6:0] ? phv_data_74 : _GEN_1951; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1953 = 7'h4b == total_offset_34[6:0] ? phv_data_75 : _GEN_1952; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1954 = 7'h4c == total_offset_34[6:0] ? phv_data_76 : _GEN_1953; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1955 = 7'h4d == total_offset_34[6:0] ? phv_data_77 : _GEN_1954; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1956 = 7'h4e == total_offset_34[6:0] ? phv_data_78 : _GEN_1955; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1957 = 7'h4f == total_offset_34[6:0] ? phv_data_79 : _GEN_1956; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1958 = 7'h50 == total_offset_34[6:0] ? phv_data_80 : _GEN_1957; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1959 = 7'h51 == total_offset_34[6:0] ? phv_data_81 : _GEN_1958; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1960 = 7'h52 == total_offset_34[6:0] ? phv_data_82 : _GEN_1959; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1961 = 7'h53 == total_offset_34[6:0] ? phv_data_83 : _GEN_1960; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1962 = 7'h54 == total_offset_34[6:0] ? phv_data_84 : _GEN_1961; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1963 = 7'h55 == total_offset_34[6:0] ? phv_data_85 : _GEN_1962; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1964 = 7'h56 == total_offset_34[6:0] ? phv_data_86 : _GEN_1963; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1965 = 7'h57 == total_offset_34[6:0] ? phv_data_87 : _GEN_1964; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1966 = 7'h58 == total_offset_34[6:0] ? phv_data_88 : _GEN_1965; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1967 = 7'h59 == total_offset_34[6:0] ? phv_data_89 : _GEN_1966; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1968 = 7'h5a == total_offset_34[6:0] ? phv_data_90 : _GEN_1967; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1969 = 7'h5b == total_offset_34[6:0] ? phv_data_91 : _GEN_1968; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1970 = 7'h5c == total_offset_34[6:0] ? phv_data_92 : _GEN_1969; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1971 = 7'h5d == total_offset_34[6:0] ? phv_data_93 : _GEN_1970; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1972 = 7'h5e == total_offset_34[6:0] ? phv_data_94 : _GEN_1971; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1973 = 7'h5f == total_offset_34[6:0] ? phv_data_95 : _GEN_1972; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_2 = 8'h2 < length_2 ? _GEN_1973 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_35 = offset_2 + 8'h3; // @[executor.scala 148:53]
  wire [7:0] _GEN_1976 = 7'h1 == total_offset_35[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1977 = 7'h2 == total_offset_35[6:0] ? phv_data_2 : _GEN_1976; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1978 = 7'h3 == total_offset_35[6:0] ? phv_data_3 : _GEN_1977; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1979 = 7'h4 == total_offset_35[6:0] ? phv_data_4 : _GEN_1978; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1980 = 7'h5 == total_offset_35[6:0] ? phv_data_5 : _GEN_1979; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1981 = 7'h6 == total_offset_35[6:0] ? phv_data_6 : _GEN_1980; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1982 = 7'h7 == total_offset_35[6:0] ? phv_data_7 : _GEN_1981; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1983 = 7'h8 == total_offset_35[6:0] ? phv_data_8 : _GEN_1982; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1984 = 7'h9 == total_offset_35[6:0] ? phv_data_9 : _GEN_1983; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1985 = 7'ha == total_offset_35[6:0] ? phv_data_10 : _GEN_1984; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1986 = 7'hb == total_offset_35[6:0] ? phv_data_11 : _GEN_1985; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1987 = 7'hc == total_offset_35[6:0] ? phv_data_12 : _GEN_1986; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1988 = 7'hd == total_offset_35[6:0] ? phv_data_13 : _GEN_1987; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1989 = 7'he == total_offset_35[6:0] ? phv_data_14 : _GEN_1988; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1990 = 7'hf == total_offset_35[6:0] ? phv_data_15 : _GEN_1989; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1991 = 7'h10 == total_offset_35[6:0] ? phv_data_16 : _GEN_1990; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1992 = 7'h11 == total_offset_35[6:0] ? phv_data_17 : _GEN_1991; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1993 = 7'h12 == total_offset_35[6:0] ? phv_data_18 : _GEN_1992; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1994 = 7'h13 == total_offset_35[6:0] ? phv_data_19 : _GEN_1993; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1995 = 7'h14 == total_offset_35[6:0] ? phv_data_20 : _GEN_1994; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1996 = 7'h15 == total_offset_35[6:0] ? phv_data_21 : _GEN_1995; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1997 = 7'h16 == total_offset_35[6:0] ? phv_data_22 : _GEN_1996; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1998 = 7'h17 == total_offset_35[6:0] ? phv_data_23 : _GEN_1997; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_1999 = 7'h18 == total_offset_35[6:0] ? phv_data_24 : _GEN_1998; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2000 = 7'h19 == total_offset_35[6:0] ? phv_data_25 : _GEN_1999; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2001 = 7'h1a == total_offset_35[6:0] ? phv_data_26 : _GEN_2000; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2002 = 7'h1b == total_offset_35[6:0] ? phv_data_27 : _GEN_2001; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2003 = 7'h1c == total_offset_35[6:0] ? phv_data_28 : _GEN_2002; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2004 = 7'h1d == total_offset_35[6:0] ? phv_data_29 : _GEN_2003; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2005 = 7'h1e == total_offset_35[6:0] ? phv_data_30 : _GEN_2004; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2006 = 7'h1f == total_offset_35[6:0] ? phv_data_31 : _GEN_2005; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2007 = 7'h20 == total_offset_35[6:0] ? phv_data_32 : _GEN_2006; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2008 = 7'h21 == total_offset_35[6:0] ? phv_data_33 : _GEN_2007; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2009 = 7'h22 == total_offset_35[6:0] ? phv_data_34 : _GEN_2008; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2010 = 7'h23 == total_offset_35[6:0] ? phv_data_35 : _GEN_2009; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2011 = 7'h24 == total_offset_35[6:0] ? phv_data_36 : _GEN_2010; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2012 = 7'h25 == total_offset_35[6:0] ? phv_data_37 : _GEN_2011; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2013 = 7'h26 == total_offset_35[6:0] ? phv_data_38 : _GEN_2012; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2014 = 7'h27 == total_offset_35[6:0] ? phv_data_39 : _GEN_2013; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2015 = 7'h28 == total_offset_35[6:0] ? phv_data_40 : _GEN_2014; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2016 = 7'h29 == total_offset_35[6:0] ? phv_data_41 : _GEN_2015; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2017 = 7'h2a == total_offset_35[6:0] ? phv_data_42 : _GEN_2016; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2018 = 7'h2b == total_offset_35[6:0] ? phv_data_43 : _GEN_2017; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2019 = 7'h2c == total_offset_35[6:0] ? phv_data_44 : _GEN_2018; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2020 = 7'h2d == total_offset_35[6:0] ? phv_data_45 : _GEN_2019; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2021 = 7'h2e == total_offset_35[6:0] ? phv_data_46 : _GEN_2020; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2022 = 7'h2f == total_offset_35[6:0] ? phv_data_47 : _GEN_2021; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2023 = 7'h30 == total_offset_35[6:0] ? phv_data_48 : _GEN_2022; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2024 = 7'h31 == total_offset_35[6:0] ? phv_data_49 : _GEN_2023; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2025 = 7'h32 == total_offset_35[6:0] ? phv_data_50 : _GEN_2024; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2026 = 7'h33 == total_offset_35[6:0] ? phv_data_51 : _GEN_2025; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2027 = 7'h34 == total_offset_35[6:0] ? phv_data_52 : _GEN_2026; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2028 = 7'h35 == total_offset_35[6:0] ? phv_data_53 : _GEN_2027; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2029 = 7'h36 == total_offset_35[6:0] ? phv_data_54 : _GEN_2028; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2030 = 7'h37 == total_offset_35[6:0] ? phv_data_55 : _GEN_2029; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2031 = 7'h38 == total_offset_35[6:0] ? phv_data_56 : _GEN_2030; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2032 = 7'h39 == total_offset_35[6:0] ? phv_data_57 : _GEN_2031; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2033 = 7'h3a == total_offset_35[6:0] ? phv_data_58 : _GEN_2032; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2034 = 7'h3b == total_offset_35[6:0] ? phv_data_59 : _GEN_2033; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2035 = 7'h3c == total_offset_35[6:0] ? phv_data_60 : _GEN_2034; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2036 = 7'h3d == total_offset_35[6:0] ? phv_data_61 : _GEN_2035; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2037 = 7'h3e == total_offset_35[6:0] ? phv_data_62 : _GEN_2036; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2038 = 7'h3f == total_offset_35[6:0] ? phv_data_63 : _GEN_2037; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2039 = 7'h40 == total_offset_35[6:0] ? phv_data_64 : _GEN_2038; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2040 = 7'h41 == total_offset_35[6:0] ? phv_data_65 : _GEN_2039; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2041 = 7'h42 == total_offset_35[6:0] ? phv_data_66 : _GEN_2040; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2042 = 7'h43 == total_offset_35[6:0] ? phv_data_67 : _GEN_2041; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2043 = 7'h44 == total_offset_35[6:0] ? phv_data_68 : _GEN_2042; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2044 = 7'h45 == total_offset_35[6:0] ? phv_data_69 : _GEN_2043; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2045 = 7'h46 == total_offset_35[6:0] ? phv_data_70 : _GEN_2044; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2046 = 7'h47 == total_offset_35[6:0] ? phv_data_71 : _GEN_2045; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2047 = 7'h48 == total_offset_35[6:0] ? phv_data_72 : _GEN_2046; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2048 = 7'h49 == total_offset_35[6:0] ? phv_data_73 : _GEN_2047; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2049 = 7'h4a == total_offset_35[6:0] ? phv_data_74 : _GEN_2048; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2050 = 7'h4b == total_offset_35[6:0] ? phv_data_75 : _GEN_2049; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2051 = 7'h4c == total_offset_35[6:0] ? phv_data_76 : _GEN_2050; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2052 = 7'h4d == total_offset_35[6:0] ? phv_data_77 : _GEN_2051; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2053 = 7'h4e == total_offset_35[6:0] ? phv_data_78 : _GEN_2052; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2054 = 7'h4f == total_offset_35[6:0] ? phv_data_79 : _GEN_2053; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2055 = 7'h50 == total_offset_35[6:0] ? phv_data_80 : _GEN_2054; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2056 = 7'h51 == total_offset_35[6:0] ? phv_data_81 : _GEN_2055; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2057 = 7'h52 == total_offset_35[6:0] ? phv_data_82 : _GEN_2056; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2058 = 7'h53 == total_offset_35[6:0] ? phv_data_83 : _GEN_2057; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2059 = 7'h54 == total_offset_35[6:0] ? phv_data_84 : _GEN_2058; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2060 = 7'h55 == total_offset_35[6:0] ? phv_data_85 : _GEN_2059; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2061 = 7'h56 == total_offset_35[6:0] ? phv_data_86 : _GEN_2060; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2062 = 7'h57 == total_offset_35[6:0] ? phv_data_87 : _GEN_2061; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2063 = 7'h58 == total_offset_35[6:0] ? phv_data_88 : _GEN_2062; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2064 = 7'h59 == total_offset_35[6:0] ? phv_data_89 : _GEN_2063; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2065 = 7'h5a == total_offset_35[6:0] ? phv_data_90 : _GEN_2064; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2066 = 7'h5b == total_offset_35[6:0] ? phv_data_91 : _GEN_2065; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2067 = 7'h5c == total_offset_35[6:0] ? phv_data_92 : _GEN_2066; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2068 = 7'h5d == total_offset_35[6:0] ? phv_data_93 : _GEN_2067; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2069 = 7'h5e == total_offset_35[6:0] ? phv_data_94 : _GEN_2068; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2070 = 7'h5f == total_offset_35[6:0] ? phv_data_95 : _GEN_2069; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_3 = 8'h3 < length_2 ? _GEN_2070 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_36 = offset_2 + 8'h4; // @[executor.scala 148:53]
  wire [7:0] _GEN_2073 = 7'h1 == total_offset_36[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2074 = 7'h2 == total_offset_36[6:0] ? phv_data_2 : _GEN_2073; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2075 = 7'h3 == total_offset_36[6:0] ? phv_data_3 : _GEN_2074; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2076 = 7'h4 == total_offset_36[6:0] ? phv_data_4 : _GEN_2075; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2077 = 7'h5 == total_offset_36[6:0] ? phv_data_5 : _GEN_2076; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2078 = 7'h6 == total_offset_36[6:0] ? phv_data_6 : _GEN_2077; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2079 = 7'h7 == total_offset_36[6:0] ? phv_data_7 : _GEN_2078; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2080 = 7'h8 == total_offset_36[6:0] ? phv_data_8 : _GEN_2079; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2081 = 7'h9 == total_offset_36[6:0] ? phv_data_9 : _GEN_2080; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2082 = 7'ha == total_offset_36[6:0] ? phv_data_10 : _GEN_2081; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2083 = 7'hb == total_offset_36[6:0] ? phv_data_11 : _GEN_2082; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2084 = 7'hc == total_offset_36[6:0] ? phv_data_12 : _GEN_2083; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2085 = 7'hd == total_offset_36[6:0] ? phv_data_13 : _GEN_2084; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2086 = 7'he == total_offset_36[6:0] ? phv_data_14 : _GEN_2085; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2087 = 7'hf == total_offset_36[6:0] ? phv_data_15 : _GEN_2086; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2088 = 7'h10 == total_offset_36[6:0] ? phv_data_16 : _GEN_2087; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2089 = 7'h11 == total_offset_36[6:0] ? phv_data_17 : _GEN_2088; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2090 = 7'h12 == total_offset_36[6:0] ? phv_data_18 : _GEN_2089; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2091 = 7'h13 == total_offset_36[6:0] ? phv_data_19 : _GEN_2090; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2092 = 7'h14 == total_offset_36[6:0] ? phv_data_20 : _GEN_2091; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2093 = 7'h15 == total_offset_36[6:0] ? phv_data_21 : _GEN_2092; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2094 = 7'h16 == total_offset_36[6:0] ? phv_data_22 : _GEN_2093; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2095 = 7'h17 == total_offset_36[6:0] ? phv_data_23 : _GEN_2094; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2096 = 7'h18 == total_offset_36[6:0] ? phv_data_24 : _GEN_2095; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2097 = 7'h19 == total_offset_36[6:0] ? phv_data_25 : _GEN_2096; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2098 = 7'h1a == total_offset_36[6:0] ? phv_data_26 : _GEN_2097; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2099 = 7'h1b == total_offset_36[6:0] ? phv_data_27 : _GEN_2098; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2100 = 7'h1c == total_offset_36[6:0] ? phv_data_28 : _GEN_2099; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2101 = 7'h1d == total_offset_36[6:0] ? phv_data_29 : _GEN_2100; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2102 = 7'h1e == total_offset_36[6:0] ? phv_data_30 : _GEN_2101; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2103 = 7'h1f == total_offset_36[6:0] ? phv_data_31 : _GEN_2102; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2104 = 7'h20 == total_offset_36[6:0] ? phv_data_32 : _GEN_2103; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2105 = 7'h21 == total_offset_36[6:0] ? phv_data_33 : _GEN_2104; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2106 = 7'h22 == total_offset_36[6:0] ? phv_data_34 : _GEN_2105; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2107 = 7'h23 == total_offset_36[6:0] ? phv_data_35 : _GEN_2106; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2108 = 7'h24 == total_offset_36[6:0] ? phv_data_36 : _GEN_2107; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2109 = 7'h25 == total_offset_36[6:0] ? phv_data_37 : _GEN_2108; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2110 = 7'h26 == total_offset_36[6:0] ? phv_data_38 : _GEN_2109; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2111 = 7'h27 == total_offset_36[6:0] ? phv_data_39 : _GEN_2110; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2112 = 7'h28 == total_offset_36[6:0] ? phv_data_40 : _GEN_2111; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2113 = 7'h29 == total_offset_36[6:0] ? phv_data_41 : _GEN_2112; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2114 = 7'h2a == total_offset_36[6:0] ? phv_data_42 : _GEN_2113; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2115 = 7'h2b == total_offset_36[6:0] ? phv_data_43 : _GEN_2114; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2116 = 7'h2c == total_offset_36[6:0] ? phv_data_44 : _GEN_2115; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2117 = 7'h2d == total_offset_36[6:0] ? phv_data_45 : _GEN_2116; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2118 = 7'h2e == total_offset_36[6:0] ? phv_data_46 : _GEN_2117; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2119 = 7'h2f == total_offset_36[6:0] ? phv_data_47 : _GEN_2118; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2120 = 7'h30 == total_offset_36[6:0] ? phv_data_48 : _GEN_2119; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2121 = 7'h31 == total_offset_36[6:0] ? phv_data_49 : _GEN_2120; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2122 = 7'h32 == total_offset_36[6:0] ? phv_data_50 : _GEN_2121; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2123 = 7'h33 == total_offset_36[6:0] ? phv_data_51 : _GEN_2122; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2124 = 7'h34 == total_offset_36[6:0] ? phv_data_52 : _GEN_2123; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2125 = 7'h35 == total_offset_36[6:0] ? phv_data_53 : _GEN_2124; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2126 = 7'h36 == total_offset_36[6:0] ? phv_data_54 : _GEN_2125; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2127 = 7'h37 == total_offset_36[6:0] ? phv_data_55 : _GEN_2126; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2128 = 7'h38 == total_offset_36[6:0] ? phv_data_56 : _GEN_2127; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2129 = 7'h39 == total_offset_36[6:0] ? phv_data_57 : _GEN_2128; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2130 = 7'h3a == total_offset_36[6:0] ? phv_data_58 : _GEN_2129; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2131 = 7'h3b == total_offset_36[6:0] ? phv_data_59 : _GEN_2130; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2132 = 7'h3c == total_offset_36[6:0] ? phv_data_60 : _GEN_2131; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2133 = 7'h3d == total_offset_36[6:0] ? phv_data_61 : _GEN_2132; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2134 = 7'h3e == total_offset_36[6:0] ? phv_data_62 : _GEN_2133; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2135 = 7'h3f == total_offset_36[6:0] ? phv_data_63 : _GEN_2134; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2136 = 7'h40 == total_offset_36[6:0] ? phv_data_64 : _GEN_2135; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2137 = 7'h41 == total_offset_36[6:0] ? phv_data_65 : _GEN_2136; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2138 = 7'h42 == total_offset_36[6:0] ? phv_data_66 : _GEN_2137; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2139 = 7'h43 == total_offset_36[6:0] ? phv_data_67 : _GEN_2138; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2140 = 7'h44 == total_offset_36[6:0] ? phv_data_68 : _GEN_2139; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2141 = 7'h45 == total_offset_36[6:0] ? phv_data_69 : _GEN_2140; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2142 = 7'h46 == total_offset_36[6:0] ? phv_data_70 : _GEN_2141; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2143 = 7'h47 == total_offset_36[6:0] ? phv_data_71 : _GEN_2142; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2144 = 7'h48 == total_offset_36[6:0] ? phv_data_72 : _GEN_2143; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2145 = 7'h49 == total_offset_36[6:0] ? phv_data_73 : _GEN_2144; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2146 = 7'h4a == total_offset_36[6:0] ? phv_data_74 : _GEN_2145; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2147 = 7'h4b == total_offset_36[6:0] ? phv_data_75 : _GEN_2146; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2148 = 7'h4c == total_offset_36[6:0] ? phv_data_76 : _GEN_2147; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2149 = 7'h4d == total_offset_36[6:0] ? phv_data_77 : _GEN_2148; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2150 = 7'h4e == total_offset_36[6:0] ? phv_data_78 : _GEN_2149; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2151 = 7'h4f == total_offset_36[6:0] ? phv_data_79 : _GEN_2150; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2152 = 7'h50 == total_offset_36[6:0] ? phv_data_80 : _GEN_2151; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2153 = 7'h51 == total_offset_36[6:0] ? phv_data_81 : _GEN_2152; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2154 = 7'h52 == total_offset_36[6:0] ? phv_data_82 : _GEN_2153; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2155 = 7'h53 == total_offset_36[6:0] ? phv_data_83 : _GEN_2154; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2156 = 7'h54 == total_offset_36[6:0] ? phv_data_84 : _GEN_2155; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2157 = 7'h55 == total_offset_36[6:0] ? phv_data_85 : _GEN_2156; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2158 = 7'h56 == total_offset_36[6:0] ? phv_data_86 : _GEN_2157; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2159 = 7'h57 == total_offset_36[6:0] ? phv_data_87 : _GEN_2158; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2160 = 7'h58 == total_offset_36[6:0] ? phv_data_88 : _GEN_2159; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2161 = 7'h59 == total_offset_36[6:0] ? phv_data_89 : _GEN_2160; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2162 = 7'h5a == total_offset_36[6:0] ? phv_data_90 : _GEN_2161; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2163 = 7'h5b == total_offset_36[6:0] ? phv_data_91 : _GEN_2162; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2164 = 7'h5c == total_offset_36[6:0] ? phv_data_92 : _GEN_2163; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2165 = 7'h5d == total_offset_36[6:0] ? phv_data_93 : _GEN_2164; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2166 = 7'h5e == total_offset_36[6:0] ? phv_data_94 : _GEN_2165; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2167 = 7'h5f == total_offset_36[6:0] ? phv_data_95 : _GEN_2166; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_4 = 8'h4 < length_2 ? _GEN_2167 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_37 = offset_2 + 8'h5; // @[executor.scala 148:53]
  wire [7:0] _GEN_2170 = 7'h1 == total_offset_37[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2171 = 7'h2 == total_offset_37[6:0] ? phv_data_2 : _GEN_2170; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2172 = 7'h3 == total_offset_37[6:0] ? phv_data_3 : _GEN_2171; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2173 = 7'h4 == total_offset_37[6:0] ? phv_data_4 : _GEN_2172; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2174 = 7'h5 == total_offset_37[6:0] ? phv_data_5 : _GEN_2173; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2175 = 7'h6 == total_offset_37[6:0] ? phv_data_6 : _GEN_2174; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2176 = 7'h7 == total_offset_37[6:0] ? phv_data_7 : _GEN_2175; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2177 = 7'h8 == total_offset_37[6:0] ? phv_data_8 : _GEN_2176; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2178 = 7'h9 == total_offset_37[6:0] ? phv_data_9 : _GEN_2177; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2179 = 7'ha == total_offset_37[6:0] ? phv_data_10 : _GEN_2178; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2180 = 7'hb == total_offset_37[6:0] ? phv_data_11 : _GEN_2179; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2181 = 7'hc == total_offset_37[6:0] ? phv_data_12 : _GEN_2180; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2182 = 7'hd == total_offset_37[6:0] ? phv_data_13 : _GEN_2181; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2183 = 7'he == total_offset_37[6:0] ? phv_data_14 : _GEN_2182; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2184 = 7'hf == total_offset_37[6:0] ? phv_data_15 : _GEN_2183; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2185 = 7'h10 == total_offset_37[6:0] ? phv_data_16 : _GEN_2184; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2186 = 7'h11 == total_offset_37[6:0] ? phv_data_17 : _GEN_2185; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2187 = 7'h12 == total_offset_37[6:0] ? phv_data_18 : _GEN_2186; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2188 = 7'h13 == total_offset_37[6:0] ? phv_data_19 : _GEN_2187; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2189 = 7'h14 == total_offset_37[6:0] ? phv_data_20 : _GEN_2188; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2190 = 7'h15 == total_offset_37[6:0] ? phv_data_21 : _GEN_2189; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2191 = 7'h16 == total_offset_37[6:0] ? phv_data_22 : _GEN_2190; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2192 = 7'h17 == total_offset_37[6:0] ? phv_data_23 : _GEN_2191; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2193 = 7'h18 == total_offset_37[6:0] ? phv_data_24 : _GEN_2192; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2194 = 7'h19 == total_offset_37[6:0] ? phv_data_25 : _GEN_2193; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2195 = 7'h1a == total_offset_37[6:0] ? phv_data_26 : _GEN_2194; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2196 = 7'h1b == total_offset_37[6:0] ? phv_data_27 : _GEN_2195; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2197 = 7'h1c == total_offset_37[6:0] ? phv_data_28 : _GEN_2196; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2198 = 7'h1d == total_offset_37[6:0] ? phv_data_29 : _GEN_2197; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2199 = 7'h1e == total_offset_37[6:0] ? phv_data_30 : _GEN_2198; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2200 = 7'h1f == total_offset_37[6:0] ? phv_data_31 : _GEN_2199; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2201 = 7'h20 == total_offset_37[6:0] ? phv_data_32 : _GEN_2200; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2202 = 7'h21 == total_offset_37[6:0] ? phv_data_33 : _GEN_2201; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2203 = 7'h22 == total_offset_37[6:0] ? phv_data_34 : _GEN_2202; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2204 = 7'h23 == total_offset_37[6:0] ? phv_data_35 : _GEN_2203; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2205 = 7'h24 == total_offset_37[6:0] ? phv_data_36 : _GEN_2204; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2206 = 7'h25 == total_offset_37[6:0] ? phv_data_37 : _GEN_2205; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2207 = 7'h26 == total_offset_37[6:0] ? phv_data_38 : _GEN_2206; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2208 = 7'h27 == total_offset_37[6:0] ? phv_data_39 : _GEN_2207; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2209 = 7'h28 == total_offset_37[6:0] ? phv_data_40 : _GEN_2208; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2210 = 7'h29 == total_offset_37[6:0] ? phv_data_41 : _GEN_2209; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2211 = 7'h2a == total_offset_37[6:0] ? phv_data_42 : _GEN_2210; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2212 = 7'h2b == total_offset_37[6:0] ? phv_data_43 : _GEN_2211; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2213 = 7'h2c == total_offset_37[6:0] ? phv_data_44 : _GEN_2212; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2214 = 7'h2d == total_offset_37[6:0] ? phv_data_45 : _GEN_2213; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2215 = 7'h2e == total_offset_37[6:0] ? phv_data_46 : _GEN_2214; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2216 = 7'h2f == total_offset_37[6:0] ? phv_data_47 : _GEN_2215; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2217 = 7'h30 == total_offset_37[6:0] ? phv_data_48 : _GEN_2216; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2218 = 7'h31 == total_offset_37[6:0] ? phv_data_49 : _GEN_2217; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2219 = 7'h32 == total_offset_37[6:0] ? phv_data_50 : _GEN_2218; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2220 = 7'h33 == total_offset_37[6:0] ? phv_data_51 : _GEN_2219; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2221 = 7'h34 == total_offset_37[6:0] ? phv_data_52 : _GEN_2220; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2222 = 7'h35 == total_offset_37[6:0] ? phv_data_53 : _GEN_2221; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2223 = 7'h36 == total_offset_37[6:0] ? phv_data_54 : _GEN_2222; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2224 = 7'h37 == total_offset_37[6:0] ? phv_data_55 : _GEN_2223; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2225 = 7'h38 == total_offset_37[6:0] ? phv_data_56 : _GEN_2224; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2226 = 7'h39 == total_offset_37[6:0] ? phv_data_57 : _GEN_2225; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2227 = 7'h3a == total_offset_37[6:0] ? phv_data_58 : _GEN_2226; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2228 = 7'h3b == total_offset_37[6:0] ? phv_data_59 : _GEN_2227; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2229 = 7'h3c == total_offset_37[6:0] ? phv_data_60 : _GEN_2228; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2230 = 7'h3d == total_offset_37[6:0] ? phv_data_61 : _GEN_2229; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2231 = 7'h3e == total_offset_37[6:0] ? phv_data_62 : _GEN_2230; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2232 = 7'h3f == total_offset_37[6:0] ? phv_data_63 : _GEN_2231; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2233 = 7'h40 == total_offset_37[6:0] ? phv_data_64 : _GEN_2232; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2234 = 7'h41 == total_offset_37[6:0] ? phv_data_65 : _GEN_2233; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2235 = 7'h42 == total_offset_37[6:0] ? phv_data_66 : _GEN_2234; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2236 = 7'h43 == total_offset_37[6:0] ? phv_data_67 : _GEN_2235; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2237 = 7'h44 == total_offset_37[6:0] ? phv_data_68 : _GEN_2236; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2238 = 7'h45 == total_offset_37[6:0] ? phv_data_69 : _GEN_2237; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2239 = 7'h46 == total_offset_37[6:0] ? phv_data_70 : _GEN_2238; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2240 = 7'h47 == total_offset_37[6:0] ? phv_data_71 : _GEN_2239; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2241 = 7'h48 == total_offset_37[6:0] ? phv_data_72 : _GEN_2240; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2242 = 7'h49 == total_offset_37[6:0] ? phv_data_73 : _GEN_2241; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2243 = 7'h4a == total_offset_37[6:0] ? phv_data_74 : _GEN_2242; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2244 = 7'h4b == total_offset_37[6:0] ? phv_data_75 : _GEN_2243; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2245 = 7'h4c == total_offset_37[6:0] ? phv_data_76 : _GEN_2244; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2246 = 7'h4d == total_offset_37[6:0] ? phv_data_77 : _GEN_2245; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2247 = 7'h4e == total_offset_37[6:0] ? phv_data_78 : _GEN_2246; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2248 = 7'h4f == total_offset_37[6:0] ? phv_data_79 : _GEN_2247; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2249 = 7'h50 == total_offset_37[6:0] ? phv_data_80 : _GEN_2248; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2250 = 7'h51 == total_offset_37[6:0] ? phv_data_81 : _GEN_2249; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2251 = 7'h52 == total_offset_37[6:0] ? phv_data_82 : _GEN_2250; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2252 = 7'h53 == total_offset_37[6:0] ? phv_data_83 : _GEN_2251; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2253 = 7'h54 == total_offset_37[6:0] ? phv_data_84 : _GEN_2252; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2254 = 7'h55 == total_offset_37[6:0] ? phv_data_85 : _GEN_2253; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2255 = 7'h56 == total_offset_37[6:0] ? phv_data_86 : _GEN_2254; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2256 = 7'h57 == total_offset_37[6:0] ? phv_data_87 : _GEN_2255; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2257 = 7'h58 == total_offset_37[6:0] ? phv_data_88 : _GEN_2256; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2258 = 7'h59 == total_offset_37[6:0] ? phv_data_89 : _GEN_2257; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2259 = 7'h5a == total_offset_37[6:0] ? phv_data_90 : _GEN_2258; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2260 = 7'h5b == total_offset_37[6:0] ? phv_data_91 : _GEN_2259; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2261 = 7'h5c == total_offset_37[6:0] ? phv_data_92 : _GEN_2260; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2262 = 7'h5d == total_offset_37[6:0] ? phv_data_93 : _GEN_2261; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2263 = 7'h5e == total_offset_37[6:0] ? phv_data_94 : _GEN_2262; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2264 = 7'h5f == total_offset_37[6:0] ? phv_data_95 : _GEN_2263; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_5 = 8'h5 < length_2 ? _GEN_2264 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_38 = offset_2 + 8'h6; // @[executor.scala 148:53]
  wire [7:0] _GEN_2267 = 7'h1 == total_offset_38[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2268 = 7'h2 == total_offset_38[6:0] ? phv_data_2 : _GEN_2267; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2269 = 7'h3 == total_offset_38[6:0] ? phv_data_3 : _GEN_2268; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2270 = 7'h4 == total_offset_38[6:0] ? phv_data_4 : _GEN_2269; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2271 = 7'h5 == total_offset_38[6:0] ? phv_data_5 : _GEN_2270; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2272 = 7'h6 == total_offset_38[6:0] ? phv_data_6 : _GEN_2271; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2273 = 7'h7 == total_offset_38[6:0] ? phv_data_7 : _GEN_2272; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2274 = 7'h8 == total_offset_38[6:0] ? phv_data_8 : _GEN_2273; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2275 = 7'h9 == total_offset_38[6:0] ? phv_data_9 : _GEN_2274; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2276 = 7'ha == total_offset_38[6:0] ? phv_data_10 : _GEN_2275; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2277 = 7'hb == total_offset_38[6:0] ? phv_data_11 : _GEN_2276; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2278 = 7'hc == total_offset_38[6:0] ? phv_data_12 : _GEN_2277; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2279 = 7'hd == total_offset_38[6:0] ? phv_data_13 : _GEN_2278; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2280 = 7'he == total_offset_38[6:0] ? phv_data_14 : _GEN_2279; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2281 = 7'hf == total_offset_38[6:0] ? phv_data_15 : _GEN_2280; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2282 = 7'h10 == total_offset_38[6:0] ? phv_data_16 : _GEN_2281; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2283 = 7'h11 == total_offset_38[6:0] ? phv_data_17 : _GEN_2282; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2284 = 7'h12 == total_offset_38[6:0] ? phv_data_18 : _GEN_2283; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2285 = 7'h13 == total_offset_38[6:0] ? phv_data_19 : _GEN_2284; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2286 = 7'h14 == total_offset_38[6:0] ? phv_data_20 : _GEN_2285; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2287 = 7'h15 == total_offset_38[6:0] ? phv_data_21 : _GEN_2286; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2288 = 7'h16 == total_offset_38[6:0] ? phv_data_22 : _GEN_2287; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2289 = 7'h17 == total_offset_38[6:0] ? phv_data_23 : _GEN_2288; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2290 = 7'h18 == total_offset_38[6:0] ? phv_data_24 : _GEN_2289; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2291 = 7'h19 == total_offset_38[6:0] ? phv_data_25 : _GEN_2290; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2292 = 7'h1a == total_offset_38[6:0] ? phv_data_26 : _GEN_2291; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2293 = 7'h1b == total_offset_38[6:0] ? phv_data_27 : _GEN_2292; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2294 = 7'h1c == total_offset_38[6:0] ? phv_data_28 : _GEN_2293; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2295 = 7'h1d == total_offset_38[6:0] ? phv_data_29 : _GEN_2294; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2296 = 7'h1e == total_offset_38[6:0] ? phv_data_30 : _GEN_2295; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2297 = 7'h1f == total_offset_38[6:0] ? phv_data_31 : _GEN_2296; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2298 = 7'h20 == total_offset_38[6:0] ? phv_data_32 : _GEN_2297; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2299 = 7'h21 == total_offset_38[6:0] ? phv_data_33 : _GEN_2298; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2300 = 7'h22 == total_offset_38[6:0] ? phv_data_34 : _GEN_2299; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2301 = 7'h23 == total_offset_38[6:0] ? phv_data_35 : _GEN_2300; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2302 = 7'h24 == total_offset_38[6:0] ? phv_data_36 : _GEN_2301; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2303 = 7'h25 == total_offset_38[6:0] ? phv_data_37 : _GEN_2302; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2304 = 7'h26 == total_offset_38[6:0] ? phv_data_38 : _GEN_2303; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2305 = 7'h27 == total_offset_38[6:0] ? phv_data_39 : _GEN_2304; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2306 = 7'h28 == total_offset_38[6:0] ? phv_data_40 : _GEN_2305; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2307 = 7'h29 == total_offset_38[6:0] ? phv_data_41 : _GEN_2306; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2308 = 7'h2a == total_offset_38[6:0] ? phv_data_42 : _GEN_2307; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2309 = 7'h2b == total_offset_38[6:0] ? phv_data_43 : _GEN_2308; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2310 = 7'h2c == total_offset_38[6:0] ? phv_data_44 : _GEN_2309; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2311 = 7'h2d == total_offset_38[6:0] ? phv_data_45 : _GEN_2310; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2312 = 7'h2e == total_offset_38[6:0] ? phv_data_46 : _GEN_2311; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2313 = 7'h2f == total_offset_38[6:0] ? phv_data_47 : _GEN_2312; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2314 = 7'h30 == total_offset_38[6:0] ? phv_data_48 : _GEN_2313; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2315 = 7'h31 == total_offset_38[6:0] ? phv_data_49 : _GEN_2314; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2316 = 7'h32 == total_offset_38[6:0] ? phv_data_50 : _GEN_2315; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2317 = 7'h33 == total_offset_38[6:0] ? phv_data_51 : _GEN_2316; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2318 = 7'h34 == total_offset_38[6:0] ? phv_data_52 : _GEN_2317; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2319 = 7'h35 == total_offset_38[6:0] ? phv_data_53 : _GEN_2318; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2320 = 7'h36 == total_offset_38[6:0] ? phv_data_54 : _GEN_2319; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2321 = 7'h37 == total_offset_38[6:0] ? phv_data_55 : _GEN_2320; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2322 = 7'h38 == total_offset_38[6:0] ? phv_data_56 : _GEN_2321; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2323 = 7'h39 == total_offset_38[6:0] ? phv_data_57 : _GEN_2322; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2324 = 7'h3a == total_offset_38[6:0] ? phv_data_58 : _GEN_2323; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2325 = 7'h3b == total_offset_38[6:0] ? phv_data_59 : _GEN_2324; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2326 = 7'h3c == total_offset_38[6:0] ? phv_data_60 : _GEN_2325; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2327 = 7'h3d == total_offset_38[6:0] ? phv_data_61 : _GEN_2326; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2328 = 7'h3e == total_offset_38[6:0] ? phv_data_62 : _GEN_2327; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2329 = 7'h3f == total_offset_38[6:0] ? phv_data_63 : _GEN_2328; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2330 = 7'h40 == total_offset_38[6:0] ? phv_data_64 : _GEN_2329; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2331 = 7'h41 == total_offset_38[6:0] ? phv_data_65 : _GEN_2330; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2332 = 7'h42 == total_offset_38[6:0] ? phv_data_66 : _GEN_2331; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2333 = 7'h43 == total_offset_38[6:0] ? phv_data_67 : _GEN_2332; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2334 = 7'h44 == total_offset_38[6:0] ? phv_data_68 : _GEN_2333; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2335 = 7'h45 == total_offset_38[6:0] ? phv_data_69 : _GEN_2334; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2336 = 7'h46 == total_offset_38[6:0] ? phv_data_70 : _GEN_2335; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2337 = 7'h47 == total_offset_38[6:0] ? phv_data_71 : _GEN_2336; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2338 = 7'h48 == total_offset_38[6:0] ? phv_data_72 : _GEN_2337; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2339 = 7'h49 == total_offset_38[6:0] ? phv_data_73 : _GEN_2338; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2340 = 7'h4a == total_offset_38[6:0] ? phv_data_74 : _GEN_2339; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2341 = 7'h4b == total_offset_38[6:0] ? phv_data_75 : _GEN_2340; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2342 = 7'h4c == total_offset_38[6:0] ? phv_data_76 : _GEN_2341; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2343 = 7'h4d == total_offset_38[6:0] ? phv_data_77 : _GEN_2342; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2344 = 7'h4e == total_offset_38[6:0] ? phv_data_78 : _GEN_2343; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2345 = 7'h4f == total_offset_38[6:0] ? phv_data_79 : _GEN_2344; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2346 = 7'h50 == total_offset_38[6:0] ? phv_data_80 : _GEN_2345; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2347 = 7'h51 == total_offset_38[6:0] ? phv_data_81 : _GEN_2346; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2348 = 7'h52 == total_offset_38[6:0] ? phv_data_82 : _GEN_2347; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2349 = 7'h53 == total_offset_38[6:0] ? phv_data_83 : _GEN_2348; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2350 = 7'h54 == total_offset_38[6:0] ? phv_data_84 : _GEN_2349; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2351 = 7'h55 == total_offset_38[6:0] ? phv_data_85 : _GEN_2350; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2352 = 7'h56 == total_offset_38[6:0] ? phv_data_86 : _GEN_2351; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2353 = 7'h57 == total_offset_38[6:0] ? phv_data_87 : _GEN_2352; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2354 = 7'h58 == total_offset_38[6:0] ? phv_data_88 : _GEN_2353; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2355 = 7'h59 == total_offset_38[6:0] ? phv_data_89 : _GEN_2354; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2356 = 7'h5a == total_offset_38[6:0] ? phv_data_90 : _GEN_2355; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2357 = 7'h5b == total_offset_38[6:0] ? phv_data_91 : _GEN_2356; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2358 = 7'h5c == total_offset_38[6:0] ? phv_data_92 : _GEN_2357; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2359 = 7'h5d == total_offset_38[6:0] ? phv_data_93 : _GEN_2358; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2360 = 7'h5e == total_offset_38[6:0] ? phv_data_94 : _GEN_2359; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2361 = 7'h5f == total_offset_38[6:0] ? phv_data_95 : _GEN_2360; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_6 = 8'h6 < length_2 ? _GEN_2361 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_39 = offset_2 + 8'h7; // @[executor.scala 148:53]
  wire [7:0] _GEN_2364 = 7'h1 == total_offset_39[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2365 = 7'h2 == total_offset_39[6:0] ? phv_data_2 : _GEN_2364; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2366 = 7'h3 == total_offset_39[6:0] ? phv_data_3 : _GEN_2365; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2367 = 7'h4 == total_offset_39[6:0] ? phv_data_4 : _GEN_2366; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2368 = 7'h5 == total_offset_39[6:0] ? phv_data_5 : _GEN_2367; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2369 = 7'h6 == total_offset_39[6:0] ? phv_data_6 : _GEN_2368; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2370 = 7'h7 == total_offset_39[6:0] ? phv_data_7 : _GEN_2369; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2371 = 7'h8 == total_offset_39[6:0] ? phv_data_8 : _GEN_2370; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2372 = 7'h9 == total_offset_39[6:0] ? phv_data_9 : _GEN_2371; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2373 = 7'ha == total_offset_39[6:0] ? phv_data_10 : _GEN_2372; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2374 = 7'hb == total_offset_39[6:0] ? phv_data_11 : _GEN_2373; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2375 = 7'hc == total_offset_39[6:0] ? phv_data_12 : _GEN_2374; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2376 = 7'hd == total_offset_39[6:0] ? phv_data_13 : _GEN_2375; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2377 = 7'he == total_offset_39[6:0] ? phv_data_14 : _GEN_2376; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2378 = 7'hf == total_offset_39[6:0] ? phv_data_15 : _GEN_2377; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2379 = 7'h10 == total_offset_39[6:0] ? phv_data_16 : _GEN_2378; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2380 = 7'h11 == total_offset_39[6:0] ? phv_data_17 : _GEN_2379; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2381 = 7'h12 == total_offset_39[6:0] ? phv_data_18 : _GEN_2380; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2382 = 7'h13 == total_offset_39[6:0] ? phv_data_19 : _GEN_2381; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2383 = 7'h14 == total_offset_39[6:0] ? phv_data_20 : _GEN_2382; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2384 = 7'h15 == total_offset_39[6:0] ? phv_data_21 : _GEN_2383; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2385 = 7'h16 == total_offset_39[6:0] ? phv_data_22 : _GEN_2384; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2386 = 7'h17 == total_offset_39[6:0] ? phv_data_23 : _GEN_2385; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2387 = 7'h18 == total_offset_39[6:0] ? phv_data_24 : _GEN_2386; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2388 = 7'h19 == total_offset_39[6:0] ? phv_data_25 : _GEN_2387; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2389 = 7'h1a == total_offset_39[6:0] ? phv_data_26 : _GEN_2388; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2390 = 7'h1b == total_offset_39[6:0] ? phv_data_27 : _GEN_2389; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2391 = 7'h1c == total_offset_39[6:0] ? phv_data_28 : _GEN_2390; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2392 = 7'h1d == total_offset_39[6:0] ? phv_data_29 : _GEN_2391; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2393 = 7'h1e == total_offset_39[6:0] ? phv_data_30 : _GEN_2392; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2394 = 7'h1f == total_offset_39[6:0] ? phv_data_31 : _GEN_2393; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2395 = 7'h20 == total_offset_39[6:0] ? phv_data_32 : _GEN_2394; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2396 = 7'h21 == total_offset_39[6:0] ? phv_data_33 : _GEN_2395; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2397 = 7'h22 == total_offset_39[6:0] ? phv_data_34 : _GEN_2396; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2398 = 7'h23 == total_offset_39[6:0] ? phv_data_35 : _GEN_2397; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2399 = 7'h24 == total_offset_39[6:0] ? phv_data_36 : _GEN_2398; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2400 = 7'h25 == total_offset_39[6:0] ? phv_data_37 : _GEN_2399; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2401 = 7'h26 == total_offset_39[6:0] ? phv_data_38 : _GEN_2400; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2402 = 7'h27 == total_offset_39[6:0] ? phv_data_39 : _GEN_2401; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2403 = 7'h28 == total_offset_39[6:0] ? phv_data_40 : _GEN_2402; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2404 = 7'h29 == total_offset_39[6:0] ? phv_data_41 : _GEN_2403; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2405 = 7'h2a == total_offset_39[6:0] ? phv_data_42 : _GEN_2404; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2406 = 7'h2b == total_offset_39[6:0] ? phv_data_43 : _GEN_2405; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2407 = 7'h2c == total_offset_39[6:0] ? phv_data_44 : _GEN_2406; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2408 = 7'h2d == total_offset_39[6:0] ? phv_data_45 : _GEN_2407; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2409 = 7'h2e == total_offset_39[6:0] ? phv_data_46 : _GEN_2408; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2410 = 7'h2f == total_offset_39[6:0] ? phv_data_47 : _GEN_2409; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2411 = 7'h30 == total_offset_39[6:0] ? phv_data_48 : _GEN_2410; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2412 = 7'h31 == total_offset_39[6:0] ? phv_data_49 : _GEN_2411; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2413 = 7'h32 == total_offset_39[6:0] ? phv_data_50 : _GEN_2412; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2414 = 7'h33 == total_offset_39[6:0] ? phv_data_51 : _GEN_2413; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2415 = 7'h34 == total_offset_39[6:0] ? phv_data_52 : _GEN_2414; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2416 = 7'h35 == total_offset_39[6:0] ? phv_data_53 : _GEN_2415; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2417 = 7'h36 == total_offset_39[6:0] ? phv_data_54 : _GEN_2416; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2418 = 7'h37 == total_offset_39[6:0] ? phv_data_55 : _GEN_2417; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2419 = 7'h38 == total_offset_39[6:0] ? phv_data_56 : _GEN_2418; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2420 = 7'h39 == total_offset_39[6:0] ? phv_data_57 : _GEN_2419; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2421 = 7'h3a == total_offset_39[6:0] ? phv_data_58 : _GEN_2420; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2422 = 7'h3b == total_offset_39[6:0] ? phv_data_59 : _GEN_2421; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2423 = 7'h3c == total_offset_39[6:0] ? phv_data_60 : _GEN_2422; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2424 = 7'h3d == total_offset_39[6:0] ? phv_data_61 : _GEN_2423; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2425 = 7'h3e == total_offset_39[6:0] ? phv_data_62 : _GEN_2424; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2426 = 7'h3f == total_offset_39[6:0] ? phv_data_63 : _GEN_2425; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2427 = 7'h40 == total_offset_39[6:0] ? phv_data_64 : _GEN_2426; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2428 = 7'h41 == total_offset_39[6:0] ? phv_data_65 : _GEN_2427; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2429 = 7'h42 == total_offset_39[6:0] ? phv_data_66 : _GEN_2428; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2430 = 7'h43 == total_offset_39[6:0] ? phv_data_67 : _GEN_2429; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2431 = 7'h44 == total_offset_39[6:0] ? phv_data_68 : _GEN_2430; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2432 = 7'h45 == total_offset_39[6:0] ? phv_data_69 : _GEN_2431; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2433 = 7'h46 == total_offset_39[6:0] ? phv_data_70 : _GEN_2432; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2434 = 7'h47 == total_offset_39[6:0] ? phv_data_71 : _GEN_2433; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2435 = 7'h48 == total_offset_39[6:0] ? phv_data_72 : _GEN_2434; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2436 = 7'h49 == total_offset_39[6:0] ? phv_data_73 : _GEN_2435; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2437 = 7'h4a == total_offset_39[6:0] ? phv_data_74 : _GEN_2436; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2438 = 7'h4b == total_offset_39[6:0] ? phv_data_75 : _GEN_2437; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2439 = 7'h4c == total_offset_39[6:0] ? phv_data_76 : _GEN_2438; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2440 = 7'h4d == total_offset_39[6:0] ? phv_data_77 : _GEN_2439; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2441 = 7'h4e == total_offset_39[6:0] ? phv_data_78 : _GEN_2440; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2442 = 7'h4f == total_offset_39[6:0] ? phv_data_79 : _GEN_2441; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2443 = 7'h50 == total_offset_39[6:0] ? phv_data_80 : _GEN_2442; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2444 = 7'h51 == total_offset_39[6:0] ? phv_data_81 : _GEN_2443; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2445 = 7'h52 == total_offset_39[6:0] ? phv_data_82 : _GEN_2444; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2446 = 7'h53 == total_offset_39[6:0] ? phv_data_83 : _GEN_2445; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2447 = 7'h54 == total_offset_39[6:0] ? phv_data_84 : _GEN_2446; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2448 = 7'h55 == total_offset_39[6:0] ? phv_data_85 : _GEN_2447; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2449 = 7'h56 == total_offset_39[6:0] ? phv_data_86 : _GEN_2448; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2450 = 7'h57 == total_offset_39[6:0] ? phv_data_87 : _GEN_2449; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2451 = 7'h58 == total_offset_39[6:0] ? phv_data_88 : _GEN_2450; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2452 = 7'h59 == total_offset_39[6:0] ? phv_data_89 : _GEN_2451; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2453 = 7'h5a == total_offset_39[6:0] ? phv_data_90 : _GEN_2452; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2454 = 7'h5b == total_offset_39[6:0] ? phv_data_91 : _GEN_2453; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2455 = 7'h5c == total_offset_39[6:0] ? phv_data_92 : _GEN_2454; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2456 = 7'h5d == total_offset_39[6:0] ? phv_data_93 : _GEN_2455; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2457 = 7'h5e == total_offset_39[6:0] ? phv_data_94 : _GEN_2456; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2458 = 7'h5f == total_offset_39[6:0] ? phv_data_95 : _GEN_2457; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_4_7 = 8'h7 < length_2 ? _GEN_2458 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [63:0] _io_field_out_2_T = {bytes_4_0,bytes_4_1,bytes_4_2,bytes_4_3,bytes_4_4,bytes_4_5,bytes_4_6,bytes_4_7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_2 = io_field_out_2_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length_2 = io_field_out_2_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_40 = {{6'd0}, args_offset_2}; // @[executor.scala 163:56]
  wire [7:0] total_offset_40 = _total_offset_T_40[7:0]; // @[executor.scala 163:56]
  wire [7:0] _GEN_3396 = {{5'd0}, args_length_2}; // @[executor.scala 164:44]
  wire [7:0] _GEN_2461 = 3'h1 == total_offset_40[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2462 = 3'h2 == total_offset_40[2:0] ? args_2 : _GEN_2461; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2463 = 3'h3 == total_offset_40[2:0] ? args_3 : _GEN_2462; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2464 = 3'h4 == total_offset_40[2:0] ? args_4 : _GEN_2463; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2465 = 3'h5 == total_offset_40[2:0] ? args_5 : _GEN_2464; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2466 = 3'h6 == total_offset_40[2:0] ? args_6 : _GEN_2465; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_5_0 = 8'h0 < _GEN_3396 ? _GEN_2466 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] _GEN_3397 = {{5'd0}, args_offset_2}; // @[executor.scala 163:56]
  wire [7:0] total_offset_41 = _GEN_3397 + 8'h1; // @[executor.scala 163:56]
  wire [7:0] _GEN_2469 = 3'h1 == total_offset_41[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2470 = 3'h2 == total_offset_41[2:0] ? args_2 : _GEN_2469; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2471 = 3'h3 == total_offset_41[2:0] ? args_3 : _GEN_2470; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2472 = 3'h4 == total_offset_41[2:0] ? args_4 : _GEN_2471; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2473 = 3'h5 == total_offset_41[2:0] ? args_5 : _GEN_2472; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2474 = 3'h6 == total_offset_41[2:0] ? args_6 : _GEN_2473; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_5_1 = 8'h1 < _GEN_3396 ? _GEN_2474 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_42 = _GEN_3397 + 8'h2; // @[executor.scala 163:56]
  wire [7:0] _GEN_2477 = 3'h1 == total_offset_42[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2478 = 3'h2 == total_offset_42[2:0] ? args_2 : _GEN_2477; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2479 = 3'h3 == total_offset_42[2:0] ? args_3 : _GEN_2478; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2480 = 3'h4 == total_offset_42[2:0] ? args_4 : _GEN_2479; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2481 = 3'h5 == total_offset_42[2:0] ? args_5 : _GEN_2480; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2482 = 3'h6 == total_offset_42[2:0] ? args_6 : _GEN_2481; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_5_2 = 8'h2 < _GEN_3396 ? _GEN_2482 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_43 = _GEN_3397 + 8'h3; // @[executor.scala 163:56]
  wire [7:0] _GEN_2485 = 3'h1 == total_offset_43[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2486 = 3'h2 == total_offset_43[2:0] ? args_2 : _GEN_2485; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2487 = 3'h3 == total_offset_43[2:0] ? args_3 : _GEN_2486; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2488 = 3'h4 == total_offset_43[2:0] ? args_4 : _GEN_2487; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2489 = 3'h5 == total_offset_43[2:0] ? args_5 : _GEN_2488; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2490 = 3'h6 == total_offset_43[2:0] ? args_6 : _GEN_2489; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_5_3 = 8'h3 < _GEN_3396 ? _GEN_2490 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_44 = _GEN_3397 + 8'h4; // @[executor.scala 163:56]
  wire [7:0] _GEN_2493 = 3'h1 == total_offset_44[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2494 = 3'h2 == total_offset_44[2:0] ? args_2 : _GEN_2493; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2495 = 3'h3 == total_offset_44[2:0] ? args_3 : _GEN_2494; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2496 = 3'h4 == total_offset_44[2:0] ? args_4 : _GEN_2495; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2497 = 3'h5 == total_offset_44[2:0] ? args_5 : _GEN_2496; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2498 = 3'h6 == total_offset_44[2:0] ? args_6 : _GEN_2497; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_5_4 = 8'h4 < _GEN_3396 ? _GEN_2498 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_45 = _GEN_3397 + 8'h5; // @[executor.scala 163:56]
  wire [7:0] _GEN_2501 = 3'h1 == total_offset_45[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2502 = 3'h2 == total_offset_45[2:0] ? args_2 : _GEN_2501; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2503 = 3'h3 == total_offset_45[2:0] ? args_3 : _GEN_2502; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2504 = 3'h4 == total_offset_45[2:0] ? args_4 : _GEN_2503; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2505 = 3'h5 == total_offset_45[2:0] ? args_5 : _GEN_2504; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2506 = 3'h6 == total_offset_45[2:0] ? args_6 : _GEN_2505; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_5_5 = 8'h5 < _GEN_3396 ? _GEN_2506 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_46 = _GEN_3397 + 8'h6; // @[executor.scala 163:56]
  wire [7:0] _GEN_2509 = 3'h1 == total_offset_46[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2510 = 3'h2 == total_offset_46[2:0] ? args_2 : _GEN_2509; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2511 = 3'h3 == total_offset_46[2:0] ? args_3 : _GEN_2510; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2512 = 3'h4 == total_offset_46[2:0] ? args_4 : _GEN_2511; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2513 = 3'h5 == total_offset_46[2:0] ? args_5 : _GEN_2512; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_2514 = 3'h6 == total_offset_46[2:0] ? args_6 : _GEN_2513; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_5_6 = 8'h6 < _GEN_3396 ? _GEN_2514 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [63:0] _io_field_out_2_T_1 = {bytes_5_0,bytes_5_1,bytes_5_2,bytes_5_3,bytes_5_4,bytes_5_5,bytes_5_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_2_hi_12 = io_field_out_2_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_2_T_4 = {io_field_out_2_hi_12,io_field_out_2_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_2524 = 4'ha == opcode_2 ? _io_field_out_2_T_1 : _io_field_out_2_T_4; // @[executor.scala 157:51 executor.scala 170:37 executor.scala 173:37]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_3_lo = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire  from_header_3 = length_3 != 8'h0; // @[executor.scala 141:41]
  wire [8:0] _total_offset_T_48 = {{1'd0}, offset_3}; // @[executor.scala 148:53]
  wire [7:0] total_offset_48 = _total_offset_T_48[7:0]; // @[executor.scala 148:53]
  wire [7:0] _GEN_2527 = 7'h1 == total_offset_48[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2528 = 7'h2 == total_offset_48[6:0] ? phv_data_2 : _GEN_2527; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2529 = 7'h3 == total_offset_48[6:0] ? phv_data_3 : _GEN_2528; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2530 = 7'h4 == total_offset_48[6:0] ? phv_data_4 : _GEN_2529; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2531 = 7'h5 == total_offset_48[6:0] ? phv_data_5 : _GEN_2530; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2532 = 7'h6 == total_offset_48[6:0] ? phv_data_6 : _GEN_2531; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2533 = 7'h7 == total_offset_48[6:0] ? phv_data_7 : _GEN_2532; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2534 = 7'h8 == total_offset_48[6:0] ? phv_data_8 : _GEN_2533; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2535 = 7'h9 == total_offset_48[6:0] ? phv_data_9 : _GEN_2534; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2536 = 7'ha == total_offset_48[6:0] ? phv_data_10 : _GEN_2535; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2537 = 7'hb == total_offset_48[6:0] ? phv_data_11 : _GEN_2536; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2538 = 7'hc == total_offset_48[6:0] ? phv_data_12 : _GEN_2537; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2539 = 7'hd == total_offset_48[6:0] ? phv_data_13 : _GEN_2538; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2540 = 7'he == total_offset_48[6:0] ? phv_data_14 : _GEN_2539; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2541 = 7'hf == total_offset_48[6:0] ? phv_data_15 : _GEN_2540; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2542 = 7'h10 == total_offset_48[6:0] ? phv_data_16 : _GEN_2541; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2543 = 7'h11 == total_offset_48[6:0] ? phv_data_17 : _GEN_2542; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2544 = 7'h12 == total_offset_48[6:0] ? phv_data_18 : _GEN_2543; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2545 = 7'h13 == total_offset_48[6:0] ? phv_data_19 : _GEN_2544; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2546 = 7'h14 == total_offset_48[6:0] ? phv_data_20 : _GEN_2545; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2547 = 7'h15 == total_offset_48[6:0] ? phv_data_21 : _GEN_2546; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2548 = 7'h16 == total_offset_48[6:0] ? phv_data_22 : _GEN_2547; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2549 = 7'h17 == total_offset_48[6:0] ? phv_data_23 : _GEN_2548; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2550 = 7'h18 == total_offset_48[6:0] ? phv_data_24 : _GEN_2549; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2551 = 7'h19 == total_offset_48[6:0] ? phv_data_25 : _GEN_2550; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2552 = 7'h1a == total_offset_48[6:0] ? phv_data_26 : _GEN_2551; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2553 = 7'h1b == total_offset_48[6:0] ? phv_data_27 : _GEN_2552; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2554 = 7'h1c == total_offset_48[6:0] ? phv_data_28 : _GEN_2553; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2555 = 7'h1d == total_offset_48[6:0] ? phv_data_29 : _GEN_2554; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2556 = 7'h1e == total_offset_48[6:0] ? phv_data_30 : _GEN_2555; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2557 = 7'h1f == total_offset_48[6:0] ? phv_data_31 : _GEN_2556; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2558 = 7'h20 == total_offset_48[6:0] ? phv_data_32 : _GEN_2557; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2559 = 7'h21 == total_offset_48[6:0] ? phv_data_33 : _GEN_2558; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2560 = 7'h22 == total_offset_48[6:0] ? phv_data_34 : _GEN_2559; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2561 = 7'h23 == total_offset_48[6:0] ? phv_data_35 : _GEN_2560; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2562 = 7'h24 == total_offset_48[6:0] ? phv_data_36 : _GEN_2561; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2563 = 7'h25 == total_offset_48[6:0] ? phv_data_37 : _GEN_2562; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2564 = 7'h26 == total_offset_48[6:0] ? phv_data_38 : _GEN_2563; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2565 = 7'h27 == total_offset_48[6:0] ? phv_data_39 : _GEN_2564; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2566 = 7'h28 == total_offset_48[6:0] ? phv_data_40 : _GEN_2565; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2567 = 7'h29 == total_offset_48[6:0] ? phv_data_41 : _GEN_2566; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2568 = 7'h2a == total_offset_48[6:0] ? phv_data_42 : _GEN_2567; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2569 = 7'h2b == total_offset_48[6:0] ? phv_data_43 : _GEN_2568; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2570 = 7'h2c == total_offset_48[6:0] ? phv_data_44 : _GEN_2569; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2571 = 7'h2d == total_offset_48[6:0] ? phv_data_45 : _GEN_2570; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2572 = 7'h2e == total_offset_48[6:0] ? phv_data_46 : _GEN_2571; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2573 = 7'h2f == total_offset_48[6:0] ? phv_data_47 : _GEN_2572; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2574 = 7'h30 == total_offset_48[6:0] ? phv_data_48 : _GEN_2573; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2575 = 7'h31 == total_offset_48[6:0] ? phv_data_49 : _GEN_2574; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2576 = 7'h32 == total_offset_48[6:0] ? phv_data_50 : _GEN_2575; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2577 = 7'h33 == total_offset_48[6:0] ? phv_data_51 : _GEN_2576; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2578 = 7'h34 == total_offset_48[6:0] ? phv_data_52 : _GEN_2577; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2579 = 7'h35 == total_offset_48[6:0] ? phv_data_53 : _GEN_2578; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2580 = 7'h36 == total_offset_48[6:0] ? phv_data_54 : _GEN_2579; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2581 = 7'h37 == total_offset_48[6:0] ? phv_data_55 : _GEN_2580; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2582 = 7'h38 == total_offset_48[6:0] ? phv_data_56 : _GEN_2581; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2583 = 7'h39 == total_offset_48[6:0] ? phv_data_57 : _GEN_2582; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2584 = 7'h3a == total_offset_48[6:0] ? phv_data_58 : _GEN_2583; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2585 = 7'h3b == total_offset_48[6:0] ? phv_data_59 : _GEN_2584; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2586 = 7'h3c == total_offset_48[6:0] ? phv_data_60 : _GEN_2585; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2587 = 7'h3d == total_offset_48[6:0] ? phv_data_61 : _GEN_2586; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2588 = 7'h3e == total_offset_48[6:0] ? phv_data_62 : _GEN_2587; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2589 = 7'h3f == total_offset_48[6:0] ? phv_data_63 : _GEN_2588; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2590 = 7'h40 == total_offset_48[6:0] ? phv_data_64 : _GEN_2589; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2591 = 7'h41 == total_offset_48[6:0] ? phv_data_65 : _GEN_2590; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2592 = 7'h42 == total_offset_48[6:0] ? phv_data_66 : _GEN_2591; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2593 = 7'h43 == total_offset_48[6:0] ? phv_data_67 : _GEN_2592; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2594 = 7'h44 == total_offset_48[6:0] ? phv_data_68 : _GEN_2593; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2595 = 7'h45 == total_offset_48[6:0] ? phv_data_69 : _GEN_2594; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2596 = 7'h46 == total_offset_48[6:0] ? phv_data_70 : _GEN_2595; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2597 = 7'h47 == total_offset_48[6:0] ? phv_data_71 : _GEN_2596; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2598 = 7'h48 == total_offset_48[6:0] ? phv_data_72 : _GEN_2597; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2599 = 7'h49 == total_offset_48[6:0] ? phv_data_73 : _GEN_2598; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2600 = 7'h4a == total_offset_48[6:0] ? phv_data_74 : _GEN_2599; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2601 = 7'h4b == total_offset_48[6:0] ? phv_data_75 : _GEN_2600; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2602 = 7'h4c == total_offset_48[6:0] ? phv_data_76 : _GEN_2601; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2603 = 7'h4d == total_offset_48[6:0] ? phv_data_77 : _GEN_2602; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2604 = 7'h4e == total_offset_48[6:0] ? phv_data_78 : _GEN_2603; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2605 = 7'h4f == total_offset_48[6:0] ? phv_data_79 : _GEN_2604; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2606 = 7'h50 == total_offset_48[6:0] ? phv_data_80 : _GEN_2605; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2607 = 7'h51 == total_offset_48[6:0] ? phv_data_81 : _GEN_2606; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2608 = 7'h52 == total_offset_48[6:0] ? phv_data_82 : _GEN_2607; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2609 = 7'h53 == total_offset_48[6:0] ? phv_data_83 : _GEN_2608; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2610 = 7'h54 == total_offset_48[6:0] ? phv_data_84 : _GEN_2609; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2611 = 7'h55 == total_offset_48[6:0] ? phv_data_85 : _GEN_2610; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2612 = 7'h56 == total_offset_48[6:0] ? phv_data_86 : _GEN_2611; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2613 = 7'h57 == total_offset_48[6:0] ? phv_data_87 : _GEN_2612; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2614 = 7'h58 == total_offset_48[6:0] ? phv_data_88 : _GEN_2613; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2615 = 7'h59 == total_offset_48[6:0] ? phv_data_89 : _GEN_2614; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2616 = 7'h5a == total_offset_48[6:0] ? phv_data_90 : _GEN_2615; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2617 = 7'h5b == total_offset_48[6:0] ? phv_data_91 : _GEN_2616; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2618 = 7'h5c == total_offset_48[6:0] ? phv_data_92 : _GEN_2617; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2619 = 7'h5d == total_offset_48[6:0] ? phv_data_93 : _GEN_2618; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2620 = 7'h5e == total_offset_48[6:0] ? phv_data_94 : _GEN_2619; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2621 = 7'h5f == total_offset_48[6:0] ? phv_data_95 : _GEN_2620; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_0 = 8'h0 < length_3 ? _GEN_2621 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_49 = offset_3 + 8'h1; // @[executor.scala 148:53]
  wire [7:0] _GEN_2624 = 7'h1 == total_offset_49[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2625 = 7'h2 == total_offset_49[6:0] ? phv_data_2 : _GEN_2624; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2626 = 7'h3 == total_offset_49[6:0] ? phv_data_3 : _GEN_2625; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2627 = 7'h4 == total_offset_49[6:0] ? phv_data_4 : _GEN_2626; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2628 = 7'h5 == total_offset_49[6:0] ? phv_data_5 : _GEN_2627; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2629 = 7'h6 == total_offset_49[6:0] ? phv_data_6 : _GEN_2628; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2630 = 7'h7 == total_offset_49[6:0] ? phv_data_7 : _GEN_2629; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2631 = 7'h8 == total_offset_49[6:0] ? phv_data_8 : _GEN_2630; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2632 = 7'h9 == total_offset_49[6:0] ? phv_data_9 : _GEN_2631; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2633 = 7'ha == total_offset_49[6:0] ? phv_data_10 : _GEN_2632; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2634 = 7'hb == total_offset_49[6:0] ? phv_data_11 : _GEN_2633; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2635 = 7'hc == total_offset_49[6:0] ? phv_data_12 : _GEN_2634; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2636 = 7'hd == total_offset_49[6:0] ? phv_data_13 : _GEN_2635; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2637 = 7'he == total_offset_49[6:0] ? phv_data_14 : _GEN_2636; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2638 = 7'hf == total_offset_49[6:0] ? phv_data_15 : _GEN_2637; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2639 = 7'h10 == total_offset_49[6:0] ? phv_data_16 : _GEN_2638; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2640 = 7'h11 == total_offset_49[6:0] ? phv_data_17 : _GEN_2639; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2641 = 7'h12 == total_offset_49[6:0] ? phv_data_18 : _GEN_2640; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2642 = 7'h13 == total_offset_49[6:0] ? phv_data_19 : _GEN_2641; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2643 = 7'h14 == total_offset_49[6:0] ? phv_data_20 : _GEN_2642; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2644 = 7'h15 == total_offset_49[6:0] ? phv_data_21 : _GEN_2643; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2645 = 7'h16 == total_offset_49[6:0] ? phv_data_22 : _GEN_2644; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2646 = 7'h17 == total_offset_49[6:0] ? phv_data_23 : _GEN_2645; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2647 = 7'h18 == total_offset_49[6:0] ? phv_data_24 : _GEN_2646; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2648 = 7'h19 == total_offset_49[6:0] ? phv_data_25 : _GEN_2647; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2649 = 7'h1a == total_offset_49[6:0] ? phv_data_26 : _GEN_2648; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2650 = 7'h1b == total_offset_49[6:0] ? phv_data_27 : _GEN_2649; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2651 = 7'h1c == total_offset_49[6:0] ? phv_data_28 : _GEN_2650; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2652 = 7'h1d == total_offset_49[6:0] ? phv_data_29 : _GEN_2651; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2653 = 7'h1e == total_offset_49[6:0] ? phv_data_30 : _GEN_2652; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2654 = 7'h1f == total_offset_49[6:0] ? phv_data_31 : _GEN_2653; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2655 = 7'h20 == total_offset_49[6:0] ? phv_data_32 : _GEN_2654; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2656 = 7'h21 == total_offset_49[6:0] ? phv_data_33 : _GEN_2655; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2657 = 7'h22 == total_offset_49[6:0] ? phv_data_34 : _GEN_2656; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2658 = 7'h23 == total_offset_49[6:0] ? phv_data_35 : _GEN_2657; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2659 = 7'h24 == total_offset_49[6:0] ? phv_data_36 : _GEN_2658; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2660 = 7'h25 == total_offset_49[6:0] ? phv_data_37 : _GEN_2659; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2661 = 7'h26 == total_offset_49[6:0] ? phv_data_38 : _GEN_2660; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2662 = 7'h27 == total_offset_49[6:0] ? phv_data_39 : _GEN_2661; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2663 = 7'h28 == total_offset_49[6:0] ? phv_data_40 : _GEN_2662; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2664 = 7'h29 == total_offset_49[6:0] ? phv_data_41 : _GEN_2663; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2665 = 7'h2a == total_offset_49[6:0] ? phv_data_42 : _GEN_2664; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2666 = 7'h2b == total_offset_49[6:0] ? phv_data_43 : _GEN_2665; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2667 = 7'h2c == total_offset_49[6:0] ? phv_data_44 : _GEN_2666; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2668 = 7'h2d == total_offset_49[6:0] ? phv_data_45 : _GEN_2667; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2669 = 7'h2e == total_offset_49[6:0] ? phv_data_46 : _GEN_2668; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2670 = 7'h2f == total_offset_49[6:0] ? phv_data_47 : _GEN_2669; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2671 = 7'h30 == total_offset_49[6:0] ? phv_data_48 : _GEN_2670; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2672 = 7'h31 == total_offset_49[6:0] ? phv_data_49 : _GEN_2671; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2673 = 7'h32 == total_offset_49[6:0] ? phv_data_50 : _GEN_2672; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2674 = 7'h33 == total_offset_49[6:0] ? phv_data_51 : _GEN_2673; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2675 = 7'h34 == total_offset_49[6:0] ? phv_data_52 : _GEN_2674; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2676 = 7'h35 == total_offset_49[6:0] ? phv_data_53 : _GEN_2675; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2677 = 7'h36 == total_offset_49[6:0] ? phv_data_54 : _GEN_2676; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2678 = 7'h37 == total_offset_49[6:0] ? phv_data_55 : _GEN_2677; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2679 = 7'h38 == total_offset_49[6:0] ? phv_data_56 : _GEN_2678; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2680 = 7'h39 == total_offset_49[6:0] ? phv_data_57 : _GEN_2679; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2681 = 7'h3a == total_offset_49[6:0] ? phv_data_58 : _GEN_2680; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2682 = 7'h3b == total_offset_49[6:0] ? phv_data_59 : _GEN_2681; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2683 = 7'h3c == total_offset_49[6:0] ? phv_data_60 : _GEN_2682; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2684 = 7'h3d == total_offset_49[6:0] ? phv_data_61 : _GEN_2683; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2685 = 7'h3e == total_offset_49[6:0] ? phv_data_62 : _GEN_2684; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2686 = 7'h3f == total_offset_49[6:0] ? phv_data_63 : _GEN_2685; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2687 = 7'h40 == total_offset_49[6:0] ? phv_data_64 : _GEN_2686; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2688 = 7'h41 == total_offset_49[6:0] ? phv_data_65 : _GEN_2687; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2689 = 7'h42 == total_offset_49[6:0] ? phv_data_66 : _GEN_2688; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2690 = 7'h43 == total_offset_49[6:0] ? phv_data_67 : _GEN_2689; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2691 = 7'h44 == total_offset_49[6:0] ? phv_data_68 : _GEN_2690; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2692 = 7'h45 == total_offset_49[6:0] ? phv_data_69 : _GEN_2691; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2693 = 7'h46 == total_offset_49[6:0] ? phv_data_70 : _GEN_2692; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2694 = 7'h47 == total_offset_49[6:0] ? phv_data_71 : _GEN_2693; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2695 = 7'h48 == total_offset_49[6:0] ? phv_data_72 : _GEN_2694; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2696 = 7'h49 == total_offset_49[6:0] ? phv_data_73 : _GEN_2695; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2697 = 7'h4a == total_offset_49[6:0] ? phv_data_74 : _GEN_2696; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2698 = 7'h4b == total_offset_49[6:0] ? phv_data_75 : _GEN_2697; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2699 = 7'h4c == total_offset_49[6:0] ? phv_data_76 : _GEN_2698; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2700 = 7'h4d == total_offset_49[6:0] ? phv_data_77 : _GEN_2699; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2701 = 7'h4e == total_offset_49[6:0] ? phv_data_78 : _GEN_2700; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2702 = 7'h4f == total_offset_49[6:0] ? phv_data_79 : _GEN_2701; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2703 = 7'h50 == total_offset_49[6:0] ? phv_data_80 : _GEN_2702; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2704 = 7'h51 == total_offset_49[6:0] ? phv_data_81 : _GEN_2703; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2705 = 7'h52 == total_offset_49[6:0] ? phv_data_82 : _GEN_2704; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2706 = 7'h53 == total_offset_49[6:0] ? phv_data_83 : _GEN_2705; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2707 = 7'h54 == total_offset_49[6:0] ? phv_data_84 : _GEN_2706; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2708 = 7'h55 == total_offset_49[6:0] ? phv_data_85 : _GEN_2707; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2709 = 7'h56 == total_offset_49[6:0] ? phv_data_86 : _GEN_2708; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2710 = 7'h57 == total_offset_49[6:0] ? phv_data_87 : _GEN_2709; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2711 = 7'h58 == total_offset_49[6:0] ? phv_data_88 : _GEN_2710; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2712 = 7'h59 == total_offset_49[6:0] ? phv_data_89 : _GEN_2711; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2713 = 7'h5a == total_offset_49[6:0] ? phv_data_90 : _GEN_2712; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2714 = 7'h5b == total_offset_49[6:0] ? phv_data_91 : _GEN_2713; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2715 = 7'h5c == total_offset_49[6:0] ? phv_data_92 : _GEN_2714; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2716 = 7'h5d == total_offset_49[6:0] ? phv_data_93 : _GEN_2715; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2717 = 7'h5e == total_offset_49[6:0] ? phv_data_94 : _GEN_2716; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2718 = 7'h5f == total_offset_49[6:0] ? phv_data_95 : _GEN_2717; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_1 = 8'h1 < length_3 ? _GEN_2718 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_50 = offset_3 + 8'h2; // @[executor.scala 148:53]
  wire [7:0] _GEN_2721 = 7'h1 == total_offset_50[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2722 = 7'h2 == total_offset_50[6:0] ? phv_data_2 : _GEN_2721; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2723 = 7'h3 == total_offset_50[6:0] ? phv_data_3 : _GEN_2722; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2724 = 7'h4 == total_offset_50[6:0] ? phv_data_4 : _GEN_2723; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2725 = 7'h5 == total_offset_50[6:0] ? phv_data_5 : _GEN_2724; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2726 = 7'h6 == total_offset_50[6:0] ? phv_data_6 : _GEN_2725; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2727 = 7'h7 == total_offset_50[6:0] ? phv_data_7 : _GEN_2726; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2728 = 7'h8 == total_offset_50[6:0] ? phv_data_8 : _GEN_2727; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2729 = 7'h9 == total_offset_50[6:0] ? phv_data_9 : _GEN_2728; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2730 = 7'ha == total_offset_50[6:0] ? phv_data_10 : _GEN_2729; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2731 = 7'hb == total_offset_50[6:0] ? phv_data_11 : _GEN_2730; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2732 = 7'hc == total_offset_50[6:0] ? phv_data_12 : _GEN_2731; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2733 = 7'hd == total_offset_50[6:0] ? phv_data_13 : _GEN_2732; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2734 = 7'he == total_offset_50[6:0] ? phv_data_14 : _GEN_2733; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2735 = 7'hf == total_offset_50[6:0] ? phv_data_15 : _GEN_2734; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2736 = 7'h10 == total_offset_50[6:0] ? phv_data_16 : _GEN_2735; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2737 = 7'h11 == total_offset_50[6:0] ? phv_data_17 : _GEN_2736; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2738 = 7'h12 == total_offset_50[6:0] ? phv_data_18 : _GEN_2737; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2739 = 7'h13 == total_offset_50[6:0] ? phv_data_19 : _GEN_2738; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2740 = 7'h14 == total_offset_50[6:0] ? phv_data_20 : _GEN_2739; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2741 = 7'h15 == total_offset_50[6:0] ? phv_data_21 : _GEN_2740; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2742 = 7'h16 == total_offset_50[6:0] ? phv_data_22 : _GEN_2741; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2743 = 7'h17 == total_offset_50[6:0] ? phv_data_23 : _GEN_2742; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2744 = 7'h18 == total_offset_50[6:0] ? phv_data_24 : _GEN_2743; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2745 = 7'h19 == total_offset_50[6:0] ? phv_data_25 : _GEN_2744; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2746 = 7'h1a == total_offset_50[6:0] ? phv_data_26 : _GEN_2745; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2747 = 7'h1b == total_offset_50[6:0] ? phv_data_27 : _GEN_2746; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2748 = 7'h1c == total_offset_50[6:0] ? phv_data_28 : _GEN_2747; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2749 = 7'h1d == total_offset_50[6:0] ? phv_data_29 : _GEN_2748; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2750 = 7'h1e == total_offset_50[6:0] ? phv_data_30 : _GEN_2749; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2751 = 7'h1f == total_offset_50[6:0] ? phv_data_31 : _GEN_2750; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2752 = 7'h20 == total_offset_50[6:0] ? phv_data_32 : _GEN_2751; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2753 = 7'h21 == total_offset_50[6:0] ? phv_data_33 : _GEN_2752; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2754 = 7'h22 == total_offset_50[6:0] ? phv_data_34 : _GEN_2753; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2755 = 7'h23 == total_offset_50[6:0] ? phv_data_35 : _GEN_2754; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2756 = 7'h24 == total_offset_50[6:0] ? phv_data_36 : _GEN_2755; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2757 = 7'h25 == total_offset_50[6:0] ? phv_data_37 : _GEN_2756; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2758 = 7'h26 == total_offset_50[6:0] ? phv_data_38 : _GEN_2757; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2759 = 7'h27 == total_offset_50[6:0] ? phv_data_39 : _GEN_2758; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2760 = 7'h28 == total_offset_50[6:0] ? phv_data_40 : _GEN_2759; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2761 = 7'h29 == total_offset_50[6:0] ? phv_data_41 : _GEN_2760; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2762 = 7'h2a == total_offset_50[6:0] ? phv_data_42 : _GEN_2761; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2763 = 7'h2b == total_offset_50[6:0] ? phv_data_43 : _GEN_2762; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2764 = 7'h2c == total_offset_50[6:0] ? phv_data_44 : _GEN_2763; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2765 = 7'h2d == total_offset_50[6:0] ? phv_data_45 : _GEN_2764; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2766 = 7'h2e == total_offset_50[6:0] ? phv_data_46 : _GEN_2765; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2767 = 7'h2f == total_offset_50[6:0] ? phv_data_47 : _GEN_2766; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2768 = 7'h30 == total_offset_50[6:0] ? phv_data_48 : _GEN_2767; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2769 = 7'h31 == total_offset_50[6:0] ? phv_data_49 : _GEN_2768; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2770 = 7'h32 == total_offset_50[6:0] ? phv_data_50 : _GEN_2769; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2771 = 7'h33 == total_offset_50[6:0] ? phv_data_51 : _GEN_2770; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2772 = 7'h34 == total_offset_50[6:0] ? phv_data_52 : _GEN_2771; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2773 = 7'h35 == total_offset_50[6:0] ? phv_data_53 : _GEN_2772; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2774 = 7'h36 == total_offset_50[6:0] ? phv_data_54 : _GEN_2773; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2775 = 7'h37 == total_offset_50[6:0] ? phv_data_55 : _GEN_2774; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2776 = 7'h38 == total_offset_50[6:0] ? phv_data_56 : _GEN_2775; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2777 = 7'h39 == total_offset_50[6:0] ? phv_data_57 : _GEN_2776; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2778 = 7'h3a == total_offset_50[6:0] ? phv_data_58 : _GEN_2777; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2779 = 7'h3b == total_offset_50[6:0] ? phv_data_59 : _GEN_2778; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2780 = 7'h3c == total_offset_50[6:0] ? phv_data_60 : _GEN_2779; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2781 = 7'h3d == total_offset_50[6:0] ? phv_data_61 : _GEN_2780; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2782 = 7'h3e == total_offset_50[6:0] ? phv_data_62 : _GEN_2781; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2783 = 7'h3f == total_offset_50[6:0] ? phv_data_63 : _GEN_2782; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2784 = 7'h40 == total_offset_50[6:0] ? phv_data_64 : _GEN_2783; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2785 = 7'h41 == total_offset_50[6:0] ? phv_data_65 : _GEN_2784; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2786 = 7'h42 == total_offset_50[6:0] ? phv_data_66 : _GEN_2785; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2787 = 7'h43 == total_offset_50[6:0] ? phv_data_67 : _GEN_2786; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2788 = 7'h44 == total_offset_50[6:0] ? phv_data_68 : _GEN_2787; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2789 = 7'h45 == total_offset_50[6:0] ? phv_data_69 : _GEN_2788; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2790 = 7'h46 == total_offset_50[6:0] ? phv_data_70 : _GEN_2789; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2791 = 7'h47 == total_offset_50[6:0] ? phv_data_71 : _GEN_2790; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2792 = 7'h48 == total_offset_50[6:0] ? phv_data_72 : _GEN_2791; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2793 = 7'h49 == total_offset_50[6:0] ? phv_data_73 : _GEN_2792; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2794 = 7'h4a == total_offset_50[6:0] ? phv_data_74 : _GEN_2793; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2795 = 7'h4b == total_offset_50[6:0] ? phv_data_75 : _GEN_2794; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2796 = 7'h4c == total_offset_50[6:0] ? phv_data_76 : _GEN_2795; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2797 = 7'h4d == total_offset_50[6:0] ? phv_data_77 : _GEN_2796; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2798 = 7'h4e == total_offset_50[6:0] ? phv_data_78 : _GEN_2797; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2799 = 7'h4f == total_offset_50[6:0] ? phv_data_79 : _GEN_2798; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2800 = 7'h50 == total_offset_50[6:0] ? phv_data_80 : _GEN_2799; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2801 = 7'h51 == total_offset_50[6:0] ? phv_data_81 : _GEN_2800; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2802 = 7'h52 == total_offset_50[6:0] ? phv_data_82 : _GEN_2801; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2803 = 7'h53 == total_offset_50[6:0] ? phv_data_83 : _GEN_2802; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2804 = 7'h54 == total_offset_50[6:0] ? phv_data_84 : _GEN_2803; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2805 = 7'h55 == total_offset_50[6:0] ? phv_data_85 : _GEN_2804; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2806 = 7'h56 == total_offset_50[6:0] ? phv_data_86 : _GEN_2805; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2807 = 7'h57 == total_offset_50[6:0] ? phv_data_87 : _GEN_2806; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2808 = 7'h58 == total_offset_50[6:0] ? phv_data_88 : _GEN_2807; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2809 = 7'h59 == total_offset_50[6:0] ? phv_data_89 : _GEN_2808; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2810 = 7'h5a == total_offset_50[6:0] ? phv_data_90 : _GEN_2809; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2811 = 7'h5b == total_offset_50[6:0] ? phv_data_91 : _GEN_2810; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2812 = 7'h5c == total_offset_50[6:0] ? phv_data_92 : _GEN_2811; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2813 = 7'h5d == total_offset_50[6:0] ? phv_data_93 : _GEN_2812; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2814 = 7'h5e == total_offset_50[6:0] ? phv_data_94 : _GEN_2813; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2815 = 7'h5f == total_offset_50[6:0] ? phv_data_95 : _GEN_2814; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_2 = 8'h2 < length_3 ? _GEN_2815 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_51 = offset_3 + 8'h3; // @[executor.scala 148:53]
  wire [7:0] _GEN_2818 = 7'h1 == total_offset_51[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2819 = 7'h2 == total_offset_51[6:0] ? phv_data_2 : _GEN_2818; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2820 = 7'h3 == total_offset_51[6:0] ? phv_data_3 : _GEN_2819; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2821 = 7'h4 == total_offset_51[6:0] ? phv_data_4 : _GEN_2820; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2822 = 7'h5 == total_offset_51[6:0] ? phv_data_5 : _GEN_2821; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2823 = 7'h6 == total_offset_51[6:0] ? phv_data_6 : _GEN_2822; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2824 = 7'h7 == total_offset_51[6:0] ? phv_data_7 : _GEN_2823; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2825 = 7'h8 == total_offset_51[6:0] ? phv_data_8 : _GEN_2824; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2826 = 7'h9 == total_offset_51[6:0] ? phv_data_9 : _GEN_2825; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2827 = 7'ha == total_offset_51[6:0] ? phv_data_10 : _GEN_2826; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2828 = 7'hb == total_offset_51[6:0] ? phv_data_11 : _GEN_2827; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2829 = 7'hc == total_offset_51[6:0] ? phv_data_12 : _GEN_2828; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2830 = 7'hd == total_offset_51[6:0] ? phv_data_13 : _GEN_2829; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2831 = 7'he == total_offset_51[6:0] ? phv_data_14 : _GEN_2830; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2832 = 7'hf == total_offset_51[6:0] ? phv_data_15 : _GEN_2831; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2833 = 7'h10 == total_offset_51[6:0] ? phv_data_16 : _GEN_2832; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2834 = 7'h11 == total_offset_51[6:0] ? phv_data_17 : _GEN_2833; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2835 = 7'h12 == total_offset_51[6:0] ? phv_data_18 : _GEN_2834; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2836 = 7'h13 == total_offset_51[6:0] ? phv_data_19 : _GEN_2835; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2837 = 7'h14 == total_offset_51[6:0] ? phv_data_20 : _GEN_2836; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2838 = 7'h15 == total_offset_51[6:0] ? phv_data_21 : _GEN_2837; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2839 = 7'h16 == total_offset_51[6:0] ? phv_data_22 : _GEN_2838; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2840 = 7'h17 == total_offset_51[6:0] ? phv_data_23 : _GEN_2839; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2841 = 7'h18 == total_offset_51[6:0] ? phv_data_24 : _GEN_2840; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2842 = 7'h19 == total_offset_51[6:0] ? phv_data_25 : _GEN_2841; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2843 = 7'h1a == total_offset_51[6:0] ? phv_data_26 : _GEN_2842; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2844 = 7'h1b == total_offset_51[6:0] ? phv_data_27 : _GEN_2843; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2845 = 7'h1c == total_offset_51[6:0] ? phv_data_28 : _GEN_2844; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2846 = 7'h1d == total_offset_51[6:0] ? phv_data_29 : _GEN_2845; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2847 = 7'h1e == total_offset_51[6:0] ? phv_data_30 : _GEN_2846; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2848 = 7'h1f == total_offset_51[6:0] ? phv_data_31 : _GEN_2847; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2849 = 7'h20 == total_offset_51[6:0] ? phv_data_32 : _GEN_2848; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2850 = 7'h21 == total_offset_51[6:0] ? phv_data_33 : _GEN_2849; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2851 = 7'h22 == total_offset_51[6:0] ? phv_data_34 : _GEN_2850; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2852 = 7'h23 == total_offset_51[6:0] ? phv_data_35 : _GEN_2851; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2853 = 7'h24 == total_offset_51[6:0] ? phv_data_36 : _GEN_2852; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2854 = 7'h25 == total_offset_51[6:0] ? phv_data_37 : _GEN_2853; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2855 = 7'h26 == total_offset_51[6:0] ? phv_data_38 : _GEN_2854; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2856 = 7'h27 == total_offset_51[6:0] ? phv_data_39 : _GEN_2855; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2857 = 7'h28 == total_offset_51[6:0] ? phv_data_40 : _GEN_2856; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2858 = 7'h29 == total_offset_51[6:0] ? phv_data_41 : _GEN_2857; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2859 = 7'h2a == total_offset_51[6:0] ? phv_data_42 : _GEN_2858; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2860 = 7'h2b == total_offset_51[6:0] ? phv_data_43 : _GEN_2859; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2861 = 7'h2c == total_offset_51[6:0] ? phv_data_44 : _GEN_2860; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2862 = 7'h2d == total_offset_51[6:0] ? phv_data_45 : _GEN_2861; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2863 = 7'h2e == total_offset_51[6:0] ? phv_data_46 : _GEN_2862; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2864 = 7'h2f == total_offset_51[6:0] ? phv_data_47 : _GEN_2863; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2865 = 7'h30 == total_offset_51[6:0] ? phv_data_48 : _GEN_2864; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2866 = 7'h31 == total_offset_51[6:0] ? phv_data_49 : _GEN_2865; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2867 = 7'h32 == total_offset_51[6:0] ? phv_data_50 : _GEN_2866; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2868 = 7'h33 == total_offset_51[6:0] ? phv_data_51 : _GEN_2867; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2869 = 7'h34 == total_offset_51[6:0] ? phv_data_52 : _GEN_2868; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2870 = 7'h35 == total_offset_51[6:0] ? phv_data_53 : _GEN_2869; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2871 = 7'h36 == total_offset_51[6:0] ? phv_data_54 : _GEN_2870; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2872 = 7'h37 == total_offset_51[6:0] ? phv_data_55 : _GEN_2871; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2873 = 7'h38 == total_offset_51[6:0] ? phv_data_56 : _GEN_2872; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2874 = 7'h39 == total_offset_51[6:0] ? phv_data_57 : _GEN_2873; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2875 = 7'h3a == total_offset_51[6:0] ? phv_data_58 : _GEN_2874; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2876 = 7'h3b == total_offset_51[6:0] ? phv_data_59 : _GEN_2875; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2877 = 7'h3c == total_offset_51[6:0] ? phv_data_60 : _GEN_2876; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2878 = 7'h3d == total_offset_51[6:0] ? phv_data_61 : _GEN_2877; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2879 = 7'h3e == total_offset_51[6:0] ? phv_data_62 : _GEN_2878; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2880 = 7'h3f == total_offset_51[6:0] ? phv_data_63 : _GEN_2879; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2881 = 7'h40 == total_offset_51[6:0] ? phv_data_64 : _GEN_2880; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2882 = 7'h41 == total_offset_51[6:0] ? phv_data_65 : _GEN_2881; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2883 = 7'h42 == total_offset_51[6:0] ? phv_data_66 : _GEN_2882; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2884 = 7'h43 == total_offset_51[6:0] ? phv_data_67 : _GEN_2883; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2885 = 7'h44 == total_offset_51[6:0] ? phv_data_68 : _GEN_2884; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2886 = 7'h45 == total_offset_51[6:0] ? phv_data_69 : _GEN_2885; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2887 = 7'h46 == total_offset_51[6:0] ? phv_data_70 : _GEN_2886; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2888 = 7'h47 == total_offset_51[6:0] ? phv_data_71 : _GEN_2887; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2889 = 7'h48 == total_offset_51[6:0] ? phv_data_72 : _GEN_2888; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2890 = 7'h49 == total_offset_51[6:0] ? phv_data_73 : _GEN_2889; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2891 = 7'h4a == total_offset_51[6:0] ? phv_data_74 : _GEN_2890; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2892 = 7'h4b == total_offset_51[6:0] ? phv_data_75 : _GEN_2891; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2893 = 7'h4c == total_offset_51[6:0] ? phv_data_76 : _GEN_2892; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2894 = 7'h4d == total_offset_51[6:0] ? phv_data_77 : _GEN_2893; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2895 = 7'h4e == total_offset_51[6:0] ? phv_data_78 : _GEN_2894; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2896 = 7'h4f == total_offset_51[6:0] ? phv_data_79 : _GEN_2895; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2897 = 7'h50 == total_offset_51[6:0] ? phv_data_80 : _GEN_2896; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2898 = 7'h51 == total_offset_51[6:0] ? phv_data_81 : _GEN_2897; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2899 = 7'h52 == total_offset_51[6:0] ? phv_data_82 : _GEN_2898; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2900 = 7'h53 == total_offset_51[6:0] ? phv_data_83 : _GEN_2899; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2901 = 7'h54 == total_offset_51[6:0] ? phv_data_84 : _GEN_2900; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2902 = 7'h55 == total_offset_51[6:0] ? phv_data_85 : _GEN_2901; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2903 = 7'h56 == total_offset_51[6:0] ? phv_data_86 : _GEN_2902; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2904 = 7'h57 == total_offset_51[6:0] ? phv_data_87 : _GEN_2903; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2905 = 7'h58 == total_offset_51[6:0] ? phv_data_88 : _GEN_2904; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2906 = 7'h59 == total_offset_51[6:0] ? phv_data_89 : _GEN_2905; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2907 = 7'h5a == total_offset_51[6:0] ? phv_data_90 : _GEN_2906; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2908 = 7'h5b == total_offset_51[6:0] ? phv_data_91 : _GEN_2907; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2909 = 7'h5c == total_offset_51[6:0] ? phv_data_92 : _GEN_2908; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2910 = 7'h5d == total_offset_51[6:0] ? phv_data_93 : _GEN_2909; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2911 = 7'h5e == total_offset_51[6:0] ? phv_data_94 : _GEN_2910; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2912 = 7'h5f == total_offset_51[6:0] ? phv_data_95 : _GEN_2911; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_3 = 8'h3 < length_3 ? _GEN_2912 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_52 = offset_3 + 8'h4; // @[executor.scala 148:53]
  wire [7:0] _GEN_2915 = 7'h1 == total_offset_52[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2916 = 7'h2 == total_offset_52[6:0] ? phv_data_2 : _GEN_2915; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2917 = 7'h3 == total_offset_52[6:0] ? phv_data_3 : _GEN_2916; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2918 = 7'h4 == total_offset_52[6:0] ? phv_data_4 : _GEN_2917; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2919 = 7'h5 == total_offset_52[6:0] ? phv_data_5 : _GEN_2918; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2920 = 7'h6 == total_offset_52[6:0] ? phv_data_6 : _GEN_2919; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2921 = 7'h7 == total_offset_52[6:0] ? phv_data_7 : _GEN_2920; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2922 = 7'h8 == total_offset_52[6:0] ? phv_data_8 : _GEN_2921; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2923 = 7'h9 == total_offset_52[6:0] ? phv_data_9 : _GEN_2922; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2924 = 7'ha == total_offset_52[6:0] ? phv_data_10 : _GEN_2923; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2925 = 7'hb == total_offset_52[6:0] ? phv_data_11 : _GEN_2924; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2926 = 7'hc == total_offset_52[6:0] ? phv_data_12 : _GEN_2925; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2927 = 7'hd == total_offset_52[6:0] ? phv_data_13 : _GEN_2926; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2928 = 7'he == total_offset_52[6:0] ? phv_data_14 : _GEN_2927; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2929 = 7'hf == total_offset_52[6:0] ? phv_data_15 : _GEN_2928; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2930 = 7'h10 == total_offset_52[6:0] ? phv_data_16 : _GEN_2929; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2931 = 7'h11 == total_offset_52[6:0] ? phv_data_17 : _GEN_2930; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2932 = 7'h12 == total_offset_52[6:0] ? phv_data_18 : _GEN_2931; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2933 = 7'h13 == total_offset_52[6:0] ? phv_data_19 : _GEN_2932; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2934 = 7'h14 == total_offset_52[6:0] ? phv_data_20 : _GEN_2933; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2935 = 7'h15 == total_offset_52[6:0] ? phv_data_21 : _GEN_2934; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2936 = 7'h16 == total_offset_52[6:0] ? phv_data_22 : _GEN_2935; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2937 = 7'h17 == total_offset_52[6:0] ? phv_data_23 : _GEN_2936; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2938 = 7'h18 == total_offset_52[6:0] ? phv_data_24 : _GEN_2937; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2939 = 7'h19 == total_offset_52[6:0] ? phv_data_25 : _GEN_2938; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2940 = 7'h1a == total_offset_52[6:0] ? phv_data_26 : _GEN_2939; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2941 = 7'h1b == total_offset_52[6:0] ? phv_data_27 : _GEN_2940; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2942 = 7'h1c == total_offset_52[6:0] ? phv_data_28 : _GEN_2941; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2943 = 7'h1d == total_offset_52[6:0] ? phv_data_29 : _GEN_2942; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2944 = 7'h1e == total_offset_52[6:0] ? phv_data_30 : _GEN_2943; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2945 = 7'h1f == total_offset_52[6:0] ? phv_data_31 : _GEN_2944; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2946 = 7'h20 == total_offset_52[6:0] ? phv_data_32 : _GEN_2945; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2947 = 7'h21 == total_offset_52[6:0] ? phv_data_33 : _GEN_2946; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2948 = 7'h22 == total_offset_52[6:0] ? phv_data_34 : _GEN_2947; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2949 = 7'h23 == total_offset_52[6:0] ? phv_data_35 : _GEN_2948; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2950 = 7'h24 == total_offset_52[6:0] ? phv_data_36 : _GEN_2949; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2951 = 7'h25 == total_offset_52[6:0] ? phv_data_37 : _GEN_2950; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2952 = 7'h26 == total_offset_52[6:0] ? phv_data_38 : _GEN_2951; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2953 = 7'h27 == total_offset_52[6:0] ? phv_data_39 : _GEN_2952; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2954 = 7'h28 == total_offset_52[6:0] ? phv_data_40 : _GEN_2953; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2955 = 7'h29 == total_offset_52[6:0] ? phv_data_41 : _GEN_2954; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2956 = 7'h2a == total_offset_52[6:0] ? phv_data_42 : _GEN_2955; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2957 = 7'h2b == total_offset_52[6:0] ? phv_data_43 : _GEN_2956; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2958 = 7'h2c == total_offset_52[6:0] ? phv_data_44 : _GEN_2957; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2959 = 7'h2d == total_offset_52[6:0] ? phv_data_45 : _GEN_2958; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2960 = 7'h2e == total_offset_52[6:0] ? phv_data_46 : _GEN_2959; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2961 = 7'h2f == total_offset_52[6:0] ? phv_data_47 : _GEN_2960; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2962 = 7'h30 == total_offset_52[6:0] ? phv_data_48 : _GEN_2961; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2963 = 7'h31 == total_offset_52[6:0] ? phv_data_49 : _GEN_2962; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2964 = 7'h32 == total_offset_52[6:0] ? phv_data_50 : _GEN_2963; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2965 = 7'h33 == total_offset_52[6:0] ? phv_data_51 : _GEN_2964; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2966 = 7'h34 == total_offset_52[6:0] ? phv_data_52 : _GEN_2965; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2967 = 7'h35 == total_offset_52[6:0] ? phv_data_53 : _GEN_2966; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2968 = 7'h36 == total_offset_52[6:0] ? phv_data_54 : _GEN_2967; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2969 = 7'h37 == total_offset_52[6:0] ? phv_data_55 : _GEN_2968; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2970 = 7'h38 == total_offset_52[6:0] ? phv_data_56 : _GEN_2969; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2971 = 7'h39 == total_offset_52[6:0] ? phv_data_57 : _GEN_2970; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2972 = 7'h3a == total_offset_52[6:0] ? phv_data_58 : _GEN_2971; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2973 = 7'h3b == total_offset_52[6:0] ? phv_data_59 : _GEN_2972; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2974 = 7'h3c == total_offset_52[6:0] ? phv_data_60 : _GEN_2973; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2975 = 7'h3d == total_offset_52[6:0] ? phv_data_61 : _GEN_2974; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2976 = 7'h3e == total_offset_52[6:0] ? phv_data_62 : _GEN_2975; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2977 = 7'h3f == total_offset_52[6:0] ? phv_data_63 : _GEN_2976; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2978 = 7'h40 == total_offset_52[6:0] ? phv_data_64 : _GEN_2977; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2979 = 7'h41 == total_offset_52[6:0] ? phv_data_65 : _GEN_2978; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2980 = 7'h42 == total_offset_52[6:0] ? phv_data_66 : _GEN_2979; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2981 = 7'h43 == total_offset_52[6:0] ? phv_data_67 : _GEN_2980; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2982 = 7'h44 == total_offset_52[6:0] ? phv_data_68 : _GEN_2981; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2983 = 7'h45 == total_offset_52[6:0] ? phv_data_69 : _GEN_2982; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2984 = 7'h46 == total_offset_52[6:0] ? phv_data_70 : _GEN_2983; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2985 = 7'h47 == total_offset_52[6:0] ? phv_data_71 : _GEN_2984; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2986 = 7'h48 == total_offset_52[6:0] ? phv_data_72 : _GEN_2985; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2987 = 7'h49 == total_offset_52[6:0] ? phv_data_73 : _GEN_2986; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2988 = 7'h4a == total_offset_52[6:0] ? phv_data_74 : _GEN_2987; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2989 = 7'h4b == total_offset_52[6:0] ? phv_data_75 : _GEN_2988; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2990 = 7'h4c == total_offset_52[6:0] ? phv_data_76 : _GEN_2989; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2991 = 7'h4d == total_offset_52[6:0] ? phv_data_77 : _GEN_2990; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2992 = 7'h4e == total_offset_52[6:0] ? phv_data_78 : _GEN_2991; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2993 = 7'h4f == total_offset_52[6:0] ? phv_data_79 : _GEN_2992; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2994 = 7'h50 == total_offset_52[6:0] ? phv_data_80 : _GEN_2993; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2995 = 7'h51 == total_offset_52[6:0] ? phv_data_81 : _GEN_2994; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2996 = 7'h52 == total_offset_52[6:0] ? phv_data_82 : _GEN_2995; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2997 = 7'h53 == total_offset_52[6:0] ? phv_data_83 : _GEN_2996; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2998 = 7'h54 == total_offset_52[6:0] ? phv_data_84 : _GEN_2997; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_2999 = 7'h55 == total_offset_52[6:0] ? phv_data_85 : _GEN_2998; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3000 = 7'h56 == total_offset_52[6:0] ? phv_data_86 : _GEN_2999; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3001 = 7'h57 == total_offset_52[6:0] ? phv_data_87 : _GEN_3000; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3002 = 7'h58 == total_offset_52[6:0] ? phv_data_88 : _GEN_3001; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3003 = 7'h59 == total_offset_52[6:0] ? phv_data_89 : _GEN_3002; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3004 = 7'h5a == total_offset_52[6:0] ? phv_data_90 : _GEN_3003; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3005 = 7'h5b == total_offset_52[6:0] ? phv_data_91 : _GEN_3004; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3006 = 7'h5c == total_offset_52[6:0] ? phv_data_92 : _GEN_3005; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3007 = 7'h5d == total_offset_52[6:0] ? phv_data_93 : _GEN_3006; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3008 = 7'h5e == total_offset_52[6:0] ? phv_data_94 : _GEN_3007; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3009 = 7'h5f == total_offset_52[6:0] ? phv_data_95 : _GEN_3008; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_4 = 8'h4 < length_3 ? _GEN_3009 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_53 = offset_3 + 8'h5; // @[executor.scala 148:53]
  wire [7:0] _GEN_3012 = 7'h1 == total_offset_53[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3013 = 7'h2 == total_offset_53[6:0] ? phv_data_2 : _GEN_3012; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3014 = 7'h3 == total_offset_53[6:0] ? phv_data_3 : _GEN_3013; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3015 = 7'h4 == total_offset_53[6:0] ? phv_data_4 : _GEN_3014; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3016 = 7'h5 == total_offset_53[6:0] ? phv_data_5 : _GEN_3015; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3017 = 7'h6 == total_offset_53[6:0] ? phv_data_6 : _GEN_3016; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3018 = 7'h7 == total_offset_53[6:0] ? phv_data_7 : _GEN_3017; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3019 = 7'h8 == total_offset_53[6:0] ? phv_data_8 : _GEN_3018; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3020 = 7'h9 == total_offset_53[6:0] ? phv_data_9 : _GEN_3019; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3021 = 7'ha == total_offset_53[6:0] ? phv_data_10 : _GEN_3020; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3022 = 7'hb == total_offset_53[6:0] ? phv_data_11 : _GEN_3021; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3023 = 7'hc == total_offset_53[6:0] ? phv_data_12 : _GEN_3022; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3024 = 7'hd == total_offset_53[6:0] ? phv_data_13 : _GEN_3023; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3025 = 7'he == total_offset_53[6:0] ? phv_data_14 : _GEN_3024; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3026 = 7'hf == total_offset_53[6:0] ? phv_data_15 : _GEN_3025; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3027 = 7'h10 == total_offset_53[6:0] ? phv_data_16 : _GEN_3026; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3028 = 7'h11 == total_offset_53[6:0] ? phv_data_17 : _GEN_3027; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3029 = 7'h12 == total_offset_53[6:0] ? phv_data_18 : _GEN_3028; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3030 = 7'h13 == total_offset_53[6:0] ? phv_data_19 : _GEN_3029; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3031 = 7'h14 == total_offset_53[6:0] ? phv_data_20 : _GEN_3030; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3032 = 7'h15 == total_offset_53[6:0] ? phv_data_21 : _GEN_3031; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3033 = 7'h16 == total_offset_53[6:0] ? phv_data_22 : _GEN_3032; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3034 = 7'h17 == total_offset_53[6:0] ? phv_data_23 : _GEN_3033; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3035 = 7'h18 == total_offset_53[6:0] ? phv_data_24 : _GEN_3034; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3036 = 7'h19 == total_offset_53[6:0] ? phv_data_25 : _GEN_3035; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3037 = 7'h1a == total_offset_53[6:0] ? phv_data_26 : _GEN_3036; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3038 = 7'h1b == total_offset_53[6:0] ? phv_data_27 : _GEN_3037; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3039 = 7'h1c == total_offset_53[6:0] ? phv_data_28 : _GEN_3038; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3040 = 7'h1d == total_offset_53[6:0] ? phv_data_29 : _GEN_3039; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3041 = 7'h1e == total_offset_53[6:0] ? phv_data_30 : _GEN_3040; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3042 = 7'h1f == total_offset_53[6:0] ? phv_data_31 : _GEN_3041; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3043 = 7'h20 == total_offset_53[6:0] ? phv_data_32 : _GEN_3042; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3044 = 7'h21 == total_offset_53[6:0] ? phv_data_33 : _GEN_3043; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3045 = 7'h22 == total_offset_53[6:0] ? phv_data_34 : _GEN_3044; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3046 = 7'h23 == total_offset_53[6:0] ? phv_data_35 : _GEN_3045; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3047 = 7'h24 == total_offset_53[6:0] ? phv_data_36 : _GEN_3046; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3048 = 7'h25 == total_offset_53[6:0] ? phv_data_37 : _GEN_3047; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3049 = 7'h26 == total_offset_53[6:0] ? phv_data_38 : _GEN_3048; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3050 = 7'h27 == total_offset_53[6:0] ? phv_data_39 : _GEN_3049; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3051 = 7'h28 == total_offset_53[6:0] ? phv_data_40 : _GEN_3050; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3052 = 7'h29 == total_offset_53[6:0] ? phv_data_41 : _GEN_3051; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3053 = 7'h2a == total_offset_53[6:0] ? phv_data_42 : _GEN_3052; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3054 = 7'h2b == total_offset_53[6:0] ? phv_data_43 : _GEN_3053; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3055 = 7'h2c == total_offset_53[6:0] ? phv_data_44 : _GEN_3054; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3056 = 7'h2d == total_offset_53[6:0] ? phv_data_45 : _GEN_3055; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3057 = 7'h2e == total_offset_53[6:0] ? phv_data_46 : _GEN_3056; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3058 = 7'h2f == total_offset_53[6:0] ? phv_data_47 : _GEN_3057; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3059 = 7'h30 == total_offset_53[6:0] ? phv_data_48 : _GEN_3058; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3060 = 7'h31 == total_offset_53[6:0] ? phv_data_49 : _GEN_3059; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3061 = 7'h32 == total_offset_53[6:0] ? phv_data_50 : _GEN_3060; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3062 = 7'h33 == total_offset_53[6:0] ? phv_data_51 : _GEN_3061; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3063 = 7'h34 == total_offset_53[6:0] ? phv_data_52 : _GEN_3062; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3064 = 7'h35 == total_offset_53[6:0] ? phv_data_53 : _GEN_3063; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3065 = 7'h36 == total_offset_53[6:0] ? phv_data_54 : _GEN_3064; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3066 = 7'h37 == total_offset_53[6:0] ? phv_data_55 : _GEN_3065; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3067 = 7'h38 == total_offset_53[6:0] ? phv_data_56 : _GEN_3066; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3068 = 7'h39 == total_offset_53[6:0] ? phv_data_57 : _GEN_3067; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3069 = 7'h3a == total_offset_53[6:0] ? phv_data_58 : _GEN_3068; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3070 = 7'h3b == total_offset_53[6:0] ? phv_data_59 : _GEN_3069; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3071 = 7'h3c == total_offset_53[6:0] ? phv_data_60 : _GEN_3070; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3072 = 7'h3d == total_offset_53[6:0] ? phv_data_61 : _GEN_3071; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3073 = 7'h3e == total_offset_53[6:0] ? phv_data_62 : _GEN_3072; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3074 = 7'h3f == total_offset_53[6:0] ? phv_data_63 : _GEN_3073; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3075 = 7'h40 == total_offset_53[6:0] ? phv_data_64 : _GEN_3074; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3076 = 7'h41 == total_offset_53[6:0] ? phv_data_65 : _GEN_3075; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3077 = 7'h42 == total_offset_53[6:0] ? phv_data_66 : _GEN_3076; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3078 = 7'h43 == total_offset_53[6:0] ? phv_data_67 : _GEN_3077; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3079 = 7'h44 == total_offset_53[6:0] ? phv_data_68 : _GEN_3078; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3080 = 7'h45 == total_offset_53[6:0] ? phv_data_69 : _GEN_3079; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3081 = 7'h46 == total_offset_53[6:0] ? phv_data_70 : _GEN_3080; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3082 = 7'h47 == total_offset_53[6:0] ? phv_data_71 : _GEN_3081; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3083 = 7'h48 == total_offset_53[6:0] ? phv_data_72 : _GEN_3082; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3084 = 7'h49 == total_offset_53[6:0] ? phv_data_73 : _GEN_3083; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3085 = 7'h4a == total_offset_53[6:0] ? phv_data_74 : _GEN_3084; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3086 = 7'h4b == total_offset_53[6:0] ? phv_data_75 : _GEN_3085; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3087 = 7'h4c == total_offset_53[6:0] ? phv_data_76 : _GEN_3086; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3088 = 7'h4d == total_offset_53[6:0] ? phv_data_77 : _GEN_3087; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3089 = 7'h4e == total_offset_53[6:0] ? phv_data_78 : _GEN_3088; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3090 = 7'h4f == total_offset_53[6:0] ? phv_data_79 : _GEN_3089; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3091 = 7'h50 == total_offset_53[6:0] ? phv_data_80 : _GEN_3090; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3092 = 7'h51 == total_offset_53[6:0] ? phv_data_81 : _GEN_3091; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3093 = 7'h52 == total_offset_53[6:0] ? phv_data_82 : _GEN_3092; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3094 = 7'h53 == total_offset_53[6:0] ? phv_data_83 : _GEN_3093; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3095 = 7'h54 == total_offset_53[6:0] ? phv_data_84 : _GEN_3094; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3096 = 7'h55 == total_offset_53[6:0] ? phv_data_85 : _GEN_3095; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3097 = 7'h56 == total_offset_53[6:0] ? phv_data_86 : _GEN_3096; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3098 = 7'h57 == total_offset_53[6:0] ? phv_data_87 : _GEN_3097; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3099 = 7'h58 == total_offset_53[6:0] ? phv_data_88 : _GEN_3098; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3100 = 7'h59 == total_offset_53[6:0] ? phv_data_89 : _GEN_3099; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3101 = 7'h5a == total_offset_53[6:0] ? phv_data_90 : _GEN_3100; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3102 = 7'h5b == total_offset_53[6:0] ? phv_data_91 : _GEN_3101; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3103 = 7'h5c == total_offset_53[6:0] ? phv_data_92 : _GEN_3102; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3104 = 7'h5d == total_offset_53[6:0] ? phv_data_93 : _GEN_3103; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3105 = 7'h5e == total_offset_53[6:0] ? phv_data_94 : _GEN_3104; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3106 = 7'h5f == total_offset_53[6:0] ? phv_data_95 : _GEN_3105; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_5 = 8'h5 < length_3 ? _GEN_3106 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_54 = offset_3 + 8'h6; // @[executor.scala 148:53]
  wire [7:0] _GEN_3109 = 7'h1 == total_offset_54[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3110 = 7'h2 == total_offset_54[6:0] ? phv_data_2 : _GEN_3109; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3111 = 7'h3 == total_offset_54[6:0] ? phv_data_3 : _GEN_3110; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3112 = 7'h4 == total_offset_54[6:0] ? phv_data_4 : _GEN_3111; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3113 = 7'h5 == total_offset_54[6:0] ? phv_data_5 : _GEN_3112; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3114 = 7'h6 == total_offset_54[6:0] ? phv_data_6 : _GEN_3113; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3115 = 7'h7 == total_offset_54[6:0] ? phv_data_7 : _GEN_3114; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3116 = 7'h8 == total_offset_54[6:0] ? phv_data_8 : _GEN_3115; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3117 = 7'h9 == total_offset_54[6:0] ? phv_data_9 : _GEN_3116; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3118 = 7'ha == total_offset_54[6:0] ? phv_data_10 : _GEN_3117; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3119 = 7'hb == total_offset_54[6:0] ? phv_data_11 : _GEN_3118; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3120 = 7'hc == total_offset_54[6:0] ? phv_data_12 : _GEN_3119; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3121 = 7'hd == total_offset_54[6:0] ? phv_data_13 : _GEN_3120; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3122 = 7'he == total_offset_54[6:0] ? phv_data_14 : _GEN_3121; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3123 = 7'hf == total_offset_54[6:0] ? phv_data_15 : _GEN_3122; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3124 = 7'h10 == total_offset_54[6:0] ? phv_data_16 : _GEN_3123; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3125 = 7'h11 == total_offset_54[6:0] ? phv_data_17 : _GEN_3124; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3126 = 7'h12 == total_offset_54[6:0] ? phv_data_18 : _GEN_3125; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3127 = 7'h13 == total_offset_54[6:0] ? phv_data_19 : _GEN_3126; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3128 = 7'h14 == total_offset_54[6:0] ? phv_data_20 : _GEN_3127; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3129 = 7'h15 == total_offset_54[6:0] ? phv_data_21 : _GEN_3128; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3130 = 7'h16 == total_offset_54[6:0] ? phv_data_22 : _GEN_3129; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3131 = 7'h17 == total_offset_54[6:0] ? phv_data_23 : _GEN_3130; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3132 = 7'h18 == total_offset_54[6:0] ? phv_data_24 : _GEN_3131; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3133 = 7'h19 == total_offset_54[6:0] ? phv_data_25 : _GEN_3132; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3134 = 7'h1a == total_offset_54[6:0] ? phv_data_26 : _GEN_3133; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3135 = 7'h1b == total_offset_54[6:0] ? phv_data_27 : _GEN_3134; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3136 = 7'h1c == total_offset_54[6:0] ? phv_data_28 : _GEN_3135; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3137 = 7'h1d == total_offset_54[6:0] ? phv_data_29 : _GEN_3136; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3138 = 7'h1e == total_offset_54[6:0] ? phv_data_30 : _GEN_3137; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3139 = 7'h1f == total_offset_54[6:0] ? phv_data_31 : _GEN_3138; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3140 = 7'h20 == total_offset_54[6:0] ? phv_data_32 : _GEN_3139; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3141 = 7'h21 == total_offset_54[6:0] ? phv_data_33 : _GEN_3140; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3142 = 7'h22 == total_offset_54[6:0] ? phv_data_34 : _GEN_3141; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3143 = 7'h23 == total_offset_54[6:0] ? phv_data_35 : _GEN_3142; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3144 = 7'h24 == total_offset_54[6:0] ? phv_data_36 : _GEN_3143; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3145 = 7'h25 == total_offset_54[6:0] ? phv_data_37 : _GEN_3144; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3146 = 7'h26 == total_offset_54[6:0] ? phv_data_38 : _GEN_3145; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3147 = 7'h27 == total_offset_54[6:0] ? phv_data_39 : _GEN_3146; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3148 = 7'h28 == total_offset_54[6:0] ? phv_data_40 : _GEN_3147; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3149 = 7'h29 == total_offset_54[6:0] ? phv_data_41 : _GEN_3148; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3150 = 7'h2a == total_offset_54[6:0] ? phv_data_42 : _GEN_3149; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3151 = 7'h2b == total_offset_54[6:0] ? phv_data_43 : _GEN_3150; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3152 = 7'h2c == total_offset_54[6:0] ? phv_data_44 : _GEN_3151; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3153 = 7'h2d == total_offset_54[6:0] ? phv_data_45 : _GEN_3152; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3154 = 7'h2e == total_offset_54[6:0] ? phv_data_46 : _GEN_3153; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3155 = 7'h2f == total_offset_54[6:0] ? phv_data_47 : _GEN_3154; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3156 = 7'h30 == total_offset_54[6:0] ? phv_data_48 : _GEN_3155; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3157 = 7'h31 == total_offset_54[6:0] ? phv_data_49 : _GEN_3156; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3158 = 7'h32 == total_offset_54[6:0] ? phv_data_50 : _GEN_3157; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3159 = 7'h33 == total_offset_54[6:0] ? phv_data_51 : _GEN_3158; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3160 = 7'h34 == total_offset_54[6:0] ? phv_data_52 : _GEN_3159; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3161 = 7'h35 == total_offset_54[6:0] ? phv_data_53 : _GEN_3160; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3162 = 7'h36 == total_offset_54[6:0] ? phv_data_54 : _GEN_3161; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3163 = 7'h37 == total_offset_54[6:0] ? phv_data_55 : _GEN_3162; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3164 = 7'h38 == total_offset_54[6:0] ? phv_data_56 : _GEN_3163; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3165 = 7'h39 == total_offset_54[6:0] ? phv_data_57 : _GEN_3164; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3166 = 7'h3a == total_offset_54[6:0] ? phv_data_58 : _GEN_3165; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3167 = 7'h3b == total_offset_54[6:0] ? phv_data_59 : _GEN_3166; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3168 = 7'h3c == total_offset_54[6:0] ? phv_data_60 : _GEN_3167; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3169 = 7'h3d == total_offset_54[6:0] ? phv_data_61 : _GEN_3168; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3170 = 7'h3e == total_offset_54[6:0] ? phv_data_62 : _GEN_3169; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3171 = 7'h3f == total_offset_54[6:0] ? phv_data_63 : _GEN_3170; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3172 = 7'h40 == total_offset_54[6:0] ? phv_data_64 : _GEN_3171; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3173 = 7'h41 == total_offset_54[6:0] ? phv_data_65 : _GEN_3172; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3174 = 7'h42 == total_offset_54[6:0] ? phv_data_66 : _GEN_3173; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3175 = 7'h43 == total_offset_54[6:0] ? phv_data_67 : _GEN_3174; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3176 = 7'h44 == total_offset_54[6:0] ? phv_data_68 : _GEN_3175; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3177 = 7'h45 == total_offset_54[6:0] ? phv_data_69 : _GEN_3176; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3178 = 7'h46 == total_offset_54[6:0] ? phv_data_70 : _GEN_3177; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3179 = 7'h47 == total_offset_54[6:0] ? phv_data_71 : _GEN_3178; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3180 = 7'h48 == total_offset_54[6:0] ? phv_data_72 : _GEN_3179; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3181 = 7'h49 == total_offset_54[6:0] ? phv_data_73 : _GEN_3180; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3182 = 7'h4a == total_offset_54[6:0] ? phv_data_74 : _GEN_3181; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3183 = 7'h4b == total_offset_54[6:0] ? phv_data_75 : _GEN_3182; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3184 = 7'h4c == total_offset_54[6:0] ? phv_data_76 : _GEN_3183; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3185 = 7'h4d == total_offset_54[6:0] ? phv_data_77 : _GEN_3184; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3186 = 7'h4e == total_offset_54[6:0] ? phv_data_78 : _GEN_3185; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3187 = 7'h4f == total_offset_54[6:0] ? phv_data_79 : _GEN_3186; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3188 = 7'h50 == total_offset_54[6:0] ? phv_data_80 : _GEN_3187; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3189 = 7'h51 == total_offset_54[6:0] ? phv_data_81 : _GEN_3188; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3190 = 7'h52 == total_offset_54[6:0] ? phv_data_82 : _GEN_3189; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3191 = 7'h53 == total_offset_54[6:0] ? phv_data_83 : _GEN_3190; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3192 = 7'h54 == total_offset_54[6:0] ? phv_data_84 : _GEN_3191; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3193 = 7'h55 == total_offset_54[6:0] ? phv_data_85 : _GEN_3192; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3194 = 7'h56 == total_offset_54[6:0] ? phv_data_86 : _GEN_3193; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3195 = 7'h57 == total_offset_54[6:0] ? phv_data_87 : _GEN_3194; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3196 = 7'h58 == total_offset_54[6:0] ? phv_data_88 : _GEN_3195; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3197 = 7'h59 == total_offset_54[6:0] ? phv_data_89 : _GEN_3196; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3198 = 7'h5a == total_offset_54[6:0] ? phv_data_90 : _GEN_3197; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3199 = 7'h5b == total_offset_54[6:0] ? phv_data_91 : _GEN_3198; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3200 = 7'h5c == total_offset_54[6:0] ? phv_data_92 : _GEN_3199; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3201 = 7'h5d == total_offset_54[6:0] ? phv_data_93 : _GEN_3200; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3202 = 7'h5e == total_offset_54[6:0] ? phv_data_94 : _GEN_3201; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3203 = 7'h5f == total_offset_54[6:0] ? phv_data_95 : _GEN_3202; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_6 = 8'h6 < length_3 ? _GEN_3203 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [7:0] total_offset_55 = offset_3 + 8'h7; // @[executor.scala 148:53]
  wire [7:0] _GEN_3206 = 7'h1 == total_offset_55[6:0] ? phv_data_1 : phv_data_0; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3207 = 7'h2 == total_offset_55[6:0] ? phv_data_2 : _GEN_3206; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3208 = 7'h3 == total_offset_55[6:0] ? phv_data_3 : _GEN_3207; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3209 = 7'h4 == total_offset_55[6:0] ? phv_data_4 : _GEN_3208; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3210 = 7'h5 == total_offset_55[6:0] ? phv_data_5 : _GEN_3209; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3211 = 7'h6 == total_offset_55[6:0] ? phv_data_6 : _GEN_3210; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3212 = 7'h7 == total_offset_55[6:0] ? phv_data_7 : _GEN_3211; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3213 = 7'h8 == total_offset_55[6:0] ? phv_data_8 : _GEN_3212; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3214 = 7'h9 == total_offset_55[6:0] ? phv_data_9 : _GEN_3213; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3215 = 7'ha == total_offset_55[6:0] ? phv_data_10 : _GEN_3214; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3216 = 7'hb == total_offset_55[6:0] ? phv_data_11 : _GEN_3215; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3217 = 7'hc == total_offset_55[6:0] ? phv_data_12 : _GEN_3216; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3218 = 7'hd == total_offset_55[6:0] ? phv_data_13 : _GEN_3217; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3219 = 7'he == total_offset_55[6:0] ? phv_data_14 : _GEN_3218; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3220 = 7'hf == total_offset_55[6:0] ? phv_data_15 : _GEN_3219; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3221 = 7'h10 == total_offset_55[6:0] ? phv_data_16 : _GEN_3220; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3222 = 7'h11 == total_offset_55[6:0] ? phv_data_17 : _GEN_3221; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3223 = 7'h12 == total_offset_55[6:0] ? phv_data_18 : _GEN_3222; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3224 = 7'h13 == total_offset_55[6:0] ? phv_data_19 : _GEN_3223; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3225 = 7'h14 == total_offset_55[6:0] ? phv_data_20 : _GEN_3224; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3226 = 7'h15 == total_offset_55[6:0] ? phv_data_21 : _GEN_3225; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3227 = 7'h16 == total_offset_55[6:0] ? phv_data_22 : _GEN_3226; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3228 = 7'h17 == total_offset_55[6:0] ? phv_data_23 : _GEN_3227; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3229 = 7'h18 == total_offset_55[6:0] ? phv_data_24 : _GEN_3228; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3230 = 7'h19 == total_offset_55[6:0] ? phv_data_25 : _GEN_3229; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3231 = 7'h1a == total_offset_55[6:0] ? phv_data_26 : _GEN_3230; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3232 = 7'h1b == total_offset_55[6:0] ? phv_data_27 : _GEN_3231; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3233 = 7'h1c == total_offset_55[6:0] ? phv_data_28 : _GEN_3232; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3234 = 7'h1d == total_offset_55[6:0] ? phv_data_29 : _GEN_3233; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3235 = 7'h1e == total_offset_55[6:0] ? phv_data_30 : _GEN_3234; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3236 = 7'h1f == total_offset_55[6:0] ? phv_data_31 : _GEN_3235; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3237 = 7'h20 == total_offset_55[6:0] ? phv_data_32 : _GEN_3236; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3238 = 7'h21 == total_offset_55[6:0] ? phv_data_33 : _GEN_3237; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3239 = 7'h22 == total_offset_55[6:0] ? phv_data_34 : _GEN_3238; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3240 = 7'h23 == total_offset_55[6:0] ? phv_data_35 : _GEN_3239; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3241 = 7'h24 == total_offset_55[6:0] ? phv_data_36 : _GEN_3240; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3242 = 7'h25 == total_offset_55[6:0] ? phv_data_37 : _GEN_3241; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3243 = 7'h26 == total_offset_55[6:0] ? phv_data_38 : _GEN_3242; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3244 = 7'h27 == total_offset_55[6:0] ? phv_data_39 : _GEN_3243; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3245 = 7'h28 == total_offset_55[6:0] ? phv_data_40 : _GEN_3244; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3246 = 7'h29 == total_offset_55[6:0] ? phv_data_41 : _GEN_3245; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3247 = 7'h2a == total_offset_55[6:0] ? phv_data_42 : _GEN_3246; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3248 = 7'h2b == total_offset_55[6:0] ? phv_data_43 : _GEN_3247; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3249 = 7'h2c == total_offset_55[6:0] ? phv_data_44 : _GEN_3248; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3250 = 7'h2d == total_offset_55[6:0] ? phv_data_45 : _GEN_3249; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3251 = 7'h2e == total_offset_55[6:0] ? phv_data_46 : _GEN_3250; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3252 = 7'h2f == total_offset_55[6:0] ? phv_data_47 : _GEN_3251; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3253 = 7'h30 == total_offset_55[6:0] ? phv_data_48 : _GEN_3252; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3254 = 7'h31 == total_offset_55[6:0] ? phv_data_49 : _GEN_3253; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3255 = 7'h32 == total_offset_55[6:0] ? phv_data_50 : _GEN_3254; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3256 = 7'h33 == total_offset_55[6:0] ? phv_data_51 : _GEN_3255; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3257 = 7'h34 == total_offset_55[6:0] ? phv_data_52 : _GEN_3256; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3258 = 7'h35 == total_offset_55[6:0] ? phv_data_53 : _GEN_3257; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3259 = 7'h36 == total_offset_55[6:0] ? phv_data_54 : _GEN_3258; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3260 = 7'h37 == total_offset_55[6:0] ? phv_data_55 : _GEN_3259; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3261 = 7'h38 == total_offset_55[6:0] ? phv_data_56 : _GEN_3260; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3262 = 7'h39 == total_offset_55[6:0] ? phv_data_57 : _GEN_3261; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3263 = 7'h3a == total_offset_55[6:0] ? phv_data_58 : _GEN_3262; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3264 = 7'h3b == total_offset_55[6:0] ? phv_data_59 : _GEN_3263; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3265 = 7'h3c == total_offset_55[6:0] ? phv_data_60 : _GEN_3264; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3266 = 7'h3d == total_offset_55[6:0] ? phv_data_61 : _GEN_3265; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3267 = 7'h3e == total_offset_55[6:0] ? phv_data_62 : _GEN_3266; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3268 = 7'h3f == total_offset_55[6:0] ? phv_data_63 : _GEN_3267; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3269 = 7'h40 == total_offset_55[6:0] ? phv_data_64 : _GEN_3268; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3270 = 7'h41 == total_offset_55[6:0] ? phv_data_65 : _GEN_3269; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3271 = 7'h42 == total_offset_55[6:0] ? phv_data_66 : _GEN_3270; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3272 = 7'h43 == total_offset_55[6:0] ? phv_data_67 : _GEN_3271; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3273 = 7'h44 == total_offset_55[6:0] ? phv_data_68 : _GEN_3272; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3274 = 7'h45 == total_offset_55[6:0] ? phv_data_69 : _GEN_3273; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3275 = 7'h46 == total_offset_55[6:0] ? phv_data_70 : _GEN_3274; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3276 = 7'h47 == total_offset_55[6:0] ? phv_data_71 : _GEN_3275; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3277 = 7'h48 == total_offset_55[6:0] ? phv_data_72 : _GEN_3276; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3278 = 7'h49 == total_offset_55[6:0] ? phv_data_73 : _GEN_3277; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3279 = 7'h4a == total_offset_55[6:0] ? phv_data_74 : _GEN_3278; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3280 = 7'h4b == total_offset_55[6:0] ? phv_data_75 : _GEN_3279; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3281 = 7'h4c == total_offset_55[6:0] ? phv_data_76 : _GEN_3280; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3282 = 7'h4d == total_offset_55[6:0] ? phv_data_77 : _GEN_3281; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3283 = 7'h4e == total_offset_55[6:0] ? phv_data_78 : _GEN_3282; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3284 = 7'h4f == total_offset_55[6:0] ? phv_data_79 : _GEN_3283; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3285 = 7'h50 == total_offset_55[6:0] ? phv_data_80 : _GEN_3284; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3286 = 7'h51 == total_offset_55[6:0] ? phv_data_81 : _GEN_3285; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3287 = 7'h52 == total_offset_55[6:0] ? phv_data_82 : _GEN_3286; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3288 = 7'h53 == total_offset_55[6:0] ? phv_data_83 : _GEN_3287; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3289 = 7'h54 == total_offset_55[6:0] ? phv_data_84 : _GEN_3288; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3290 = 7'h55 == total_offset_55[6:0] ? phv_data_85 : _GEN_3289; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3291 = 7'h56 == total_offset_55[6:0] ? phv_data_86 : _GEN_3290; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3292 = 7'h57 == total_offset_55[6:0] ? phv_data_87 : _GEN_3291; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3293 = 7'h58 == total_offset_55[6:0] ? phv_data_88 : _GEN_3292; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3294 = 7'h59 == total_offset_55[6:0] ? phv_data_89 : _GEN_3293; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3295 = 7'h5a == total_offset_55[6:0] ? phv_data_90 : _GEN_3294; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3296 = 7'h5b == total_offset_55[6:0] ? phv_data_91 : _GEN_3295; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3297 = 7'h5c == total_offset_55[6:0] ? phv_data_92 : _GEN_3296; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3298 = 7'h5d == total_offset_55[6:0] ? phv_data_93 : _GEN_3297; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3299 = 7'h5e == total_offset_55[6:0] ? phv_data_94 : _GEN_3298; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] _GEN_3300 = 7'h5f == total_offset_55[6:0] ? phv_data_95 : _GEN_3299; // @[executor.scala 150:34 executor.scala 150:34]
  wire [7:0] bytes_6_7 = 8'h7 < length_3 ? _GEN_3300 : 8'h0; // @[executor.scala 149:56 executor.scala 150:34 executor.scala 152:34]
  wire [63:0] _io_field_out_3_T = {bytes_6_0,bytes_6_1,bytes_6_2,bytes_6_3,bytes_6_4,bytes_6_5,bytes_6_6,bytes_6_7}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_3 = io_field_out_3_lo[13:11]; // @[primitive.scala 34:52]
  wire [2:0] args_length_3 = io_field_out_3_lo[10:8]; // @[primitive.scala 35:52]
  wire [8:0] _total_offset_T_56 = {{6'd0}, args_offset_3}; // @[executor.scala 163:56]
  wire [7:0] total_offset_56 = _total_offset_T_56[7:0]; // @[executor.scala 163:56]
  wire [7:0] _GEN_3410 = {{5'd0}, args_length_3}; // @[executor.scala 164:44]
  wire [7:0] _GEN_3303 = 3'h1 == total_offset_56[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3304 = 3'h2 == total_offset_56[2:0] ? args_2 : _GEN_3303; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3305 = 3'h3 == total_offset_56[2:0] ? args_3 : _GEN_3304; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3306 = 3'h4 == total_offset_56[2:0] ? args_4 : _GEN_3305; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3307 = 3'h5 == total_offset_56[2:0] ? args_5 : _GEN_3306; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3308 = 3'h6 == total_offset_56[2:0] ? args_6 : _GEN_3307; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_7_0 = 8'h0 < _GEN_3410 ? _GEN_3308 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] _GEN_3411 = {{5'd0}, args_offset_3}; // @[executor.scala 163:56]
  wire [7:0] total_offset_57 = _GEN_3411 + 8'h1; // @[executor.scala 163:56]
  wire [7:0] _GEN_3311 = 3'h1 == total_offset_57[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3312 = 3'h2 == total_offset_57[2:0] ? args_2 : _GEN_3311; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3313 = 3'h3 == total_offset_57[2:0] ? args_3 : _GEN_3312; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3314 = 3'h4 == total_offset_57[2:0] ? args_4 : _GEN_3313; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3315 = 3'h5 == total_offset_57[2:0] ? args_5 : _GEN_3314; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3316 = 3'h6 == total_offset_57[2:0] ? args_6 : _GEN_3315; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_7_1 = 8'h1 < _GEN_3410 ? _GEN_3316 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_58 = _GEN_3411 + 8'h2; // @[executor.scala 163:56]
  wire [7:0] _GEN_3319 = 3'h1 == total_offset_58[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3320 = 3'h2 == total_offset_58[2:0] ? args_2 : _GEN_3319; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3321 = 3'h3 == total_offset_58[2:0] ? args_3 : _GEN_3320; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3322 = 3'h4 == total_offset_58[2:0] ? args_4 : _GEN_3321; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3323 = 3'h5 == total_offset_58[2:0] ? args_5 : _GEN_3322; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3324 = 3'h6 == total_offset_58[2:0] ? args_6 : _GEN_3323; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_7_2 = 8'h2 < _GEN_3410 ? _GEN_3324 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_59 = _GEN_3411 + 8'h3; // @[executor.scala 163:56]
  wire [7:0] _GEN_3327 = 3'h1 == total_offset_59[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3328 = 3'h2 == total_offset_59[2:0] ? args_2 : _GEN_3327; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3329 = 3'h3 == total_offset_59[2:0] ? args_3 : _GEN_3328; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3330 = 3'h4 == total_offset_59[2:0] ? args_4 : _GEN_3329; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3331 = 3'h5 == total_offset_59[2:0] ? args_5 : _GEN_3330; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3332 = 3'h6 == total_offset_59[2:0] ? args_6 : _GEN_3331; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_7_3 = 8'h3 < _GEN_3410 ? _GEN_3332 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_60 = _GEN_3411 + 8'h4; // @[executor.scala 163:56]
  wire [7:0] _GEN_3335 = 3'h1 == total_offset_60[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3336 = 3'h2 == total_offset_60[2:0] ? args_2 : _GEN_3335; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3337 = 3'h3 == total_offset_60[2:0] ? args_3 : _GEN_3336; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3338 = 3'h4 == total_offset_60[2:0] ? args_4 : _GEN_3337; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3339 = 3'h5 == total_offset_60[2:0] ? args_5 : _GEN_3338; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3340 = 3'h6 == total_offset_60[2:0] ? args_6 : _GEN_3339; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_7_4 = 8'h4 < _GEN_3410 ? _GEN_3340 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_61 = _GEN_3411 + 8'h5; // @[executor.scala 163:56]
  wire [7:0] _GEN_3343 = 3'h1 == total_offset_61[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3344 = 3'h2 == total_offset_61[2:0] ? args_2 : _GEN_3343; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3345 = 3'h3 == total_offset_61[2:0] ? args_3 : _GEN_3344; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3346 = 3'h4 == total_offset_61[2:0] ? args_4 : _GEN_3345; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3347 = 3'h5 == total_offset_61[2:0] ? args_5 : _GEN_3346; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3348 = 3'h6 == total_offset_61[2:0] ? args_6 : _GEN_3347; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_7_5 = 8'h5 < _GEN_3410 ? _GEN_3348 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [7:0] total_offset_62 = _GEN_3411 + 8'h6; // @[executor.scala 163:56]
  wire [7:0] _GEN_3351 = 3'h1 == total_offset_62[2:0] ? args_1 : args_0; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3352 = 3'h2 == total_offset_62[2:0] ? args_2 : _GEN_3351; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3353 = 3'h3 == total_offset_62[2:0] ? args_3 : _GEN_3352; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3354 = 3'h4 == total_offset_62[2:0] ? args_4 : _GEN_3353; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3355 = 3'h5 == total_offset_62[2:0] ? args_5 : _GEN_3354; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] _GEN_3356 = 3'h6 == total_offset_62[2:0] ? args_6 : _GEN_3355; // @[executor.scala 165:38 executor.scala 165:38]
  wire [7:0] bytes_7_6 = 8'h6 < _GEN_3410 ? _GEN_3356 : 8'h0; // @[executor.scala 164:59 executor.scala 165:38 executor.scala 167:38]
  wire [63:0] _io_field_out_3_T_1 = {bytes_7_0,bytes_7_1,bytes_7_2,bytes_7_3,bytes_7_4,bytes_7_5,bytes_7_6,8'h0}; // @[Cat.scala 30:58]
  wire [49:0] io_field_out_3_hi_12 = io_field_out_3_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_field_out_3_T_4 = {io_field_out_3_hi_12,io_field_out_3_lo}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_3366 = 4'ha == opcode_3 ? _io_field_out_3_T_1 : _io_field_out_3_T_4; // @[executor.scala 157:51 executor.scala 170:37 executor.scala 173:37]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 121:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 121:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 121:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 121:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 121:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 121:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 121:25]
  assign io_vliw_out_0 = vliw_0; // @[executor.scala 128:21]
  assign io_vliw_out_1 = vliw_1; // @[executor.scala 128:21]
  assign io_vliw_out_2 = vliw_2; // @[executor.scala 128:21]
  assign io_vliw_out_3 = vliw_3; // @[executor.scala 128:21]
  assign io_field_out_0 = from_header ? _io_field_out_0_T : _GEN_840; // @[executor.scala 142:32 executor.scala 155:33]
  assign io_field_out_1 = from_header_1 ? _io_field_out_1_T : _GEN_1682; // @[executor.scala 142:32 executor.scala 155:33]
  assign io_field_out_2 = from_header_2 ? _io_field_out_2_T : _GEN_2524; // @[executor.scala 142:32 executor.scala 155:33]
  assign io_field_out_3 = from_header_3 ? _io_field_out_3_T : _GEN_3366; // @[executor.scala 142:32 executor.scala 155:33]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 120:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 120:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 120:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 120:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 120:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 120:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 120:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 120:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 120:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 120:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 120:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 120:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 120:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 120:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 120:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 120:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 120:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 120:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 120:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 120:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 120:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 120:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 120:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 120:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 120:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 120:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 120:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 120:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 120:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 120:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 120:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 120:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 120:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 120:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 120:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 120:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 120:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 120:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 120:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 120:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 120:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 120:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 120:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 120:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 120:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 120:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 120:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 120:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 120:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 120:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 120:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 120:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 120:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 120:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 120:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 120:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 120:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 120:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 120:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 120:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 120:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 120:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 120:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 120:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 120:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 120:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 120:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 120:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 120:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 120:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 120:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 120:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 120:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 120:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 120:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 120:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 120:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 120:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 120:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 120:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 120:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 120:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 120:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 120:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 120:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 120:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 120:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 120:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 120:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 120:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 120:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 120:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 120:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 120:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 120:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 120:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 120:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 120:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 120:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 120:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 120:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 120:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 120:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 120:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 120:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 120:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 120:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 120:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 120:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 120:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 120:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 120:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 120:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 120:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 120:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 120:13]
    args_0 <= io_args_in_0; // @[executor.scala 124:14]
    args_1 <= io_args_in_1; // @[executor.scala 124:14]
    args_2 <= io_args_in_2; // @[executor.scala 124:14]
    args_3 <= io_args_in_3; // @[executor.scala 124:14]
    args_4 <= io_args_in_4; // @[executor.scala 124:14]
    args_5 <= io_args_in_5; // @[executor.scala 124:14]
    args_6 <= io_args_in_6; // @[executor.scala 124:14]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 127:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 127:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 127:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 127:14]
    offset_0 <= io_offset_in_0; // @[executor.scala 132:16]
    offset_1 <= io_offset_in_1; // @[executor.scala 132:16]
    offset_2 <= io_offset_in_2; // @[executor.scala 132:16]
    offset_3 <= io_offset_in_3; // @[executor.scala 132:16]
    length_0 <= io_length_in_0; // @[executor.scala 133:16]
    length_1 <= io_length_in_1; // @[executor.scala 133:16]
    length_2 <= io_length_in_2; // @[executor.scala 133:16]
    length_3 <= io_length_in_3; // @[executor.scala 133:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  args_0 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  args_1 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  args_2 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  args_3 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  args_4 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  args_5 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  args_6 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  vliw_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  vliw_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  vliw_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  vliw_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  offset_0 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  offset_1 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  offset_2 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  offset_3 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  length_0 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  length_1 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  length_2 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  length_3 = _RAND_134[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PrimitiveALU(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [63:0] io_field_in_0,
  input  [63:0] io_field_in_1,
  input  [63:0] io_field_in_2,
  input  [63:0] io_field_in_3,
  output [31:0] io_vliw_out_0,
  output [31:0] io_vliw_out_1,
  output [31:0] io_vliw_out_2,
  output [31:0] io_vliw_out_3,
  output [63:0] io_field_out_0,
  output [63:0] io_field_out_1,
  output [63:0] io_field_out_2,
  output [63:0] io_field_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 190:22]
  reg [7:0] phv_data_1; // @[executor.scala 190:22]
  reg [7:0] phv_data_2; // @[executor.scala 190:22]
  reg [7:0] phv_data_3; // @[executor.scala 190:22]
  reg [7:0] phv_data_4; // @[executor.scala 190:22]
  reg [7:0] phv_data_5; // @[executor.scala 190:22]
  reg [7:0] phv_data_6; // @[executor.scala 190:22]
  reg [7:0] phv_data_7; // @[executor.scala 190:22]
  reg [7:0] phv_data_8; // @[executor.scala 190:22]
  reg [7:0] phv_data_9; // @[executor.scala 190:22]
  reg [7:0] phv_data_10; // @[executor.scala 190:22]
  reg [7:0] phv_data_11; // @[executor.scala 190:22]
  reg [7:0] phv_data_12; // @[executor.scala 190:22]
  reg [7:0] phv_data_13; // @[executor.scala 190:22]
  reg [7:0] phv_data_14; // @[executor.scala 190:22]
  reg [7:0] phv_data_15; // @[executor.scala 190:22]
  reg [7:0] phv_data_16; // @[executor.scala 190:22]
  reg [7:0] phv_data_17; // @[executor.scala 190:22]
  reg [7:0] phv_data_18; // @[executor.scala 190:22]
  reg [7:0] phv_data_19; // @[executor.scala 190:22]
  reg [7:0] phv_data_20; // @[executor.scala 190:22]
  reg [7:0] phv_data_21; // @[executor.scala 190:22]
  reg [7:0] phv_data_22; // @[executor.scala 190:22]
  reg [7:0] phv_data_23; // @[executor.scala 190:22]
  reg [7:0] phv_data_24; // @[executor.scala 190:22]
  reg [7:0] phv_data_25; // @[executor.scala 190:22]
  reg [7:0] phv_data_26; // @[executor.scala 190:22]
  reg [7:0] phv_data_27; // @[executor.scala 190:22]
  reg [7:0] phv_data_28; // @[executor.scala 190:22]
  reg [7:0] phv_data_29; // @[executor.scala 190:22]
  reg [7:0] phv_data_30; // @[executor.scala 190:22]
  reg [7:0] phv_data_31; // @[executor.scala 190:22]
  reg [7:0] phv_data_32; // @[executor.scala 190:22]
  reg [7:0] phv_data_33; // @[executor.scala 190:22]
  reg [7:0] phv_data_34; // @[executor.scala 190:22]
  reg [7:0] phv_data_35; // @[executor.scala 190:22]
  reg [7:0] phv_data_36; // @[executor.scala 190:22]
  reg [7:0] phv_data_37; // @[executor.scala 190:22]
  reg [7:0] phv_data_38; // @[executor.scala 190:22]
  reg [7:0] phv_data_39; // @[executor.scala 190:22]
  reg [7:0] phv_data_40; // @[executor.scala 190:22]
  reg [7:0] phv_data_41; // @[executor.scala 190:22]
  reg [7:0] phv_data_42; // @[executor.scala 190:22]
  reg [7:0] phv_data_43; // @[executor.scala 190:22]
  reg [7:0] phv_data_44; // @[executor.scala 190:22]
  reg [7:0] phv_data_45; // @[executor.scala 190:22]
  reg [7:0] phv_data_46; // @[executor.scala 190:22]
  reg [7:0] phv_data_47; // @[executor.scala 190:22]
  reg [7:0] phv_data_48; // @[executor.scala 190:22]
  reg [7:0] phv_data_49; // @[executor.scala 190:22]
  reg [7:0] phv_data_50; // @[executor.scala 190:22]
  reg [7:0] phv_data_51; // @[executor.scala 190:22]
  reg [7:0] phv_data_52; // @[executor.scala 190:22]
  reg [7:0] phv_data_53; // @[executor.scala 190:22]
  reg [7:0] phv_data_54; // @[executor.scala 190:22]
  reg [7:0] phv_data_55; // @[executor.scala 190:22]
  reg [7:0] phv_data_56; // @[executor.scala 190:22]
  reg [7:0] phv_data_57; // @[executor.scala 190:22]
  reg [7:0] phv_data_58; // @[executor.scala 190:22]
  reg [7:0] phv_data_59; // @[executor.scala 190:22]
  reg [7:0] phv_data_60; // @[executor.scala 190:22]
  reg [7:0] phv_data_61; // @[executor.scala 190:22]
  reg [7:0] phv_data_62; // @[executor.scala 190:22]
  reg [7:0] phv_data_63; // @[executor.scala 190:22]
  reg [7:0] phv_data_64; // @[executor.scala 190:22]
  reg [7:0] phv_data_65; // @[executor.scala 190:22]
  reg [7:0] phv_data_66; // @[executor.scala 190:22]
  reg [7:0] phv_data_67; // @[executor.scala 190:22]
  reg [7:0] phv_data_68; // @[executor.scala 190:22]
  reg [7:0] phv_data_69; // @[executor.scala 190:22]
  reg [7:0] phv_data_70; // @[executor.scala 190:22]
  reg [7:0] phv_data_71; // @[executor.scala 190:22]
  reg [7:0] phv_data_72; // @[executor.scala 190:22]
  reg [7:0] phv_data_73; // @[executor.scala 190:22]
  reg [7:0] phv_data_74; // @[executor.scala 190:22]
  reg [7:0] phv_data_75; // @[executor.scala 190:22]
  reg [7:0] phv_data_76; // @[executor.scala 190:22]
  reg [7:0] phv_data_77; // @[executor.scala 190:22]
  reg [7:0] phv_data_78; // @[executor.scala 190:22]
  reg [7:0] phv_data_79; // @[executor.scala 190:22]
  reg [7:0] phv_data_80; // @[executor.scala 190:22]
  reg [7:0] phv_data_81; // @[executor.scala 190:22]
  reg [7:0] phv_data_82; // @[executor.scala 190:22]
  reg [7:0] phv_data_83; // @[executor.scala 190:22]
  reg [7:0] phv_data_84; // @[executor.scala 190:22]
  reg [7:0] phv_data_85; // @[executor.scala 190:22]
  reg [7:0] phv_data_86; // @[executor.scala 190:22]
  reg [7:0] phv_data_87; // @[executor.scala 190:22]
  reg [7:0] phv_data_88; // @[executor.scala 190:22]
  reg [7:0] phv_data_89; // @[executor.scala 190:22]
  reg [7:0] phv_data_90; // @[executor.scala 190:22]
  reg [7:0] phv_data_91; // @[executor.scala 190:22]
  reg [7:0] phv_data_92; // @[executor.scala 190:22]
  reg [7:0] phv_data_93; // @[executor.scala 190:22]
  reg [7:0] phv_data_94; // @[executor.scala 190:22]
  reg [7:0] phv_data_95; // @[executor.scala 190:22]
  reg [15:0] phv_header_0; // @[executor.scala 190:22]
  reg [15:0] phv_header_1; // @[executor.scala 190:22]
  reg [15:0] phv_header_2; // @[executor.scala 190:22]
  reg [15:0] phv_header_3; // @[executor.scala 190:22]
  reg [15:0] phv_header_4; // @[executor.scala 190:22]
  reg [15:0] phv_header_5; // @[executor.scala 190:22]
  reg [15:0] phv_header_6; // @[executor.scala 190:22]
  reg [15:0] phv_header_7; // @[executor.scala 190:22]
  reg [15:0] phv_header_8; // @[executor.scala 190:22]
  reg [15:0] phv_header_9; // @[executor.scala 190:22]
  reg [15:0] phv_header_10; // @[executor.scala 190:22]
  reg [15:0] phv_header_11; // @[executor.scala 190:22]
  reg [15:0] phv_header_12; // @[executor.scala 190:22]
  reg [15:0] phv_header_13; // @[executor.scala 190:22]
  reg [15:0] phv_header_14; // @[executor.scala 190:22]
  reg [15:0] phv_header_15; // @[executor.scala 190:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 190:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 190:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 190:22]
  reg [1:0] phv_next_processor_id; // @[executor.scala 190:22]
  reg [31:0] vliw_0; // @[executor.scala 194:23]
  reg [31:0] vliw_1; // @[executor.scala 194:23]
  reg [31:0] vliw_2; // @[executor.scala 194:23]
  reg [31:0] vliw_3; // @[executor.scala 194:23]
  reg [63:0] field_0; // @[executor.scala 198:24]
  reg [63:0] field_1; // @[executor.scala 198:24]
  reg [63:0] field_2; // @[executor.scala 198:24]
  reg [63:0] field_3; // @[executor.scala 198:24]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] imm_lo = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire [49:0] imm_hi = imm_lo[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] imm = {imm_hi,imm_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_field_out_0_T_1 = field_0 + imm; // @[executor.scala 208:45]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] imm_lo_1 = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire [49:0] imm_hi_1 = imm_lo_1[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] imm_1 = {imm_hi_1,imm_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _io_field_out_1_T_1 = field_1 + imm_1; // @[executor.scala 208:45]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] imm_lo_2 = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire [49:0] imm_hi_2 = imm_lo_2[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] imm_2 = {imm_hi_2,imm_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_field_out_2_T_1 = field_2 + imm_2; // @[executor.scala 208:45]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] imm_lo_3 = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire [49:0] imm_hi_3 = imm_lo_3[13] ? 50'h3ffffffffffff : 50'h0; // @[Bitwise.scala 72:12]
  wire [63:0] imm_3 = {imm_hi_3,imm_lo_3}; // @[Cat.scala 30:58]
  wire [63:0] _io_field_out_3_T_1 = field_3 + imm_3; // @[executor.scala 208:45]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 192:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 192:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 192:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 192:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 192:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 192:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 192:25]
  assign io_vliw_out_0 = vliw_0; // @[executor.scala 196:21]
  assign io_vliw_out_1 = vliw_1; // @[executor.scala 196:21]
  assign io_vliw_out_2 = vliw_2; // @[executor.scala 196:21]
  assign io_vliw_out_3 = vliw_3; // @[executor.scala 196:21]
  assign io_field_out_0 = 4'h8 == opcode ? _io_field_out_0_T_1 : field_0; // @[executor.scala 206:48 executor.scala 208:33 executor.scala 210:33]
  assign io_field_out_1 = 4'h8 == opcode_1 ? _io_field_out_1_T_1 : field_1; // @[executor.scala 206:48 executor.scala 208:33 executor.scala 210:33]
  assign io_field_out_2 = 4'h8 == opcode_2 ? _io_field_out_2_T_1 : field_2; // @[executor.scala 206:48 executor.scala 208:33 executor.scala 210:33]
  assign io_field_out_3 = 4'h8 == opcode_3 ? _io_field_out_3_T_1 : field_3; // @[executor.scala 206:48 executor.scala 208:33 executor.scala 210:33]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 191:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 191:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 191:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 191:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 191:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 191:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 191:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 191:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 191:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 191:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 191:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 191:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 191:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 191:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 191:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 191:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 191:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 191:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 191:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 191:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 191:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 191:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 191:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 191:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 191:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 191:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 191:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 191:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 191:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 191:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 191:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 191:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 191:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 191:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 191:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 191:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 191:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 191:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 191:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 191:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 191:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 191:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 191:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 191:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 191:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 191:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 191:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 191:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 191:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 191:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 191:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 191:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 191:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 191:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 191:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 191:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 191:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 191:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 191:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 191:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 191:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 191:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 191:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 191:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 191:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 191:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 191:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 191:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 191:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 191:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 191:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 191:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 191:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 191:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 191:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 191:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 191:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 191:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 191:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 191:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 191:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 191:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 191:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 191:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 191:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 191:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 191:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 191:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 191:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 191:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 191:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 191:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 191:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 191:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 191:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 191:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 191:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 191:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 191:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 191:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 191:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 191:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 191:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 191:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 191:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 191:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 191:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 191:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 191:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 191:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 191:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 191:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 191:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 191:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 191:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 191:13]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 195:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 195:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 195:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 195:14]
    field_0 <= io_field_in_0; // @[executor.scala 199:15]
    field_1 <= io_field_in_1; // @[executor.scala 199:15]
    field_2 <= io_field_in_2; // @[executor.scala 199:15]
    field_3 <= io_field_in_3; // @[executor.scala 199:15]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  vliw_0 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  vliw_1 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  vliw_2 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  vliw_3 = _RAND_119[31:0];
  _RAND_120 = {2{`RANDOM}};
  field_0 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  field_1 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  field_2 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  field_3 = _RAND_123[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PrimitiveGetWriteBackOffset(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [63:0] io_field_in_0,
  input  [63:0] io_field_in_1,
  input  [63:0] io_field_in_2,
  input  [63:0] io_field_in_3,
  output [7:0]  io_offset_out_0,
  output [7:0]  io_offset_out_1,
  output [7:0]  io_offset_out_2,
  output [7:0]  io_offset_out_3,
  output [7:0]  io_length_out_0,
  output [7:0]  io_length_out_1,
  output [7:0]  io_length_out_2,
  output [7:0]  io_length_out_3,
  output [63:0] io_field_out_0,
  output [63:0] io_field_out_1,
  output [63:0] io_field_out_2,
  output [63:0] io_field_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 227:22]
  reg [7:0] phv_data_1; // @[executor.scala 227:22]
  reg [7:0] phv_data_2; // @[executor.scala 227:22]
  reg [7:0] phv_data_3; // @[executor.scala 227:22]
  reg [7:0] phv_data_4; // @[executor.scala 227:22]
  reg [7:0] phv_data_5; // @[executor.scala 227:22]
  reg [7:0] phv_data_6; // @[executor.scala 227:22]
  reg [7:0] phv_data_7; // @[executor.scala 227:22]
  reg [7:0] phv_data_8; // @[executor.scala 227:22]
  reg [7:0] phv_data_9; // @[executor.scala 227:22]
  reg [7:0] phv_data_10; // @[executor.scala 227:22]
  reg [7:0] phv_data_11; // @[executor.scala 227:22]
  reg [7:0] phv_data_12; // @[executor.scala 227:22]
  reg [7:0] phv_data_13; // @[executor.scala 227:22]
  reg [7:0] phv_data_14; // @[executor.scala 227:22]
  reg [7:0] phv_data_15; // @[executor.scala 227:22]
  reg [7:0] phv_data_16; // @[executor.scala 227:22]
  reg [7:0] phv_data_17; // @[executor.scala 227:22]
  reg [7:0] phv_data_18; // @[executor.scala 227:22]
  reg [7:0] phv_data_19; // @[executor.scala 227:22]
  reg [7:0] phv_data_20; // @[executor.scala 227:22]
  reg [7:0] phv_data_21; // @[executor.scala 227:22]
  reg [7:0] phv_data_22; // @[executor.scala 227:22]
  reg [7:0] phv_data_23; // @[executor.scala 227:22]
  reg [7:0] phv_data_24; // @[executor.scala 227:22]
  reg [7:0] phv_data_25; // @[executor.scala 227:22]
  reg [7:0] phv_data_26; // @[executor.scala 227:22]
  reg [7:0] phv_data_27; // @[executor.scala 227:22]
  reg [7:0] phv_data_28; // @[executor.scala 227:22]
  reg [7:0] phv_data_29; // @[executor.scala 227:22]
  reg [7:0] phv_data_30; // @[executor.scala 227:22]
  reg [7:0] phv_data_31; // @[executor.scala 227:22]
  reg [7:0] phv_data_32; // @[executor.scala 227:22]
  reg [7:0] phv_data_33; // @[executor.scala 227:22]
  reg [7:0] phv_data_34; // @[executor.scala 227:22]
  reg [7:0] phv_data_35; // @[executor.scala 227:22]
  reg [7:0] phv_data_36; // @[executor.scala 227:22]
  reg [7:0] phv_data_37; // @[executor.scala 227:22]
  reg [7:0] phv_data_38; // @[executor.scala 227:22]
  reg [7:0] phv_data_39; // @[executor.scala 227:22]
  reg [7:0] phv_data_40; // @[executor.scala 227:22]
  reg [7:0] phv_data_41; // @[executor.scala 227:22]
  reg [7:0] phv_data_42; // @[executor.scala 227:22]
  reg [7:0] phv_data_43; // @[executor.scala 227:22]
  reg [7:0] phv_data_44; // @[executor.scala 227:22]
  reg [7:0] phv_data_45; // @[executor.scala 227:22]
  reg [7:0] phv_data_46; // @[executor.scala 227:22]
  reg [7:0] phv_data_47; // @[executor.scala 227:22]
  reg [7:0] phv_data_48; // @[executor.scala 227:22]
  reg [7:0] phv_data_49; // @[executor.scala 227:22]
  reg [7:0] phv_data_50; // @[executor.scala 227:22]
  reg [7:0] phv_data_51; // @[executor.scala 227:22]
  reg [7:0] phv_data_52; // @[executor.scala 227:22]
  reg [7:0] phv_data_53; // @[executor.scala 227:22]
  reg [7:0] phv_data_54; // @[executor.scala 227:22]
  reg [7:0] phv_data_55; // @[executor.scala 227:22]
  reg [7:0] phv_data_56; // @[executor.scala 227:22]
  reg [7:0] phv_data_57; // @[executor.scala 227:22]
  reg [7:0] phv_data_58; // @[executor.scala 227:22]
  reg [7:0] phv_data_59; // @[executor.scala 227:22]
  reg [7:0] phv_data_60; // @[executor.scala 227:22]
  reg [7:0] phv_data_61; // @[executor.scala 227:22]
  reg [7:0] phv_data_62; // @[executor.scala 227:22]
  reg [7:0] phv_data_63; // @[executor.scala 227:22]
  reg [7:0] phv_data_64; // @[executor.scala 227:22]
  reg [7:0] phv_data_65; // @[executor.scala 227:22]
  reg [7:0] phv_data_66; // @[executor.scala 227:22]
  reg [7:0] phv_data_67; // @[executor.scala 227:22]
  reg [7:0] phv_data_68; // @[executor.scala 227:22]
  reg [7:0] phv_data_69; // @[executor.scala 227:22]
  reg [7:0] phv_data_70; // @[executor.scala 227:22]
  reg [7:0] phv_data_71; // @[executor.scala 227:22]
  reg [7:0] phv_data_72; // @[executor.scala 227:22]
  reg [7:0] phv_data_73; // @[executor.scala 227:22]
  reg [7:0] phv_data_74; // @[executor.scala 227:22]
  reg [7:0] phv_data_75; // @[executor.scala 227:22]
  reg [7:0] phv_data_76; // @[executor.scala 227:22]
  reg [7:0] phv_data_77; // @[executor.scala 227:22]
  reg [7:0] phv_data_78; // @[executor.scala 227:22]
  reg [7:0] phv_data_79; // @[executor.scala 227:22]
  reg [7:0] phv_data_80; // @[executor.scala 227:22]
  reg [7:0] phv_data_81; // @[executor.scala 227:22]
  reg [7:0] phv_data_82; // @[executor.scala 227:22]
  reg [7:0] phv_data_83; // @[executor.scala 227:22]
  reg [7:0] phv_data_84; // @[executor.scala 227:22]
  reg [7:0] phv_data_85; // @[executor.scala 227:22]
  reg [7:0] phv_data_86; // @[executor.scala 227:22]
  reg [7:0] phv_data_87; // @[executor.scala 227:22]
  reg [7:0] phv_data_88; // @[executor.scala 227:22]
  reg [7:0] phv_data_89; // @[executor.scala 227:22]
  reg [7:0] phv_data_90; // @[executor.scala 227:22]
  reg [7:0] phv_data_91; // @[executor.scala 227:22]
  reg [7:0] phv_data_92; // @[executor.scala 227:22]
  reg [7:0] phv_data_93; // @[executor.scala 227:22]
  reg [7:0] phv_data_94; // @[executor.scala 227:22]
  reg [7:0] phv_data_95; // @[executor.scala 227:22]
  reg [15:0] phv_header_0; // @[executor.scala 227:22]
  reg [15:0] phv_header_1; // @[executor.scala 227:22]
  reg [15:0] phv_header_2; // @[executor.scala 227:22]
  reg [15:0] phv_header_3; // @[executor.scala 227:22]
  reg [15:0] phv_header_4; // @[executor.scala 227:22]
  reg [15:0] phv_header_5; // @[executor.scala 227:22]
  reg [15:0] phv_header_6; // @[executor.scala 227:22]
  reg [15:0] phv_header_7; // @[executor.scala 227:22]
  reg [15:0] phv_header_8; // @[executor.scala 227:22]
  reg [15:0] phv_header_9; // @[executor.scala 227:22]
  reg [15:0] phv_header_10; // @[executor.scala 227:22]
  reg [15:0] phv_header_11; // @[executor.scala 227:22]
  reg [15:0] phv_header_12; // @[executor.scala 227:22]
  reg [15:0] phv_header_13; // @[executor.scala 227:22]
  reg [15:0] phv_header_14; // @[executor.scala 227:22]
  reg [15:0] phv_header_15; // @[executor.scala 227:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 227:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 227:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 227:22]
  reg [1:0] phv_next_processor_id; // @[executor.scala 227:22]
  reg [31:0] vliw_0; // @[executor.scala 231:23]
  reg [31:0] vliw_1; // @[executor.scala 231:23]
  reg [31:0] vliw_2; // @[executor.scala 231:23]
  reg [31:0] vliw_3; // @[executor.scala 231:23]
  reg [63:0] field_0; // @[executor.scala 234:24]
  reg [63:0] field_1; // @[executor.scala 234:24]
  reg [63:0] field_2; // @[executor.scala 234:24]
  reg [63:0] field_3; // @[executor.scala 234:24]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1 = vliw_0[27:14]; // @[primitive.scala 10:44]
  wire [3:0] field_header_id = parameter_1[13:10]; // @[primitive.scala 27:52]
  wire [4:0] field_internal_offset = parameter_1[9:5]; // @[primitive.scala 28:52]
  wire [4:0] field_length = parameter_1[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_1 = 4'h1 == field_header_id ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_2 = 4'h2 == field_header_id ? phv_header_2 : _GEN_1; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_3 = 4'h3 == field_header_id ? phv_header_3 : _GEN_2; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_4 = 4'h4 == field_header_id ? phv_header_4 : _GEN_3; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_5 = 4'h5 == field_header_id ? phv_header_5 : _GEN_4; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_6 = 4'h6 == field_header_id ? phv_header_6 : _GEN_5; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_7 = 4'h7 == field_header_id ? phv_header_7 : _GEN_6; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_8 = 4'h8 == field_header_id ? phv_header_8 : _GEN_7; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_9 = 4'h9 == field_header_id ? phv_header_9 : _GEN_8; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_10 = 4'ha == field_header_id ? phv_header_10 : _GEN_9; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_11 = 4'hb == field_header_id ? phv_header_11 : _GEN_10; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_12 = 4'hc == field_header_id ? phv_header_12 : _GEN_11; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_13 = 4'hd == field_header_id ? phv_header_13 : _GEN_12; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_14 = 4'he == field_header_id ? phv_header_14 : _GEN_13; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_15 = 4'hf == field_header_id ? phv_header_15 : _GEN_14; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] field_header_offset = _GEN_15[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_68 = {{3'd0}, field_internal_offset}; // @[executor.scala 247:61]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_1 = vliw_1[27:14]; // @[primitive.scala 10:44]
  wire [3:0] field_header_id_1 = parameter_1_1[13:10]; // @[primitive.scala 27:52]
  wire [4:0] field_internal_offset_1 = parameter_1_1[9:5]; // @[primitive.scala 28:52]
  wire [4:0] field_length_1 = parameter_1_1[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_18 = 4'h1 == field_header_id_1 ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_19 = 4'h2 == field_header_id_1 ? phv_header_2 : _GEN_18; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_20 = 4'h3 == field_header_id_1 ? phv_header_3 : _GEN_19; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_21 = 4'h4 == field_header_id_1 ? phv_header_4 : _GEN_20; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_22 = 4'h5 == field_header_id_1 ? phv_header_5 : _GEN_21; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_23 = 4'h6 == field_header_id_1 ? phv_header_6 : _GEN_22; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_24 = 4'h7 == field_header_id_1 ? phv_header_7 : _GEN_23; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_25 = 4'h8 == field_header_id_1 ? phv_header_8 : _GEN_24; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_26 = 4'h9 == field_header_id_1 ? phv_header_9 : _GEN_25; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_27 = 4'ha == field_header_id_1 ? phv_header_10 : _GEN_26; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_28 = 4'hb == field_header_id_1 ? phv_header_11 : _GEN_27; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_29 = 4'hc == field_header_id_1 ? phv_header_12 : _GEN_28; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_30 = 4'hd == field_header_id_1 ? phv_header_13 : _GEN_29; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_31 = 4'he == field_header_id_1 ? phv_header_14 : _GEN_30; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_32 = 4'hf == field_header_id_1 ? phv_header_15 : _GEN_31; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] field_header_offset_1 = _GEN_32[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_69 = {{3'd0}, field_internal_offset_1}; // @[executor.scala 247:61]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_2 = vliw_2[27:14]; // @[primitive.scala 10:44]
  wire [3:0] field_header_id_2 = parameter_1_2[13:10]; // @[primitive.scala 27:52]
  wire [4:0] field_internal_offset_2 = parameter_1_2[9:5]; // @[primitive.scala 28:52]
  wire [4:0] field_length_2 = parameter_1_2[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_35 = 4'h1 == field_header_id_2 ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_36 = 4'h2 == field_header_id_2 ? phv_header_2 : _GEN_35; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_37 = 4'h3 == field_header_id_2 ? phv_header_3 : _GEN_36; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_38 = 4'h4 == field_header_id_2 ? phv_header_4 : _GEN_37; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_39 = 4'h5 == field_header_id_2 ? phv_header_5 : _GEN_38; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_40 = 4'h6 == field_header_id_2 ? phv_header_6 : _GEN_39; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_41 = 4'h7 == field_header_id_2 ? phv_header_7 : _GEN_40; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_42 = 4'h8 == field_header_id_2 ? phv_header_8 : _GEN_41; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_43 = 4'h9 == field_header_id_2 ? phv_header_9 : _GEN_42; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_44 = 4'ha == field_header_id_2 ? phv_header_10 : _GEN_43; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_45 = 4'hb == field_header_id_2 ? phv_header_11 : _GEN_44; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_46 = 4'hc == field_header_id_2 ? phv_header_12 : _GEN_45; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_47 = 4'hd == field_header_id_2 ? phv_header_13 : _GEN_46; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_48 = 4'he == field_header_id_2 ? phv_header_14 : _GEN_47; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_49 = 4'hf == field_header_id_2 ? phv_header_15 : _GEN_48; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] field_header_offset_2 = _GEN_49[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_70 = {{3'd0}, field_internal_offset_2}; // @[executor.scala 247:61]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_3 = vliw_3[27:14]; // @[primitive.scala 10:44]
  wire [3:0] field_header_id_3 = parameter_1_3[13:10]; // @[primitive.scala 27:52]
  wire [4:0] field_internal_offset_3 = parameter_1_3[9:5]; // @[primitive.scala 28:52]
  wire [4:0] field_length_3 = parameter_1_3[4:0]; // @[primitive.scala 29:52]
  wire [15:0] _GEN_52 = 4'h1 == field_header_id_3 ? phv_header_1 : phv_header_0; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_53 = 4'h2 == field_header_id_3 ? phv_header_2 : _GEN_52; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_54 = 4'h3 == field_header_id_3 ? phv_header_3 : _GEN_53; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_55 = 4'h4 == field_header_id_3 ? phv_header_4 : _GEN_54; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_56 = 4'h5 == field_header_id_3 ? phv_header_5 : _GEN_55; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_57 = 4'h6 == field_header_id_3 ? phv_header_6 : _GEN_56; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_58 = 4'h7 == field_header_id_3 ? phv_header_7 : _GEN_57; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_59 = 4'h8 == field_header_id_3 ? phv_header_8 : _GEN_58; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_60 = 4'h9 == field_header_id_3 ? phv_header_9 : _GEN_59; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_61 = 4'ha == field_header_id_3 ? phv_header_10 : _GEN_60; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_62 = 4'hb == field_header_id_3 ? phv_header_11 : _GEN_61; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_63 = 4'hc == field_header_id_3 ? phv_header_12 : _GEN_62; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_64 = 4'hd == field_header_id_3 ? phv_header_13 : _GEN_63; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_65 = 4'he == field_header_id_3 ? phv_header_14 : _GEN_64; // @[const.scala 29:43 const.scala 29:43]
  wire [15:0] _GEN_66 = 4'hf == field_header_id_3 ? phv_header_15 : _GEN_65; // @[const.scala 29:43 const.scala 29:43]
  wire [7:0] field_header_offset_3 = _GEN_66[15:8]; // @[const.scala 29:43]
  wire [7:0] _GEN_71 = {{3'd0}, field_internal_offset_3}; // @[executor.scala 247:61]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 229:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 229:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 229:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 229:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 229:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 229:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 229:25]
  assign io_offset_out_0 = field_header_offset + _GEN_68; // @[executor.scala 247:61]
  assign io_offset_out_1 = field_header_offset_1 + _GEN_69; // @[executor.scala 247:61]
  assign io_offset_out_2 = field_header_offset_2 + _GEN_70; // @[executor.scala 247:61]
  assign io_offset_out_3 = field_header_offset_3 + _GEN_71; // @[executor.scala 247:61]
  assign io_length_out_0 = 4'hf == opcode ? 8'h0 : {{3'd0}, field_length}; // @[executor.scala 250:48 executor.scala 251:34 executor.scala 253:34]
  assign io_length_out_1 = 4'hf == opcode_1 ? 8'h0 : {{3'd0}, field_length_1}; // @[executor.scala 250:48 executor.scala 251:34 executor.scala 253:34]
  assign io_length_out_2 = 4'hf == opcode_2 ? 8'h0 : {{3'd0}, field_length_2}; // @[executor.scala 250:48 executor.scala 251:34 executor.scala 253:34]
  assign io_length_out_3 = 4'hf == opcode_3 ? 8'h0 : {{3'd0}, field_length_3}; // @[executor.scala 250:48 executor.scala 251:34 executor.scala 253:34]
  assign io_field_out_0 = field_0; // @[executor.scala 236:22]
  assign io_field_out_1 = field_1; // @[executor.scala 236:22]
  assign io_field_out_2 = field_2; // @[executor.scala 236:22]
  assign io_field_out_3 = field_3; // @[executor.scala 236:22]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 228:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 228:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 228:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 228:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 228:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 228:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 228:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 228:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 228:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 228:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 228:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 228:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 228:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 228:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 228:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 228:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 228:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 228:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 228:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 228:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 228:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 228:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 228:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 228:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 228:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 228:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 228:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 228:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 228:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 228:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 228:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 228:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 228:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 228:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 228:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 228:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 228:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 228:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 228:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 228:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 228:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 228:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 228:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 228:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 228:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 228:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 228:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 228:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 228:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 228:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 228:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 228:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 228:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 228:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 228:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 228:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 228:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 228:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 228:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 228:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 228:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 228:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 228:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 228:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 228:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 228:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 228:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 228:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 228:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 228:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 228:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 228:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 228:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 228:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 228:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 228:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 228:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 228:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 228:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 228:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 228:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 228:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 228:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 228:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 228:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 228:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 228:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 228:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 228:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 228:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 228:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 228:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 228:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 228:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 228:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 228:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 228:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 228:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 228:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 228:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 228:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 228:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 228:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 228:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 228:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 228:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 228:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 228:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 228:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 228:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 228:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 228:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 228:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 228:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 228:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 228:13]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 232:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 232:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 232:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 232:14]
    field_0 <= io_field_in_0; // @[executor.scala 235:15]
    field_1 <= io_field_in_1; // @[executor.scala 235:15]
    field_2 <= io_field_in_2; // @[executor.scala 235:15]
    field_3 <= io_field_in_3; // @[executor.scala 235:15]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  vliw_0 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  vliw_1 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  vliw_2 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  vliw_3 = _RAND_119[31:0];
  _RAND_120 = {2{`RANDOM}};
  field_0 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  field_1 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  field_2 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  field_3 = _RAND_123[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PrimitiveWriteBack(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  input  [7:0]  io_offset_in_0,
  input  [7:0]  io_offset_in_1,
  input  [7:0]  io_offset_in_2,
  input  [7:0]  io_offset_in_3,
  input  [7:0]  io_length_in_0,
  input  [7:0]  io_length_in_1,
  input  [7:0]  io_length_in_2,
  input  [7:0]  io_length_in_3,
  input  [63:0] io_field_in_0,
  input  [63:0] io_field_in_1,
  input  [63:0] io_field_in_2,
  input  [63:0] io_field_in_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 268:22]
  reg [7:0] phv_data_1; // @[executor.scala 268:22]
  reg [7:0] phv_data_2; // @[executor.scala 268:22]
  reg [7:0] phv_data_3; // @[executor.scala 268:22]
  reg [7:0] phv_data_4; // @[executor.scala 268:22]
  reg [7:0] phv_data_5; // @[executor.scala 268:22]
  reg [7:0] phv_data_6; // @[executor.scala 268:22]
  reg [7:0] phv_data_7; // @[executor.scala 268:22]
  reg [7:0] phv_data_8; // @[executor.scala 268:22]
  reg [7:0] phv_data_9; // @[executor.scala 268:22]
  reg [7:0] phv_data_10; // @[executor.scala 268:22]
  reg [7:0] phv_data_11; // @[executor.scala 268:22]
  reg [7:0] phv_data_12; // @[executor.scala 268:22]
  reg [7:0] phv_data_13; // @[executor.scala 268:22]
  reg [7:0] phv_data_14; // @[executor.scala 268:22]
  reg [7:0] phv_data_15; // @[executor.scala 268:22]
  reg [7:0] phv_data_16; // @[executor.scala 268:22]
  reg [7:0] phv_data_17; // @[executor.scala 268:22]
  reg [7:0] phv_data_18; // @[executor.scala 268:22]
  reg [7:0] phv_data_19; // @[executor.scala 268:22]
  reg [7:0] phv_data_20; // @[executor.scala 268:22]
  reg [7:0] phv_data_21; // @[executor.scala 268:22]
  reg [7:0] phv_data_22; // @[executor.scala 268:22]
  reg [7:0] phv_data_23; // @[executor.scala 268:22]
  reg [7:0] phv_data_24; // @[executor.scala 268:22]
  reg [7:0] phv_data_25; // @[executor.scala 268:22]
  reg [7:0] phv_data_26; // @[executor.scala 268:22]
  reg [7:0] phv_data_27; // @[executor.scala 268:22]
  reg [7:0] phv_data_28; // @[executor.scala 268:22]
  reg [7:0] phv_data_29; // @[executor.scala 268:22]
  reg [7:0] phv_data_30; // @[executor.scala 268:22]
  reg [7:0] phv_data_31; // @[executor.scala 268:22]
  reg [7:0] phv_data_32; // @[executor.scala 268:22]
  reg [7:0] phv_data_33; // @[executor.scala 268:22]
  reg [7:0] phv_data_34; // @[executor.scala 268:22]
  reg [7:0] phv_data_35; // @[executor.scala 268:22]
  reg [7:0] phv_data_36; // @[executor.scala 268:22]
  reg [7:0] phv_data_37; // @[executor.scala 268:22]
  reg [7:0] phv_data_38; // @[executor.scala 268:22]
  reg [7:0] phv_data_39; // @[executor.scala 268:22]
  reg [7:0] phv_data_40; // @[executor.scala 268:22]
  reg [7:0] phv_data_41; // @[executor.scala 268:22]
  reg [7:0] phv_data_42; // @[executor.scala 268:22]
  reg [7:0] phv_data_43; // @[executor.scala 268:22]
  reg [7:0] phv_data_44; // @[executor.scala 268:22]
  reg [7:0] phv_data_45; // @[executor.scala 268:22]
  reg [7:0] phv_data_46; // @[executor.scala 268:22]
  reg [7:0] phv_data_47; // @[executor.scala 268:22]
  reg [7:0] phv_data_48; // @[executor.scala 268:22]
  reg [7:0] phv_data_49; // @[executor.scala 268:22]
  reg [7:0] phv_data_50; // @[executor.scala 268:22]
  reg [7:0] phv_data_51; // @[executor.scala 268:22]
  reg [7:0] phv_data_52; // @[executor.scala 268:22]
  reg [7:0] phv_data_53; // @[executor.scala 268:22]
  reg [7:0] phv_data_54; // @[executor.scala 268:22]
  reg [7:0] phv_data_55; // @[executor.scala 268:22]
  reg [7:0] phv_data_56; // @[executor.scala 268:22]
  reg [7:0] phv_data_57; // @[executor.scala 268:22]
  reg [7:0] phv_data_58; // @[executor.scala 268:22]
  reg [7:0] phv_data_59; // @[executor.scala 268:22]
  reg [7:0] phv_data_60; // @[executor.scala 268:22]
  reg [7:0] phv_data_61; // @[executor.scala 268:22]
  reg [7:0] phv_data_62; // @[executor.scala 268:22]
  reg [7:0] phv_data_63; // @[executor.scala 268:22]
  reg [7:0] phv_data_64; // @[executor.scala 268:22]
  reg [7:0] phv_data_65; // @[executor.scala 268:22]
  reg [7:0] phv_data_66; // @[executor.scala 268:22]
  reg [7:0] phv_data_67; // @[executor.scala 268:22]
  reg [7:0] phv_data_68; // @[executor.scala 268:22]
  reg [7:0] phv_data_69; // @[executor.scala 268:22]
  reg [7:0] phv_data_70; // @[executor.scala 268:22]
  reg [7:0] phv_data_71; // @[executor.scala 268:22]
  reg [7:0] phv_data_72; // @[executor.scala 268:22]
  reg [7:0] phv_data_73; // @[executor.scala 268:22]
  reg [7:0] phv_data_74; // @[executor.scala 268:22]
  reg [7:0] phv_data_75; // @[executor.scala 268:22]
  reg [7:0] phv_data_76; // @[executor.scala 268:22]
  reg [7:0] phv_data_77; // @[executor.scala 268:22]
  reg [7:0] phv_data_78; // @[executor.scala 268:22]
  reg [7:0] phv_data_79; // @[executor.scala 268:22]
  reg [7:0] phv_data_80; // @[executor.scala 268:22]
  reg [7:0] phv_data_81; // @[executor.scala 268:22]
  reg [7:0] phv_data_82; // @[executor.scala 268:22]
  reg [7:0] phv_data_83; // @[executor.scala 268:22]
  reg [7:0] phv_data_84; // @[executor.scala 268:22]
  reg [7:0] phv_data_85; // @[executor.scala 268:22]
  reg [7:0] phv_data_86; // @[executor.scala 268:22]
  reg [7:0] phv_data_87; // @[executor.scala 268:22]
  reg [7:0] phv_data_88; // @[executor.scala 268:22]
  reg [7:0] phv_data_89; // @[executor.scala 268:22]
  reg [7:0] phv_data_90; // @[executor.scala 268:22]
  reg [7:0] phv_data_91; // @[executor.scala 268:22]
  reg [7:0] phv_data_92; // @[executor.scala 268:22]
  reg [7:0] phv_data_93; // @[executor.scala 268:22]
  reg [7:0] phv_data_94; // @[executor.scala 268:22]
  reg [7:0] phv_data_95; // @[executor.scala 268:22]
  reg [15:0] phv_header_0; // @[executor.scala 268:22]
  reg [15:0] phv_header_1; // @[executor.scala 268:22]
  reg [15:0] phv_header_2; // @[executor.scala 268:22]
  reg [15:0] phv_header_3; // @[executor.scala 268:22]
  reg [15:0] phv_header_4; // @[executor.scala 268:22]
  reg [15:0] phv_header_5; // @[executor.scala 268:22]
  reg [15:0] phv_header_6; // @[executor.scala 268:22]
  reg [15:0] phv_header_7; // @[executor.scala 268:22]
  reg [15:0] phv_header_8; // @[executor.scala 268:22]
  reg [15:0] phv_header_9; // @[executor.scala 268:22]
  reg [15:0] phv_header_10; // @[executor.scala 268:22]
  reg [15:0] phv_header_11; // @[executor.scala 268:22]
  reg [15:0] phv_header_12; // @[executor.scala 268:22]
  reg [15:0] phv_header_13; // @[executor.scala 268:22]
  reg [15:0] phv_header_14; // @[executor.scala 268:22]
  reg [15:0] phv_header_15; // @[executor.scala 268:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 268:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 268:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 268:22]
  reg [1:0] phv_next_processor_id; // @[executor.scala 268:22]
  reg [7:0] offset_0; // @[executor.scala 272:25]
  reg [7:0] offset_1; // @[executor.scala 272:25]
  reg [7:0] offset_2; // @[executor.scala 272:25]
  reg [7:0] offset_3; // @[executor.scala 272:25]
  reg [7:0] length_0; // @[executor.scala 273:25]
  reg [7:0] length_1; // @[executor.scala 273:25]
  reg [7:0] length_2; // @[executor.scala 273:25]
  reg [7:0] length_3; // @[executor.scala 273:25]
  reg [63:0] field_0; // @[executor.scala 274:25]
  reg [63:0] field_1; // @[executor.scala 274:25]
  reg [63:0] field_2; // @[executor.scala 274:25]
  reg [63:0] field_3; // @[executor.scala 274:25]
  wire [7:0] field_byte = field_0[63:56]; // @[executor.scala 287:53]
  wire [8:0] _total_offset_T = {{1'd0}, offset_0}; // @[executor.scala 289:53]
  wire [7:0] total_offset = _total_offset_T[7:0]; // @[executor.scala 289:53]
  wire [7:0] _GEN_0 = 7'h0 == total_offset[6:0] ? field_byte : phv_data_0; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_1 = 7'h1 == total_offset[6:0] ? field_byte : phv_data_1; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_2 = 7'h2 == total_offset[6:0] ? field_byte : phv_data_2; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_3 = 7'h3 == total_offset[6:0] ? field_byte : phv_data_3; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_4 = 7'h4 == total_offset[6:0] ? field_byte : phv_data_4; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_5 = 7'h5 == total_offset[6:0] ? field_byte : phv_data_5; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_6 = 7'h6 == total_offset[6:0] ? field_byte : phv_data_6; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_7 = 7'h7 == total_offset[6:0] ? field_byte : phv_data_7; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_8 = 7'h8 == total_offset[6:0] ? field_byte : phv_data_8; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_9 = 7'h9 == total_offset[6:0] ? field_byte : phv_data_9; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_10 = 7'ha == total_offset[6:0] ? field_byte : phv_data_10; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_11 = 7'hb == total_offset[6:0] ? field_byte : phv_data_11; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_12 = 7'hc == total_offset[6:0] ? field_byte : phv_data_12; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_13 = 7'hd == total_offset[6:0] ? field_byte : phv_data_13; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_14 = 7'he == total_offset[6:0] ? field_byte : phv_data_14; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_15 = 7'hf == total_offset[6:0] ? field_byte : phv_data_15; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_16 = 7'h10 == total_offset[6:0] ? field_byte : phv_data_16; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_17 = 7'h11 == total_offset[6:0] ? field_byte : phv_data_17; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_18 = 7'h12 == total_offset[6:0] ? field_byte : phv_data_18; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_19 = 7'h13 == total_offset[6:0] ? field_byte : phv_data_19; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_20 = 7'h14 == total_offset[6:0] ? field_byte : phv_data_20; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_21 = 7'h15 == total_offset[6:0] ? field_byte : phv_data_21; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_22 = 7'h16 == total_offset[6:0] ? field_byte : phv_data_22; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_23 = 7'h17 == total_offset[6:0] ? field_byte : phv_data_23; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_24 = 7'h18 == total_offset[6:0] ? field_byte : phv_data_24; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_25 = 7'h19 == total_offset[6:0] ? field_byte : phv_data_25; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_26 = 7'h1a == total_offset[6:0] ? field_byte : phv_data_26; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_27 = 7'h1b == total_offset[6:0] ? field_byte : phv_data_27; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_28 = 7'h1c == total_offset[6:0] ? field_byte : phv_data_28; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_29 = 7'h1d == total_offset[6:0] ? field_byte : phv_data_29; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_30 = 7'h1e == total_offset[6:0] ? field_byte : phv_data_30; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_31 = 7'h1f == total_offset[6:0] ? field_byte : phv_data_31; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_32 = 7'h20 == total_offset[6:0] ? field_byte : phv_data_32; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_33 = 7'h21 == total_offset[6:0] ? field_byte : phv_data_33; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_34 = 7'h22 == total_offset[6:0] ? field_byte : phv_data_34; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_35 = 7'h23 == total_offset[6:0] ? field_byte : phv_data_35; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_36 = 7'h24 == total_offset[6:0] ? field_byte : phv_data_36; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_37 = 7'h25 == total_offset[6:0] ? field_byte : phv_data_37; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_38 = 7'h26 == total_offset[6:0] ? field_byte : phv_data_38; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_39 = 7'h27 == total_offset[6:0] ? field_byte : phv_data_39; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_40 = 7'h28 == total_offset[6:0] ? field_byte : phv_data_40; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_41 = 7'h29 == total_offset[6:0] ? field_byte : phv_data_41; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_42 = 7'h2a == total_offset[6:0] ? field_byte : phv_data_42; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_43 = 7'h2b == total_offset[6:0] ? field_byte : phv_data_43; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_44 = 7'h2c == total_offset[6:0] ? field_byte : phv_data_44; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_45 = 7'h2d == total_offset[6:0] ? field_byte : phv_data_45; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_46 = 7'h2e == total_offset[6:0] ? field_byte : phv_data_46; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_47 = 7'h2f == total_offset[6:0] ? field_byte : phv_data_47; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_48 = 7'h30 == total_offset[6:0] ? field_byte : phv_data_48; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_49 = 7'h31 == total_offset[6:0] ? field_byte : phv_data_49; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_50 = 7'h32 == total_offset[6:0] ? field_byte : phv_data_50; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_51 = 7'h33 == total_offset[6:0] ? field_byte : phv_data_51; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_52 = 7'h34 == total_offset[6:0] ? field_byte : phv_data_52; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_53 = 7'h35 == total_offset[6:0] ? field_byte : phv_data_53; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_54 = 7'h36 == total_offset[6:0] ? field_byte : phv_data_54; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_55 = 7'h37 == total_offset[6:0] ? field_byte : phv_data_55; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_56 = 7'h38 == total_offset[6:0] ? field_byte : phv_data_56; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_57 = 7'h39 == total_offset[6:0] ? field_byte : phv_data_57; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_58 = 7'h3a == total_offset[6:0] ? field_byte : phv_data_58; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_59 = 7'h3b == total_offset[6:0] ? field_byte : phv_data_59; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_60 = 7'h3c == total_offset[6:0] ? field_byte : phv_data_60; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_61 = 7'h3d == total_offset[6:0] ? field_byte : phv_data_61; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_62 = 7'h3e == total_offset[6:0] ? field_byte : phv_data_62; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_63 = 7'h3f == total_offset[6:0] ? field_byte : phv_data_63; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_64 = 7'h40 == total_offset[6:0] ? field_byte : phv_data_64; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_65 = 7'h41 == total_offset[6:0] ? field_byte : phv_data_65; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_66 = 7'h42 == total_offset[6:0] ? field_byte : phv_data_66; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_67 = 7'h43 == total_offset[6:0] ? field_byte : phv_data_67; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_68 = 7'h44 == total_offset[6:0] ? field_byte : phv_data_68; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_69 = 7'h45 == total_offset[6:0] ? field_byte : phv_data_69; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_70 = 7'h46 == total_offset[6:0] ? field_byte : phv_data_70; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_71 = 7'h47 == total_offset[6:0] ? field_byte : phv_data_71; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_72 = 7'h48 == total_offset[6:0] ? field_byte : phv_data_72; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_73 = 7'h49 == total_offset[6:0] ? field_byte : phv_data_73; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_74 = 7'h4a == total_offset[6:0] ? field_byte : phv_data_74; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_75 = 7'h4b == total_offset[6:0] ? field_byte : phv_data_75; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_76 = 7'h4c == total_offset[6:0] ? field_byte : phv_data_76; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_77 = 7'h4d == total_offset[6:0] ? field_byte : phv_data_77; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_78 = 7'h4e == total_offset[6:0] ? field_byte : phv_data_78; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_79 = 7'h4f == total_offset[6:0] ? field_byte : phv_data_79; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_80 = 7'h50 == total_offset[6:0] ? field_byte : phv_data_80; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_81 = 7'h51 == total_offset[6:0] ? field_byte : phv_data_81; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_82 = 7'h52 == total_offset[6:0] ? field_byte : phv_data_82; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_83 = 7'h53 == total_offset[6:0] ? field_byte : phv_data_83; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_84 = 7'h54 == total_offset[6:0] ? field_byte : phv_data_84; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_85 = 7'h55 == total_offset[6:0] ? field_byte : phv_data_85; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_86 = 7'h56 == total_offset[6:0] ? field_byte : phv_data_86; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_87 = 7'h57 == total_offset[6:0] ? field_byte : phv_data_87; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_88 = 7'h58 == total_offset[6:0] ? field_byte : phv_data_88; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_89 = 7'h59 == total_offset[6:0] ? field_byte : phv_data_89; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_90 = 7'h5a == total_offset[6:0] ? field_byte : phv_data_90; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_91 = 7'h5b == total_offset[6:0] ? field_byte : phv_data_91; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_92 = 7'h5c == total_offset[6:0] ? field_byte : phv_data_92; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_93 = 7'h5d == total_offset[6:0] ? field_byte : phv_data_93; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_94 = 7'h5e == total_offset[6:0] ? field_byte : phv_data_94; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_95 = 7'h5f == total_offset[6:0] ? field_byte : phv_data_95; // @[executor.scala 291:60 executor.scala 291:60 executor.scala 270:25]
  wire [7:0] _GEN_96 = 8'h0 < length_0 ? _GEN_0 : phv_data_0; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_97 = 8'h0 < length_0 ? _GEN_1 : phv_data_1; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_98 = 8'h0 < length_0 ? _GEN_2 : phv_data_2; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_99 = 8'h0 < length_0 ? _GEN_3 : phv_data_3; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_100 = 8'h0 < length_0 ? _GEN_4 : phv_data_4; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_101 = 8'h0 < length_0 ? _GEN_5 : phv_data_5; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_102 = 8'h0 < length_0 ? _GEN_6 : phv_data_6; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_103 = 8'h0 < length_0 ? _GEN_7 : phv_data_7; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_104 = 8'h0 < length_0 ? _GEN_8 : phv_data_8; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_105 = 8'h0 < length_0 ? _GEN_9 : phv_data_9; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_106 = 8'h0 < length_0 ? _GEN_10 : phv_data_10; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_107 = 8'h0 < length_0 ? _GEN_11 : phv_data_11; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_108 = 8'h0 < length_0 ? _GEN_12 : phv_data_12; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_109 = 8'h0 < length_0 ? _GEN_13 : phv_data_13; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_110 = 8'h0 < length_0 ? _GEN_14 : phv_data_14; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_111 = 8'h0 < length_0 ? _GEN_15 : phv_data_15; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_112 = 8'h0 < length_0 ? _GEN_16 : phv_data_16; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_113 = 8'h0 < length_0 ? _GEN_17 : phv_data_17; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_114 = 8'h0 < length_0 ? _GEN_18 : phv_data_18; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_115 = 8'h0 < length_0 ? _GEN_19 : phv_data_19; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_116 = 8'h0 < length_0 ? _GEN_20 : phv_data_20; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_117 = 8'h0 < length_0 ? _GEN_21 : phv_data_21; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_118 = 8'h0 < length_0 ? _GEN_22 : phv_data_22; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_119 = 8'h0 < length_0 ? _GEN_23 : phv_data_23; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_120 = 8'h0 < length_0 ? _GEN_24 : phv_data_24; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_121 = 8'h0 < length_0 ? _GEN_25 : phv_data_25; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_122 = 8'h0 < length_0 ? _GEN_26 : phv_data_26; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_123 = 8'h0 < length_0 ? _GEN_27 : phv_data_27; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_124 = 8'h0 < length_0 ? _GEN_28 : phv_data_28; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_125 = 8'h0 < length_0 ? _GEN_29 : phv_data_29; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_126 = 8'h0 < length_0 ? _GEN_30 : phv_data_30; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_127 = 8'h0 < length_0 ? _GEN_31 : phv_data_31; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_128 = 8'h0 < length_0 ? _GEN_32 : phv_data_32; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_129 = 8'h0 < length_0 ? _GEN_33 : phv_data_33; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_130 = 8'h0 < length_0 ? _GEN_34 : phv_data_34; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_131 = 8'h0 < length_0 ? _GEN_35 : phv_data_35; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_132 = 8'h0 < length_0 ? _GEN_36 : phv_data_36; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_133 = 8'h0 < length_0 ? _GEN_37 : phv_data_37; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_134 = 8'h0 < length_0 ? _GEN_38 : phv_data_38; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_135 = 8'h0 < length_0 ? _GEN_39 : phv_data_39; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_136 = 8'h0 < length_0 ? _GEN_40 : phv_data_40; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_137 = 8'h0 < length_0 ? _GEN_41 : phv_data_41; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_138 = 8'h0 < length_0 ? _GEN_42 : phv_data_42; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_139 = 8'h0 < length_0 ? _GEN_43 : phv_data_43; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_140 = 8'h0 < length_0 ? _GEN_44 : phv_data_44; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_141 = 8'h0 < length_0 ? _GEN_45 : phv_data_45; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_142 = 8'h0 < length_0 ? _GEN_46 : phv_data_46; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_143 = 8'h0 < length_0 ? _GEN_47 : phv_data_47; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_144 = 8'h0 < length_0 ? _GEN_48 : phv_data_48; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_145 = 8'h0 < length_0 ? _GEN_49 : phv_data_49; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_146 = 8'h0 < length_0 ? _GEN_50 : phv_data_50; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_147 = 8'h0 < length_0 ? _GEN_51 : phv_data_51; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_148 = 8'h0 < length_0 ? _GEN_52 : phv_data_52; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_149 = 8'h0 < length_0 ? _GEN_53 : phv_data_53; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_150 = 8'h0 < length_0 ? _GEN_54 : phv_data_54; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_151 = 8'h0 < length_0 ? _GEN_55 : phv_data_55; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_152 = 8'h0 < length_0 ? _GEN_56 : phv_data_56; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_153 = 8'h0 < length_0 ? _GEN_57 : phv_data_57; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_154 = 8'h0 < length_0 ? _GEN_58 : phv_data_58; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_155 = 8'h0 < length_0 ? _GEN_59 : phv_data_59; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_156 = 8'h0 < length_0 ? _GEN_60 : phv_data_60; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_157 = 8'h0 < length_0 ? _GEN_61 : phv_data_61; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_158 = 8'h0 < length_0 ? _GEN_62 : phv_data_62; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_159 = 8'h0 < length_0 ? _GEN_63 : phv_data_63; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_160 = 8'h0 < length_0 ? _GEN_64 : phv_data_64; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_161 = 8'h0 < length_0 ? _GEN_65 : phv_data_65; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_162 = 8'h0 < length_0 ? _GEN_66 : phv_data_66; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_163 = 8'h0 < length_0 ? _GEN_67 : phv_data_67; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_164 = 8'h0 < length_0 ? _GEN_68 : phv_data_68; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_165 = 8'h0 < length_0 ? _GEN_69 : phv_data_69; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_166 = 8'h0 < length_0 ? _GEN_70 : phv_data_70; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_167 = 8'h0 < length_0 ? _GEN_71 : phv_data_71; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_168 = 8'h0 < length_0 ? _GEN_72 : phv_data_72; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_169 = 8'h0 < length_0 ? _GEN_73 : phv_data_73; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_170 = 8'h0 < length_0 ? _GEN_74 : phv_data_74; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_171 = 8'h0 < length_0 ? _GEN_75 : phv_data_75; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_172 = 8'h0 < length_0 ? _GEN_76 : phv_data_76; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_173 = 8'h0 < length_0 ? _GEN_77 : phv_data_77; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_174 = 8'h0 < length_0 ? _GEN_78 : phv_data_78; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_175 = 8'h0 < length_0 ? _GEN_79 : phv_data_79; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_176 = 8'h0 < length_0 ? _GEN_80 : phv_data_80; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_177 = 8'h0 < length_0 ? _GEN_81 : phv_data_81; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_178 = 8'h0 < length_0 ? _GEN_82 : phv_data_82; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_179 = 8'h0 < length_0 ? _GEN_83 : phv_data_83; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_180 = 8'h0 < length_0 ? _GEN_84 : phv_data_84; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_181 = 8'h0 < length_0 ? _GEN_85 : phv_data_85; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_182 = 8'h0 < length_0 ? _GEN_86 : phv_data_86; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_183 = 8'h0 < length_0 ? _GEN_87 : phv_data_87; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_184 = 8'h0 < length_0 ? _GEN_88 : phv_data_88; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_185 = 8'h0 < length_0 ? _GEN_89 : phv_data_89; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_186 = 8'h0 < length_0 ? _GEN_90 : phv_data_90; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_187 = 8'h0 < length_0 ? _GEN_91 : phv_data_91; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_188 = 8'h0 < length_0 ? _GEN_92 : phv_data_92; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_189 = 8'h0 < length_0 ? _GEN_93 : phv_data_93; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_190 = 8'h0 < length_0 ? _GEN_94 : phv_data_94; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] _GEN_191 = 8'h0 < length_0 ? _GEN_95 : phv_data_95; // @[executor.scala 290:56 executor.scala 270:25]
  wire [7:0] field_byte_1 = field_0[55:48]; // @[executor.scala 287:53]
  wire [7:0] total_offset_1 = offset_0 + 8'h1; // @[executor.scala 289:53]
  wire [7:0] _GEN_192 = 7'h0 == total_offset_1[6:0] ? field_byte_1 : _GEN_96; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_193 = 7'h1 == total_offset_1[6:0] ? field_byte_1 : _GEN_97; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_194 = 7'h2 == total_offset_1[6:0] ? field_byte_1 : _GEN_98; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_195 = 7'h3 == total_offset_1[6:0] ? field_byte_1 : _GEN_99; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_196 = 7'h4 == total_offset_1[6:0] ? field_byte_1 : _GEN_100; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_197 = 7'h5 == total_offset_1[6:0] ? field_byte_1 : _GEN_101; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_198 = 7'h6 == total_offset_1[6:0] ? field_byte_1 : _GEN_102; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_199 = 7'h7 == total_offset_1[6:0] ? field_byte_1 : _GEN_103; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_200 = 7'h8 == total_offset_1[6:0] ? field_byte_1 : _GEN_104; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_201 = 7'h9 == total_offset_1[6:0] ? field_byte_1 : _GEN_105; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_202 = 7'ha == total_offset_1[6:0] ? field_byte_1 : _GEN_106; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_203 = 7'hb == total_offset_1[6:0] ? field_byte_1 : _GEN_107; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_204 = 7'hc == total_offset_1[6:0] ? field_byte_1 : _GEN_108; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_205 = 7'hd == total_offset_1[6:0] ? field_byte_1 : _GEN_109; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_206 = 7'he == total_offset_1[6:0] ? field_byte_1 : _GEN_110; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_207 = 7'hf == total_offset_1[6:0] ? field_byte_1 : _GEN_111; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_208 = 7'h10 == total_offset_1[6:0] ? field_byte_1 : _GEN_112; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_209 = 7'h11 == total_offset_1[6:0] ? field_byte_1 : _GEN_113; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_210 = 7'h12 == total_offset_1[6:0] ? field_byte_1 : _GEN_114; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_211 = 7'h13 == total_offset_1[6:0] ? field_byte_1 : _GEN_115; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_212 = 7'h14 == total_offset_1[6:0] ? field_byte_1 : _GEN_116; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_213 = 7'h15 == total_offset_1[6:0] ? field_byte_1 : _GEN_117; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_214 = 7'h16 == total_offset_1[6:0] ? field_byte_1 : _GEN_118; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_215 = 7'h17 == total_offset_1[6:0] ? field_byte_1 : _GEN_119; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_216 = 7'h18 == total_offset_1[6:0] ? field_byte_1 : _GEN_120; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_217 = 7'h19 == total_offset_1[6:0] ? field_byte_1 : _GEN_121; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_218 = 7'h1a == total_offset_1[6:0] ? field_byte_1 : _GEN_122; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_219 = 7'h1b == total_offset_1[6:0] ? field_byte_1 : _GEN_123; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_220 = 7'h1c == total_offset_1[6:0] ? field_byte_1 : _GEN_124; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_221 = 7'h1d == total_offset_1[6:0] ? field_byte_1 : _GEN_125; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_222 = 7'h1e == total_offset_1[6:0] ? field_byte_1 : _GEN_126; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_223 = 7'h1f == total_offset_1[6:0] ? field_byte_1 : _GEN_127; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_224 = 7'h20 == total_offset_1[6:0] ? field_byte_1 : _GEN_128; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_225 = 7'h21 == total_offset_1[6:0] ? field_byte_1 : _GEN_129; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_226 = 7'h22 == total_offset_1[6:0] ? field_byte_1 : _GEN_130; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_227 = 7'h23 == total_offset_1[6:0] ? field_byte_1 : _GEN_131; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_228 = 7'h24 == total_offset_1[6:0] ? field_byte_1 : _GEN_132; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_229 = 7'h25 == total_offset_1[6:0] ? field_byte_1 : _GEN_133; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_230 = 7'h26 == total_offset_1[6:0] ? field_byte_1 : _GEN_134; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_231 = 7'h27 == total_offset_1[6:0] ? field_byte_1 : _GEN_135; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_232 = 7'h28 == total_offset_1[6:0] ? field_byte_1 : _GEN_136; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_233 = 7'h29 == total_offset_1[6:0] ? field_byte_1 : _GEN_137; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_234 = 7'h2a == total_offset_1[6:0] ? field_byte_1 : _GEN_138; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_235 = 7'h2b == total_offset_1[6:0] ? field_byte_1 : _GEN_139; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_236 = 7'h2c == total_offset_1[6:0] ? field_byte_1 : _GEN_140; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_237 = 7'h2d == total_offset_1[6:0] ? field_byte_1 : _GEN_141; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_238 = 7'h2e == total_offset_1[6:0] ? field_byte_1 : _GEN_142; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_239 = 7'h2f == total_offset_1[6:0] ? field_byte_1 : _GEN_143; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_240 = 7'h30 == total_offset_1[6:0] ? field_byte_1 : _GEN_144; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_241 = 7'h31 == total_offset_1[6:0] ? field_byte_1 : _GEN_145; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_242 = 7'h32 == total_offset_1[6:0] ? field_byte_1 : _GEN_146; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_243 = 7'h33 == total_offset_1[6:0] ? field_byte_1 : _GEN_147; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_244 = 7'h34 == total_offset_1[6:0] ? field_byte_1 : _GEN_148; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_245 = 7'h35 == total_offset_1[6:0] ? field_byte_1 : _GEN_149; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_246 = 7'h36 == total_offset_1[6:0] ? field_byte_1 : _GEN_150; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_247 = 7'h37 == total_offset_1[6:0] ? field_byte_1 : _GEN_151; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_248 = 7'h38 == total_offset_1[6:0] ? field_byte_1 : _GEN_152; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_249 = 7'h39 == total_offset_1[6:0] ? field_byte_1 : _GEN_153; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_250 = 7'h3a == total_offset_1[6:0] ? field_byte_1 : _GEN_154; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_251 = 7'h3b == total_offset_1[6:0] ? field_byte_1 : _GEN_155; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_252 = 7'h3c == total_offset_1[6:0] ? field_byte_1 : _GEN_156; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_253 = 7'h3d == total_offset_1[6:0] ? field_byte_1 : _GEN_157; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_254 = 7'h3e == total_offset_1[6:0] ? field_byte_1 : _GEN_158; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_255 = 7'h3f == total_offset_1[6:0] ? field_byte_1 : _GEN_159; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_256 = 7'h40 == total_offset_1[6:0] ? field_byte_1 : _GEN_160; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_257 = 7'h41 == total_offset_1[6:0] ? field_byte_1 : _GEN_161; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_258 = 7'h42 == total_offset_1[6:0] ? field_byte_1 : _GEN_162; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_259 = 7'h43 == total_offset_1[6:0] ? field_byte_1 : _GEN_163; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_260 = 7'h44 == total_offset_1[6:0] ? field_byte_1 : _GEN_164; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_261 = 7'h45 == total_offset_1[6:0] ? field_byte_1 : _GEN_165; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_262 = 7'h46 == total_offset_1[6:0] ? field_byte_1 : _GEN_166; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_263 = 7'h47 == total_offset_1[6:0] ? field_byte_1 : _GEN_167; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_264 = 7'h48 == total_offset_1[6:0] ? field_byte_1 : _GEN_168; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_265 = 7'h49 == total_offset_1[6:0] ? field_byte_1 : _GEN_169; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_266 = 7'h4a == total_offset_1[6:0] ? field_byte_1 : _GEN_170; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_267 = 7'h4b == total_offset_1[6:0] ? field_byte_1 : _GEN_171; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_268 = 7'h4c == total_offset_1[6:0] ? field_byte_1 : _GEN_172; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_269 = 7'h4d == total_offset_1[6:0] ? field_byte_1 : _GEN_173; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_270 = 7'h4e == total_offset_1[6:0] ? field_byte_1 : _GEN_174; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_271 = 7'h4f == total_offset_1[6:0] ? field_byte_1 : _GEN_175; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_272 = 7'h50 == total_offset_1[6:0] ? field_byte_1 : _GEN_176; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_273 = 7'h51 == total_offset_1[6:0] ? field_byte_1 : _GEN_177; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_274 = 7'h52 == total_offset_1[6:0] ? field_byte_1 : _GEN_178; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_275 = 7'h53 == total_offset_1[6:0] ? field_byte_1 : _GEN_179; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_276 = 7'h54 == total_offset_1[6:0] ? field_byte_1 : _GEN_180; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_277 = 7'h55 == total_offset_1[6:0] ? field_byte_1 : _GEN_181; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_278 = 7'h56 == total_offset_1[6:0] ? field_byte_1 : _GEN_182; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_279 = 7'h57 == total_offset_1[6:0] ? field_byte_1 : _GEN_183; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_280 = 7'h58 == total_offset_1[6:0] ? field_byte_1 : _GEN_184; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_281 = 7'h59 == total_offset_1[6:0] ? field_byte_1 : _GEN_185; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_282 = 7'h5a == total_offset_1[6:0] ? field_byte_1 : _GEN_186; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_283 = 7'h5b == total_offset_1[6:0] ? field_byte_1 : _GEN_187; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_284 = 7'h5c == total_offset_1[6:0] ? field_byte_1 : _GEN_188; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_285 = 7'h5d == total_offset_1[6:0] ? field_byte_1 : _GEN_189; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_286 = 7'h5e == total_offset_1[6:0] ? field_byte_1 : _GEN_190; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_287 = 7'h5f == total_offset_1[6:0] ? field_byte_1 : _GEN_191; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_288 = 8'h1 < length_0 ? _GEN_192 : _GEN_96; // @[executor.scala 290:56]
  wire [7:0] _GEN_289 = 8'h1 < length_0 ? _GEN_193 : _GEN_97; // @[executor.scala 290:56]
  wire [7:0] _GEN_290 = 8'h1 < length_0 ? _GEN_194 : _GEN_98; // @[executor.scala 290:56]
  wire [7:0] _GEN_291 = 8'h1 < length_0 ? _GEN_195 : _GEN_99; // @[executor.scala 290:56]
  wire [7:0] _GEN_292 = 8'h1 < length_0 ? _GEN_196 : _GEN_100; // @[executor.scala 290:56]
  wire [7:0] _GEN_293 = 8'h1 < length_0 ? _GEN_197 : _GEN_101; // @[executor.scala 290:56]
  wire [7:0] _GEN_294 = 8'h1 < length_0 ? _GEN_198 : _GEN_102; // @[executor.scala 290:56]
  wire [7:0] _GEN_295 = 8'h1 < length_0 ? _GEN_199 : _GEN_103; // @[executor.scala 290:56]
  wire [7:0] _GEN_296 = 8'h1 < length_0 ? _GEN_200 : _GEN_104; // @[executor.scala 290:56]
  wire [7:0] _GEN_297 = 8'h1 < length_0 ? _GEN_201 : _GEN_105; // @[executor.scala 290:56]
  wire [7:0] _GEN_298 = 8'h1 < length_0 ? _GEN_202 : _GEN_106; // @[executor.scala 290:56]
  wire [7:0] _GEN_299 = 8'h1 < length_0 ? _GEN_203 : _GEN_107; // @[executor.scala 290:56]
  wire [7:0] _GEN_300 = 8'h1 < length_0 ? _GEN_204 : _GEN_108; // @[executor.scala 290:56]
  wire [7:0] _GEN_301 = 8'h1 < length_0 ? _GEN_205 : _GEN_109; // @[executor.scala 290:56]
  wire [7:0] _GEN_302 = 8'h1 < length_0 ? _GEN_206 : _GEN_110; // @[executor.scala 290:56]
  wire [7:0] _GEN_303 = 8'h1 < length_0 ? _GEN_207 : _GEN_111; // @[executor.scala 290:56]
  wire [7:0] _GEN_304 = 8'h1 < length_0 ? _GEN_208 : _GEN_112; // @[executor.scala 290:56]
  wire [7:0] _GEN_305 = 8'h1 < length_0 ? _GEN_209 : _GEN_113; // @[executor.scala 290:56]
  wire [7:0] _GEN_306 = 8'h1 < length_0 ? _GEN_210 : _GEN_114; // @[executor.scala 290:56]
  wire [7:0] _GEN_307 = 8'h1 < length_0 ? _GEN_211 : _GEN_115; // @[executor.scala 290:56]
  wire [7:0] _GEN_308 = 8'h1 < length_0 ? _GEN_212 : _GEN_116; // @[executor.scala 290:56]
  wire [7:0] _GEN_309 = 8'h1 < length_0 ? _GEN_213 : _GEN_117; // @[executor.scala 290:56]
  wire [7:0] _GEN_310 = 8'h1 < length_0 ? _GEN_214 : _GEN_118; // @[executor.scala 290:56]
  wire [7:0] _GEN_311 = 8'h1 < length_0 ? _GEN_215 : _GEN_119; // @[executor.scala 290:56]
  wire [7:0] _GEN_312 = 8'h1 < length_0 ? _GEN_216 : _GEN_120; // @[executor.scala 290:56]
  wire [7:0] _GEN_313 = 8'h1 < length_0 ? _GEN_217 : _GEN_121; // @[executor.scala 290:56]
  wire [7:0] _GEN_314 = 8'h1 < length_0 ? _GEN_218 : _GEN_122; // @[executor.scala 290:56]
  wire [7:0] _GEN_315 = 8'h1 < length_0 ? _GEN_219 : _GEN_123; // @[executor.scala 290:56]
  wire [7:0] _GEN_316 = 8'h1 < length_0 ? _GEN_220 : _GEN_124; // @[executor.scala 290:56]
  wire [7:0] _GEN_317 = 8'h1 < length_0 ? _GEN_221 : _GEN_125; // @[executor.scala 290:56]
  wire [7:0] _GEN_318 = 8'h1 < length_0 ? _GEN_222 : _GEN_126; // @[executor.scala 290:56]
  wire [7:0] _GEN_319 = 8'h1 < length_0 ? _GEN_223 : _GEN_127; // @[executor.scala 290:56]
  wire [7:0] _GEN_320 = 8'h1 < length_0 ? _GEN_224 : _GEN_128; // @[executor.scala 290:56]
  wire [7:0] _GEN_321 = 8'h1 < length_0 ? _GEN_225 : _GEN_129; // @[executor.scala 290:56]
  wire [7:0] _GEN_322 = 8'h1 < length_0 ? _GEN_226 : _GEN_130; // @[executor.scala 290:56]
  wire [7:0] _GEN_323 = 8'h1 < length_0 ? _GEN_227 : _GEN_131; // @[executor.scala 290:56]
  wire [7:0] _GEN_324 = 8'h1 < length_0 ? _GEN_228 : _GEN_132; // @[executor.scala 290:56]
  wire [7:0] _GEN_325 = 8'h1 < length_0 ? _GEN_229 : _GEN_133; // @[executor.scala 290:56]
  wire [7:0] _GEN_326 = 8'h1 < length_0 ? _GEN_230 : _GEN_134; // @[executor.scala 290:56]
  wire [7:0] _GEN_327 = 8'h1 < length_0 ? _GEN_231 : _GEN_135; // @[executor.scala 290:56]
  wire [7:0] _GEN_328 = 8'h1 < length_0 ? _GEN_232 : _GEN_136; // @[executor.scala 290:56]
  wire [7:0] _GEN_329 = 8'h1 < length_0 ? _GEN_233 : _GEN_137; // @[executor.scala 290:56]
  wire [7:0] _GEN_330 = 8'h1 < length_0 ? _GEN_234 : _GEN_138; // @[executor.scala 290:56]
  wire [7:0] _GEN_331 = 8'h1 < length_0 ? _GEN_235 : _GEN_139; // @[executor.scala 290:56]
  wire [7:0] _GEN_332 = 8'h1 < length_0 ? _GEN_236 : _GEN_140; // @[executor.scala 290:56]
  wire [7:0] _GEN_333 = 8'h1 < length_0 ? _GEN_237 : _GEN_141; // @[executor.scala 290:56]
  wire [7:0] _GEN_334 = 8'h1 < length_0 ? _GEN_238 : _GEN_142; // @[executor.scala 290:56]
  wire [7:0] _GEN_335 = 8'h1 < length_0 ? _GEN_239 : _GEN_143; // @[executor.scala 290:56]
  wire [7:0] _GEN_336 = 8'h1 < length_0 ? _GEN_240 : _GEN_144; // @[executor.scala 290:56]
  wire [7:0] _GEN_337 = 8'h1 < length_0 ? _GEN_241 : _GEN_145; // @[executor.scala 290:56]
  wire [7:0] _GEN_338 = 8'h1 < length_0 ? _GEN_242 : _GEN_146; // @[executor.scala 290:56]
  wire [7:0] _GEN_339 = 8'h1 < length_0 ? _GEN_243 : _GEN_147; // @[executor.scala 290:56]
  wire [7:0] _GEN_340 = 8'h1 < length_0 ? _GEN_244 : _GEN_148; // @[executor.scala 290:56]
  wire [7:0] _GEN_341 = 8'h1 < length_0 ? _GEN_245 : _GEN_149; // @[executor.scala 290:56]
  wire [7:0] _GEN_342 = 8'h1 < length_0 ? _GEN_246 : _GEN_150; // @[executor.scala 290:56]
  wire [7:0] _GEN_343 = 8'h1 < length_0 ? _GEN_247 : _GEN_151; // @[executor.scala 290:56]
  wire [7:0] _GEN_344 = 8'h1 < length_0 ? _GEN_248 : _GEN_152; // @[executor.scala 290:56]
  wire [7:0] _GEN_345 = 8'h1 < length_0 ? _GEN_249 : _GEN_153; // @[executor.scala 290:56]
  wire [7:0] _GEN_346 = 8'h1 < length_0 ? _GEN_250 : _GEN_154; // @[executor.scala 290:56]
  wire [7:0] _GEN_347 = 8'h1 < length_0 ? _GEN_251 : _GEN_155; // @[executor.scala 290:56]
  wire [7:0] _GEN_348 = 8'h1 < length_0 ? _GEN_252 : _GEN_156; // @[executor.scala 290:56]
  wire [7:0] _GEN_349 = 8'h1 < length_0 ? _GEN_253 : _GEN_157; // @[executor.scala 290:56]
  wire [7:0] _GEN_350 = 8'h1 < length_0 ? _GEN_254 : _GEN_158; // @[executor.scala 290:56]
  wire [7:0] _GEN_351 = 8'h1 < length_0 ? _GEN_255 : _GEN_159; // @[executor.scala 290:56]
  wire [7:0] _GEN_352 = 8'h1 < length_0 ? _GEN_256 : _GEN_160; // @[executor.scala 290:56]
  wire [7:0] _GEN_353 = 8'h1 < length_0 ? _GEN_257 : _GEN_161; // @[executor.scala 290:56]
  wire [7:0] _GEN_354 = 8'h1 < length_0 ? _GEN_258 : _GEN_162; // @[executor.scala 290:56]
  wire [7:0] _GEN_355 = 8'h1 < length_0 ? _GEN_259 : _GEN_163; // @[executor.scala 290:56]
  wire [7:0] _GEN_356 = 8'h1 < length_0 ? _GEN_260 : _GEN_164; // @[executor.scala 290:56]
  wire [7:0] _GEN_357 = 8'h1 < length_0 ? _GEN_261 : _GEN_165; // @[executor.scala 290:56]
  wire [7:0] _GEN_358 = 8'h1 < length_0 ? _GEN_262 : _GEN_166; // @[executor.scala 290:56]
  wire [7:0] _GEN_359 = 8'h1 < length_0 ? _GEN_263 : _GEN_167; // @[executor.scala 290:56]
  wire [7:0] _GEN_360 = 8'h1 < length_0 ? _GEN_264 : _GEN_168; // @[executor.scala 290:56]
  wire [7:0] _GEN_361 = 8'h1 < length_0 ? _GEN_265 : _GEN_169; // @[executor.scala 290:56]
  wire [7:0] _GEN_362 = 8'h1 < length_0 ? _GEN_266 : _GEN_170; // @[executor.scala 290:56]
  wire [7:0] _GEN_363 = 8'h1 < length_0 ? _GEN_267 : _GEN_171; // @[executor.scala 290:56]
  wire [7:0] _GEN_364 = 8'h1 < length_0 ? _GEN_268 : _GEN_172; // @[executor.scala 290:56]
  wire [7:0] _GEN_365 = 8'h1 < length_0 ? _GEN_269 : _GEN_173; // @[executor.scala 290:56]
  wire [7:0] _GEN_366 = 8'h1 < length_0 ? _GEN_270 : _GEN_174; // @[executor.scala 290:56]
  wire [7:0] _GEN_367 = 8'h1 < length_0 ? _GEN_271 : _GEN_175; // @[executor.scala 290:56]
  wire [7:0] _GEN_368 = 8'h1 < length_0 ? _GEN_272 : _GEN_176; // @[executor.scala 290:56]
  wire [7:0] _GEN_369 = 8'h1 < length_0 ? _GEN_273 : _GEN_177; // @[executor.scala 290:56]
  wire [7:0] _GEN_370 = 8'h1 < length_0 ? _GEN_274 : _GEN_178; // @[executor.scala 290:56]
  wire [7:0] _GEN_371 = 8'h1 < length_0 ? _GEN_275 : _GEN_179; // @[executor.scala 290:56]
  wire [7:0] _GEN_372 = 8'h1 < length_0 ? _GEN_276 : _GEN_180; // @[executor.scala 290:56]
  wire [7:0] _GEN_373 = 8'h1 < length_0 ? _GEN_277 : _GEN_181; // @[executor.scala 290:56]
  wire [7:0] _GEN_374 = 8'h1 < length_0 ? _GEN_278 : _GEN_182; // @[executor.scala 290:56]
  wire [7:0] _GEN_375 = 8'h1 < length_0 ? _GEN_279 : _GEN_183; // @[executor.scala 290:56]
  wire [7:0] _GEN_376 = 8'h1 < length_0 ? _GEN_280 : _GEN_184; // @[executor.scala 290:56]
  wire [7:0] _GEN_377 = 8'h1 < length_0 ? _GEN_281 : _GEN_185; // @[executor.scala 290:56]
  wire [7:0] _GEN_378 = 8'h1 < length_0 ? _GEN_282 : _GEN_186; // @[executor.scala 290:56]
  wire [7:0] _GEN_379 = 8'h1 < length_0 ? _GEN_283 : _GEN_187; // @[executor.scala 290:56]
  wire [7:0] _GEN_380 = 8'h1 < length_0 ? _GEN_284 : _GEN_188; // @[executor.scala 290:56]
  wire [7:0] _GEN_381 = 8'h1 < length_0 ? _GEN_285 : _GEN_189; // @[executor.scala 290:56]
  wire [7:0] _GEN_382 = 8'h1 < length_0 ? _GEN_286 : _GEN_190; // @[executor.scala 290:56]
  wire [7:0] _GEN_383 = 8'h1 < length_0 ? _GEN_287 : _GEN_191; // @[executor.scala 290:56]
  wire [7:0] field_byte_2 = field_0[47:40]; // @[executor.scala 287:53]
  wire [7:0] total_offset_2 = offset_0 + 8'h2; // @[executor.scala 289:53]
  wire [7:0] _GEN_384 = 7'h0 == total_offset_2[6:0] ? field_byte_2 : _GEN_288; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_385 = 7'h1 == total_offset_2[6:0] ? field_byte_2 : _GEN_289; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_386 = 7'h2 == total_offset_2[6:0] ? field_byte_2 : _GEN_290; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_387 = 7'h3 == total_offset_2[6:0] ? field_byte_2 : _GEN_291; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_388 = 7'h4 == total_offset_2[6:0] ? field_byte_2 : _GEN_292; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_389 = 7'h5 == total_offset_2[6:0] ? field_byte_2 : _GEN_293; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_390 = 7'h6 == total_offset_2[6:0] ? field_byte_2 : _GEN_294; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_391 = 7'h7 == total_offset_2[6:0] ? field_byte_2 : _GEN_295; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_392 = 7'h8 == total_offset_2[6:0] ? field_byte_2 : _GEN_296; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_393 = 7'h9 == total_offset_2[6:0] ? field_byte_2 : _GEN_297; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_394 = 7'ha == total_offset_2[6:0] ? field_byte_2 : _GEN_298; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_395 = 7'hb == total_offset_2[6:0] ? field_byte_2 : _GEN_299; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_396 = 7'hc == total_offset_2[6:0] ? field_byte_2 : _GEN_300; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_397 = 7'hd == total_offset_2[6:0] ? field_byte_2 : _GEN_301; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_398 = 7'he == total_offset_2[6:0] ? field_byte_2 : _GEN_302; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_399 = 7'hf == total_offset_2[6:0] ? field_byte_2 : _GEN_303; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_400 = 7'h10 == total_offset_2[6:0] ? field_byte_2 : _GEN_304; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_401 = 7'h11 == total_offset_2[6:0] ? field_byte_2 : _GEN_305; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_402 = 7'h12 == total_offset_2[6:0] ? field_byte_2 : _GEN_306; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_403 = 7'h13 == total_offset_2[6:0] ? field_byte_2 : _GEN_307; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_404 = 7'h14 == total_offset_2[6:0] ? field_byte_2 : _GEN_308; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_405 = 7'h15 == total_offset_2[6:0] ? field_byte_2 : _GEN_309; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_406 = 7'h16 == total_offset_2[6:0] ? field_byte_2 : _GEN_310; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_407 = 7'h17 == total_offset_2[6:0] ? field_byte_2 : _GEN_311; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_408 = 7'h18 == total_offset_2[6:0] ? field_byte_2 : _GEN_312; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_409 = 7'h19 == total_offset_2[6:0] ? field_byte_2 : _GEN_313; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_410 = 7'h1a == total_offset_2[6:0] ? field_byte_2 : _GEN_314; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_411 = 7'h1b == total_offset_2[6:0] ? field_byte_2 : _GEN_315; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_412 = 7'h1c == total_offset_2[6:0] ? field_byte_2 : _GEN_316; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_413 = 7'h1d == total_offset_2[6:0] ? field_byte_2 : _GEN_317; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_414 = 7'h1e == total_offset_2[6:0] ? field_byte_2 : _GEN_318; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_415 = 7'h1f == total_offset_2[6:0] ? field_byte_2 : _GEN_319; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_416 = 7'h20 == total_offset_2[6:0] ? field_byte_2 : _GEN_320; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_417 = 7'h21 == total_offset_2[6:0] ? field_byte_2 : _GEN_321; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_418 = 7'h22 == total_offset_2[6:0] ? field_byte_2 : _GEN_322; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_419 = 7'h23 == total_offset_2[6:0] ? field_byte_2 : _GEN_323; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_420 = 7'h24 == total_offset_2[6:0] ? field_byte_2 : _GEN_324; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_421 = 7'h25 == total_offset_2[6:0] ? field_byte_2 : _GEN_325; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_422 = 7'h26 == total_offset_2[6:0] ? field_byte_2 : _GEN_326; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_423 = 7'h27 == total_offset_2[6:0] ? field_byte_2 : _GEN_327; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_424 = 7'h28 == total_offset_2[6:0] ? field_byte_2 : _GEN_328; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_425 = 7'h29 == total_offset_2[6:0] ? field_byte_2 : _GEN_329; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_426 = 7'h2a == total_offset_2[6:0] ? field_byte_2 : _GEN_330; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_427 = 7'h2b == total_offset_2[6:0] ? field_byte_2 : _GEN_331; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_428 = 7'h2c == total_offset_2[6:0] ? field_byte_2 : _GEN_332; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_429 = 7'h2d == total_offset_2[6:0] ? field_byte_2 : _GEN_333; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_430 = 7'h2e == total_offset_2[6:0] ? field_byte_2 : _GEN_334; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_431 = 7'h2f == total_offset_2[6:0] ? field_byte_2 : _GEN_335; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_432 = 7'h30 == total_offset_2[6:0] ? field_byte_2 : _GEN_336; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_433 = 7'h31 == total_offset_2[6:0] ? field_byte_2 : _GEN_337; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_434 = 7'h32 == total_offset_2[6:0] ? field_byte_2 : _GEN_338; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_435 = 7'h33 == total_offset_2[6:0] ? field_byte_2 : _GEN_339; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_436 = 7'h34 == total_offset_2[6:0] ? field_byte_2 : _GEN_340; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_437 = 7'h35 == total_offset_2[6:0] ? field_byte_2 : _GEN_341; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_438 = 7'h36 == total_offset_2[6:0] ? field_byte_2 : _GEN_342; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_439 = 7'h37 == total_offset_2[6:0] ? field_byte_2 : _GEN_343; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_440 = 7'h38 == total_offset_2[6:0] ? field_byte_2 : _GEN_344; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_441 = 7'h39 == total_offset_2[6:0] ? field_byte_2 : _GEN_345; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_442 = 7'h3a == total_offset_2[6:0] ? field_byte_2 : _GEN_346; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_443 = 7'h3b == total_offset_2[6:0] ? field_byte_2 : _GEN_347; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_444 = 7'h3c == total_offset_2[6:0] ? field_byte_2 : _GEN_348; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_445 = 7'h3d == total_offset_2[6:0] ? field_byte_2 : _GEN_349; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_446 = 7'h3e == total_offset_2[6:0] ? field_byte_2 : _GEN_350; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_447 = 7'h3f == total_offset_2[6:0] ? field_byte_2 : _GEN_351; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_448 = 7'h40 == total_offset_2[6:0] ? field_byte_2 : _GEN_352; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_449 = 7'h41 == total_offset_2[6:0] ? field_byte_2 : _GEN_353; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_450 = 7'h42 == total_offset_2[6:0] ? field_byte_2 : _GEN_354; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_451 = 7'h43 == total_offset_2[6:0] ? field_byte_2 : _GEN_355; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_452 = 7'h44 == total_offset_2[6:0] ? field_byte_2 : _GEN_356; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_453 = 7'h45 == total_offset_2[6:0] ? field_byte_2 : _GEN_357; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_454 = 7'h46 == total_offset_2[6:0] ? field_byte_2 : _GEN_358; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_455 = 7'h47 == total_offset_2[6:0] ? field_byte_2 : _GEN_359; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_456 = 7'h48 == total_offset_2[6:0] ? field_byte_2 : _GEN_360; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_457 = 7'h49 == total_offset_2[6:0] ? field_byte_2 : _GEN_361; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_458 = 7'h4a == total_offset_2[6:0] ? field_byte_2 : _GEN_362; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_459 = 7'h4b == total_offset_2[6:0] ? field_byte_2 : _GEN_363; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_460 = 7'h4c == total_offset_2[6:0] ? field_byte_2 : _GEN_364; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_461 = 7'h4d == total_offset_2[6:0] ? field_byte_2 : _GEN_365; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_462 = 7'h4e == total_offset_2[6:0] ? field_byte_2 : _GEN_366; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_463 = 7'h4f == total_offset_2[6:0] ? field_byte_2 : _GEN_367; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_464 = 7'h50 == total_offset_2[6:0] ? field_byte_2 : _GEN_368; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_465 = 7'h51 == total_offset_2[6:0] ? field_byte_2 : _GEN_369; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_466 = 7'h52 == total_offset_2[6:0] ? field_byte_2 : _GEN_370; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_467 = 7'h53 == total_offset_2[6:0] ? field_byte_2 : _GEN_371; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_468 = 7'h54 == total_offset_2[6:0] ? field_byte_2 : _GEN_372; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_469 = 7'h55 == total_offset_2[6:0] ? field_byte_2 : _GEN_373; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_470 = 7'h56 == total_offset_2[6:0] ? field_byte_2 : _GEN_374; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_471 = 7'h57 == total_offset_2[6:0] ? field_byte_2 : _GEN_375; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_472 = 7'h58 == total_offset_2[6:0] ? field_byte_2 : _GEN_376; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_473 = 7'h59 == total_offset_2[6:0] ? field_byte_2 : _GEN_377; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_474 = 7'h5a == total_offset_2[6:0] ? field_byte_2 : _GEN_378; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_475 = 7'h5b == total_offset_2[6:0] ? field_byte_2 : _GEN_379; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_476 = 7'h5c == total_offset_2[6:0] ? field_byte_2 : _GEN_380; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_477 = 7'h5d == total_offset_2[6:0] ? field_byte_2 : _GEN_381; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_478 = 7'h5e == total_offset_2[6:0] ? field_byte_2 : _GEN_382; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_479 = 7'h5f == total_offset_2[6:0] ? field_byte_2 : _GEN_383; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_480 = 8'h2 < length_0 ? _GEN_384 : _GEN_288; // @[executor.scala 290:56]
  wire [7:0] _GEN_481 = 8'h2 < length_0 ? _GEN_385 : _GEN_289; // @[executor.scala 290:56]
  wire [7:0] _GEN_482 = 8'h2 < length_0 ? _GEN_386 : _GEN_290; // @[executor.scala 290:56]
  wire [7:0] _GEN_483 = 8'h2 < length_0 ? _GEN_387 : _GEN_291; // @[executor.scala 290:56]
  wire [7:0] _GEN_484 = 8'h2 < length_0 ? _GEN_388 : _GEN_292; // @[executor.scala 290:56]
  wire [7:0] _GEN_485 = 8'h2 < length_0 ? _GEN_389 : _GEN_293; // @[executor.scala 290:56]
  wire [7:0] _GEN_486 = 8'h2 < length_0 ? _GEN_390 : _GEN_294; // @[executor.scala 290:56]
  wire [7:0] _GEN_487 = 8'h2 < length_0 ? _GEN_391 : _GEN_295; // @[executor.scala 290:56]
  wire [7:0] _GEN_488 = 8'h2 < length_0 ? _GEN_392 : _GEN_296; // @[executor.scala 290:56]
  wire [7:0] _GEN_489 = 8'h2 < length_0 ? _GEN_393 : _GEN_297; // @[executor.scala 290:56]
  wire [7:0] _GEN_490 = 8'h2 < length_0 ? _GEN_394 : _GEN_298; // @[executor.scala 290:56]
  wire [7:0] _GEN_491 = 8'h2 < length_0 ? _GEN_395 : _GEN_299; // @[executor.scala 290:56]
  wire [7:0] _GEN_492 = 8'h2 < length_0 ? _GEN_396 : _GEN_300; // @[executor.scala 290:56]
  wire [7:0] _GEN_493 = 8'h2 < length_0 ? _GEN_397 : _GEN_301; // @[executor.scala 290:56]
  wire [7:0] _GEN_494 = 8'h2 < length_0 ? _GEN_398 : _GEN_302; // @[executor.scala 290:56]
  wire [7:0] _GEN_495 = 8'h2 < length_0 ? _GEN_399 : _GEN_303; // @[executor.scala 290:56]
  wire [7:0] _GEN_496 = 8'h2 < length_0 ? _GEN_400 : _GEN_304; // @[executor.scala 290:56]
  wire [7:0] _GEN_497 = 8'h2 < length_0 ? _GEN_401 : _GEN_305; // @[executor.scala 290:56]
  wire [7:0] _GEN_498 = 8'h2 < length_0 ? _GEN_402 : _GEN_306; // @[executor.scala 290:56]
  wire [7:0] _GEN_499 = 8'h2 < length_0 ? _GEN_403 : _GEN_307; // @[executor.scala 290:56]
  wire [7:0] _GEN_500 = 8'h2 < length_0 ? _GEN_404 : _GEN_308; // @[executor.scala 290:56]
  wire [7:0] _GEN_501 = 8'h2 < length_0 ? _GEN_405 : _GEN_309; // @[executor.scala 290:56]
  wire [7:0] _GEN_502 = 8'h2 < length_0 ? _GEN_406 : _GEN_310; // @[executor.scala 290:56]
  wire [7:0] _GEN_503 = 8'h2 < length_0 ? _GEN_407 : _GEN_311; // @[executor.scala 290:56]
  wire [7:0] _GEN_504 = 8'h2 < length_0 ? _GEN_408 : _GEN_312; // @[executor.scala 290:56]
  wire [7:0] _GEN_505 = 8'h2 < length_0 ? _GEN_409 : _GEN_313; // @[executor.scala 290:56]
  wire [7:0] _GEN_506 = 8'h2 < length_0 ? _GEN_410 : _GEN_314; // @[executor.scala 290:56]
  wire [7:0] _GEN_507 = 8'h2 < length_0 ? _GEN_411 : _GEN_315; // @[executor.scala 290:56]
  wire [7:0] _GEN_508 = 8'h2 < length_0 ? _GEN_412 : _GEN_316; // @[executor.scala 290:56]
  wire [7:0] _GEN_509 = 8'h2 < length_0 ? _GEN_413 : _GEN_317; // @[executor.scala 290:56]
  wire [7:0] _GEN_510 = 8'h2 < length_0 ? _GEN_414 : _GEN_318; // @[executor.scala 290:56]
  wire [7:0] _GEN_511 = 8'h2 < length_0 ? _GEN_415 : _GEN_319; // @[executor.scala 290:56]
  wire [7:0] _GEN_512 = 8'h2 < length_0 ? _GEN_416 : _GEN_320; // @[executor.scala 290:56]
  wire [7:0] _GEN_513 = 8'h2 < length_0 ? _GEN_417 : _GEN_321; // @[executor.scala 290:56]
  wire [7:0] _GEN_514 = 8'h2 < length_0 ? _GEN_418 : _GEN_322; // @[executor.scala 290:56]
  wire [7:0] _GEN_515 = 8'h2 < length_0 ? _GEN_419 : _GEN_323; // @[executor.scala 290:56]
  wire [7:0] _GEN_516 = 8'h2 < length_0 ? _GEN_420 : _GEN_324; // @[executor.scala 290:56]
  wire [7:0] _GEN_517 = 8'h2 < length_0 ? _GEN_421 : _GEN_325; // @[executor.scala 290:56]
  wire [7:0] _GEN_518 = 8'h2 < length_0 ? _GEN_422 : _GEN_326; // @[executor.scala 290:56]
  wire [7:0] _GEN_519 = 8'h2 < length_0 ? _GEN_423 : _GEN_327; // @[executor.scala 290:56]
  wire [7:0] _GEN_520 = 8'h2 < length_0 ? _GEN_424 : _GEN_328; // @[executor.scala 290:56]
  wire [7:0] _GEN_521 = 8'h2 < length_0 ? _GEN_425 : _GEN_329; // @[executor.scala 290:56]
  wire [7:0] _GEN_522 = 8'h2 < length_0 ? _GEN_426 : _GEN_330; // @[executor.scala 290:56]
  wire [7:0] _GEN_523 = 8'h2 < length_0 ? _GEN_427 : _GEN_331; // @[executor.scala 290:56]
  wire [7:0] _GEN_524 = 8'h2 < length_0 ? _GEN_428 : _GEN_332; // @[executor.scala 290:56]
  wire [7:0] _GEN_525 = 8'h2 < length_0 ? _GEN_429 : _GEN_333; // @[executor.scala 290:56]
  wire [7:0] _GEN_526 = 8'h2 < length_0 ? _GEN_430 : _GEN_334; // @[executor.scala 290:56]
  wire [7:0] _GEN_527 = 8'h2 < length_0 ? _GEN_431 : _GEN_335; // @[executor.scala 290:56]
  wire [7:0] _GEN_528 = 8'h2 < length_0 ? _GEN_432 : _GEN_336; // @[executor.scala 290:56]
  wire [7:0] _GEN_529 = 8'h2 < length_0 ? _GEN_433 : _GEN_337; // @[executor.scala 290:56]
  wire [7:0] _GEN_530 = 8'h2 < length_0 ? _GEN_434 : _GEN_338; // @[executor.scala 290:56]
  wire [7:0] _GEN_531 = 8'h2 < length_0 ? _GEN_435 : _GEN_339; // @[executor.scala 290:56]
  wire [7:0] _GEN_532 = 8'h2 < length_0 ? _GEN_436 : _GEN_340; // @[executor.scala 290:56]
  wire [7:0] _GEN_533 = 8'h2 < length_0 ? _GEN_437 : _GEN_341; // @[executor.scala 290:56]
  wire [7:0] _GEN_534 = 8'h2 < length_0 ? _GEN_438 : _GEN_342; // @[executor.scala 290:56]
  wire [7:0] _GEN_535 = 8'h2 < length_0 ? _GEN_439 : _GEN_343; // @[executor.scala 290:56]
  wire [7:0] _GEN_536 = 8'h2 < length_0 ? _GEN_440 : _GEN_344; // @[executor.scala 290:56]
  wire [7:0] _GEN_537 = 8'h2 < length_0 ? _GEN_441 : _GEN_345; // @[executor.scala 290:56]
  wire [7:0] _GEN_538 = 8'h2 < length_0 ? _GEN_442 : _GEN_346; // @[executor.scala 290:56]
  wire [7:0] _GEN_539 = 8'h2 < length_0 ? _GEN_443 : _GEN_347; // @[executor.scala 290:56]
  wire [7:0] _GEN_540 = 8'h2 < length_0 ? _GEN_444 : _GEN_348; // @[executor.scala 290:56]
  wire [7:0] _GEN_541 = 8'h2 < length_0 ? _GEN_445 : _GEN_349; // @[executor.scala 290:56]
  wire [7:0] _GEN_542 = 8'h2 < length_0 ? _GEN_446 : _GEN_350; // @[executor.scala 290:56]
  wire [7:0] _GEN_543 = 8'h2 < length_0 ? _GEN_447 : _GEN_351; // @[executor.scala 290:56]
  wire [7:0] _GEN_544 = 8'h2 < length_0 ? _GEN_448 : _GEN_352; // @[executor.scala 290:56]
  wire [7:0] _GEN_545 = 8'h2 < length_0 ? _GEN_449 : _GEN_353; // @[executor.scala 290:56]
  wire [7:0] _GEN_546 = 8'h2 < length_0 ? _GEN_450 : _GEN_354; // @[executor.scala 290:56]
  wire [7:0] _GEN_547 = 8'h2 < length_0 ? _GEN_451 : _GEN_355; // @[executor.scala 290:56]
  wire [7:0] _GEN_548 = 8'h2 < length_0 ? _GEN_452 : _GEN_356; // @[executor.scala 290:56]
  wire [7:0] _GEN_549 = 8'h2 < length_0 ? _GEN_453 : _GEN_357; // @[executor.scala 290:56]
  wire [7:0] _GEN_550 = 8'h2 < length_0 ? _GEN_454 : _GEN_358; // @[executor.scala 290:56]
  wire [7:0] _GEN_551 = 8'h2 < length_0 ? _GEN_455 : _GEN_359; // @[executor.scala 290:56]
  wire [7:0] _GEN_552 = 8'h2 < length_0 ? _GEN_456 : _GEN_360; // @[executor.scala 290:56]
  wire [7:0] _GEN_553 = 8'h2 < length_0 ? _GEN_457 : _GEN_361; // @[executor.scala 290:56]
  wire [7:0] _GEN_554 = 8'h2 < length_0 ? _GEN_458 : _GEN_362; // @[executor.scala 290:56]
  wire [7:0] _GEN_555 = 8'h2 < length_0 ? _GEN_459 : _GEN_363; // @[executor.scala 290:56]
  wire [7:0] _GEN_556 = 8'h2 < length_0 ? _GEN_460 : _GEN_364; // @[executor.scala 290:56]
  wire [7:0] _GEN_557 = 8'h2 < length_0 ? _GEN_461 : _GEN_365; // @[executor.scala 290:56]
  wire [7:0] _GEN_558 = 8'h2 < length_0 ? _GEN_462 : _GEN_366; // @[executor.scala 290:56]
  wire [7:0] _GEN_559 = 8'h2 < length_0 ? _GEN_463 : _GEN_367; // @[executor.scala 290:56]
  wire [7:0] _GEN_560 = 8'h2 < length_0 ? _GEN_464 : _GEN_368; // @[executor.scala 290:56]
  wire [7:0] _GEN_561 = 8'h2 < length_0 ? _GEN_465 : _GEN_369; // @[executor.scala 290:56]
  wire [7:0] _GEN_562 = 8'h2 < length_0 ? _GEN_466 : _GEN_370; // @[executor.scala 290:56]
  wire [7:0] _GEN_563 = 8'h2 < length_0 ? _GEN_467 : _GEN_371; // @[executor.scala 290:56]
  wire [7:0] _GEN_564 = 8'h2 < length_0 ? _GEN_468 : _GEN_372; // @[executor.scala 290:56]
  wire [7:0] _GEN_565 = 8'h2 < length_0 ? _GEN_469 : _GEN_373; // @[executor.scala 290:56]
  wire [7:0] _GEN_566 = 8'h2 < length_0 ? _GEN_470 : _GEN_374; // @[executor.scala 290:56]
  wire [7:0] _GEN_567 = 8'h2 < length_0 ? _GEN_471 : _GEN_375; // @[executor.scala 290:56]
  wire [7:0] _GEN_568 = 8'h2 < length_0 ? _GEN_472 : _GEN_376; // @[executor.scala 290:56]
  wire [7:0] _GEN_569 = 8'h2 < length_0 ? _GEN_473 : _GEN_377; // @[executor.scala 290:56]
  wire [7:0] _GEN_570 = 8'h2 < length_0 ? _GEN_474 : _GEN_378; // @[executor.scala 290:56]
  wire [7:0] _GEN_571 = 8'h2 < length_0 ? _GEN_475 : _GEN_379; // @[executor.scala 290:56]
  wire [7:0] _GEN_572 = 8'h2 < length_0 ? _GEN_476 : _GEN_380; // @[executor.scala 290:56]
  wire [7:0] _GEN_573 = 8'h2 < length_0 ? _GEN_477 : _GEN_381; // @[executor.scala 290:56]
  wire [7:0] _GEN_574 = 8'h2 < length_0 ? _GEN_478 : _GEN_382; // @[executor.scala 290:56]
  wire [7:0] _GEN_575 = 8'h2 < length_0 ? _GEN_479 : _GEN_383; // @[executor.scala 290:56]
  wire [7:0] field_byte_3 = field_0[39:32]; // @[executor.scala 287:53]
  wire [7:0] total_offset_3 = offset_0 + 8'h3; // @[executor.scala 289:53]
  wire [7:0] _GEN_576 = 7'h0 == total_offset_3[6:0] ? field_byte_3 : _GEN_480; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_577 = 7'h1 == total_offset_3[6:0] ? field_byte_3 : _GEN_481; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_578 = 7'h2 == total_offset_3[6:0] ? field_byte_3 : _GEN_482; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_579 = 7'h3 == total_offset_3[6:0] ? field_byte_3 : _GEN_483; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_580 = 7'h4 == total_offset_3[6:0] ? field_byte_3 : _GEN_484; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_581 = 7'h5 == total_offset_3[6:0] ? field_byte_3 : _GEN_485; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_582 = 7'h6 == total_offset_3[6:0] ? field_byte_3 : _GEN_486; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_583 = 7'h7 == total_offset_3[6:0] ? field_byte_3 : _GEN_487; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_584 = 7'h8 == total_offset_3[6:0] ? field_byte_3 : _GEN_488; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_585 = 7'h9 == total_offset_3[6:0] ? field_byte_3 : _GEN_489; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_586 = 7'ha == total_offset_3[6:0] ? field_byte_3 : _GEN_490; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_587 = 7'hb == total_offset_3[6:0] ? field_byte_3 : _GEN_491; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_588 = 7'hc == total_offset_3[6:0] ? field_byte_3 : _GEN_492; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_589 = 7'hd == total_offset_3[6:0] ? field_byte_3 : _GEN_493; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_590 = 7'he == total_offset_3[6:0] ? field_byte_3 : _GEN_494; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_591 = 7'hf == total_offset_3[6:0] ? field_byte_3 : _GEN_495; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_592 = 7'h10 == total_offset_3[6:0] ? field_byte_3 : _GEN_496; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_593 = 7'h11 == total_offset_3[6:0] ? field_byte_3 : _GEN_497; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_594 = 7'h12 == total_offset_3[6:0] ? field_byte_3 : _GEN_498; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_595 = 7'h13 == total_offset_3[6:0] ? field_byte_3 : _GEN_499; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_596 = 7'h14 == total_offset_3[6:0] ? field_byte_3 : _GEN_500; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_597 = 7'h15 == total_offset_3[6:0] ? field_byte_3 : _GEN_501; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_598 = 7'h16 == total_offset_3[6:0] ? field_byte_3 : _GEN_502; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_599 = 7'h17 == total_offset_3[6:0] ? field_byte_3 : _GEN_503; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_600 = 7'h18 == total_offset_3[6:0] ? field_byte_3 : _GEN_504; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_601 = 7'h19 == total_offset_3[6:0] ? field_byte_3 : _GEN_505; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_602 = 7'h1a == total_offset_3[6:0] ? field_byte_3 : _GEN_506; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_603 = 7'h1b == total_offset_3[6:0] ? field_byte_3 : _GEN_507; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_604 = 7'h1c == total_offset_3[6:0] ? field_byte_3 : _GEN_508; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_605 = 7'h1d == total_offset_3[6:0] ? field_byte_3 : _GEN_509; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_606 = 7'h1e == total_offset_3[6:0] ? field_byte_3 : _GEN_510; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_607 = 7'h1f == total_offset_3[6:0] ? field_byte_3 : _GEN_511; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_608 = 7'h20 == total_offset_3[6:0] ? field_byte_3 : _GEN_512; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_609 = 7'h21 == total_offset_3[6:0] ? field_byte_3 : _GEN_513; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_610 = 7'h22 == total_offset_3[6:0] ? field_byte_3 : _GEN_514; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_611 = 7'h23 == total_offset_3[6:0] ? field_byte_3 : _GEN_515; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_612 = 7'h24 == total_offset_3[6:0] ? field_byte_3 : _GEN_516; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_613 = 7'h25 == total_offset_3[6:0] ? field_byte_3 : _GEN_517; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_614 = 7'h26 == total_offset_3[6:0] ? field_byte_3 : _GEN_518; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_615 = 7'h27 == total_offset_3[6:0] ? field_byte_3 : _GEN_519; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_616 = 7'h28 == total_offset_3[6:0] ? field_byte_3 : _GEN_520; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_617 = 7'h29 == total_offset_3[6:0] ? field_byte_3 : _GEN_521; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_618 = 7'h2a == total_offset_3[6:0] ? field_byte_3 : _GEN_522; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_619 = 7'h2b == total_offset_3[6:0] ? field_byte_3 : _GEN_523; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_620 = 7'h2c == total_offset_3[6:0] ? field_byte_3 : _GEN_524; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_621 = 7'h2d == total_offset_3[6:0] ? field_byte_3 : _GEN_525; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_622 = 7'h2e == total_offset_3[6:0] ? field_byte_3 : _GEN_526; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_623 = 7'h2f == total_offset_3[6:0] ? field_byte_3 : _GEN_527; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_624 = 7'h30 == total_offset_3[6:0] ? field_byte_3 : _GEN_528; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_625 = 7'h31 == total_offset_3[6:0] ? field_byte_3 : _GEN_529; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_626 = 7'h32 == total_offset_3[6:0] ? field_byte_3 : _GEN_530; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_627 = 7'h33 == total_offset_3[6:0] ? field_byte_3 : _GEN_531; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_628 = 7'h34 == total_offset_3[6:0] ? field_byte_3 : _GEN_532; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_629 = 7'h35 == total_offset_3[6:0] ? field_byte_3 : _GEN_533; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_630 = 7'h36 == total_offset_3[6:0] ? field_byte_3 : _GEN_534; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_631 = 7'h37 == total_offset_3[6:0] ? field_byte_3 : _GEN_535; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_632 = 7'h38 == total_offset_3[6:0] ? field_byte_3 : _GEN_536; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_633 = 7'h39 == total_offset_3[6:0] ? field_byte_3 : _GEN_537; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_634 = 7'h3a == total_offset_3[6:0] ? field_byte_3 : _GEN_538; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_635 = 7'h3b == total_offset_3[6:0] ? field_byte_3 : _GEN_539; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_636 = 7'h3c == total_offset_3[6:0] ? field_byte_3 : _GEN_540; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_637 = 7'h3d == total_offset_3[6:0] ? field_byte_3 : _GEN_541; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_638 = 7'h3e == total_offset_3[6:0] ? field_byte_3 : _GEN_542; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_639 = 7'h3f == total_offset_3[6:0] ? field_byte_3 : _GEN_543; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_640 = 7'h40 == total_offset_3[6:0] ? field_byte_3 : _GEN_544; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_641 = 7'h41 == total_offset_3[6:0] ? field_byte_3 : _GEN_545; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_642 = 7'h42 == total_offset_3[6:0] ? field_byte_3 : _GEN_546; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_643 = 7'h43 == total_offset_3[6:0] ? field_byte_3 : _GEN_547; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_644 = 7'h44 == total_offset_3[6:0] ? field_byte_3 : _GEN_548; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_645 = 7'h45 == total_offset_3[6:0] ? field_byte_3 : _GEN_549; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_646 = 7'h46 == total_offset_3[6:0] ? field_byte_3 : _GEN_550; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_647 = 7'h47 == total_offset_3[6:0] ? field_byte_3 : _GEN_551; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_648 = 7'h48 == total_offset_3[6:0] ? field_byte_3 : _GEN_552; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_649 = 7'h49 == total_offset_3[6:0] ? field_byte_3 : _GEN_553; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_650 = 7'h4a == total_offset_3[6:0] ? field_byte_3 : _GEN_554; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_651 = 7'h4b == total_offset_3[6:0] ? field_byte_3 : _GEN_555; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_652 = 7'h4c == total_offset_3[6:0] ? field_byte_3 : _GEN_556; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_653 = 7'h4d == total_offset_3[6:0] ? field_byte_3 : _GEN_557; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_654 = 7'h4e == total_offset_3[6:0] ? field_byte_3 : _GEN_558; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_655 = 7'h4f == total_offset_3[6:0] ? field_byte_3 : _GEN_559; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_656 = 7'h50 == total_offset_3[6:0] ? field_byte_3 : _GEN_560; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_657 = 7'h51 == total_offset_3[6:0] ? field_byte_3 : _GEN_561; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_658 = 7'h52 == total_offset_3[6:0] ? field_byte_3 : _GEN_562; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_659 = 7'h53 == total_offset_3[6:0] ? field_byte_3 : _GEN_563; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_660 = 7'h54 == total_offset_3[6:0] ? field_byte_3 : _GEN_564; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_661 = 7'h55 == total_offset_3[6:0] ? field_byte_3 : _GEN_565; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_662 = 7'h56 == total_offset_3[6:0] ? field_byte_3 : _GEN_566; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_663 = 7'h57 == total_offset_3[6:0] ? field_byte_3 : _GEN_567; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_664 = 7'h58 == total_offset_3[6:0] ? field_byte_3 : _GEN_568; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_665 = 7'h59 == total_offset_3[6:0] ? field_byte_3 : _GEN_569; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_666 = 7'h5a == total_offset_3[6:0] ? field_byte_3 : _GEN_570; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_667 = 7'h5b == total_offset_3[6:0] ? field_byte_3 : _GEN_571; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_668 = 7'h5c == total_offset_3[6:0] ? field_byte_3 : _GEN_572; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_669 = 7'h5d == total_offset_3[6:0] ? field_byte_3 : _GEN_573; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_670 = 7'h5e == total_offset_3[6:0] ? field_byte_3 : _GEN_574; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_671 = 7'h5f == total_offset_3[6:0] ? field_byte_3 : _GEN_575; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_672 = 8'h3 < length_0 ? _GEN_576 : _GEN_480; // @[executor.scala 290:56]
  wire [7:0] _GEN_673 = 8'h3 < length_0 ? _GEN_577 : _GEN_481; // @[executor.scala 290:56]
  wire [7:0] _GEN_674 = 8'h3 < length_0 ? _GEN_578 : _GEN_482; // @[executor.scala 290:56]
  wire [7:0] _GEN_675 = 8'h3 < length_0 ? _GEN_579 : _GEN_483; // @[executor.scala 290:56]
  wire [7:0] _GEN_676 = 8'h3 < length_0 ? _GEN_580 : _GEN_484; // @[executor.scala 290:56]
  wire [7:0] _GEN_677 = 8'h3 < length_0 ? _GEN_581 : _GEN_485; // @[executor.scala 290:56]
  wire [7:0] _GEN_678 = 8'h3 < length_0 ? _GEN_582 : _GEN_486; // @[executor.scala 290:56]
  wire [7:0] _GEN_679 = 8'h3 < length_0 ? _GEN_583 : _GEN_487; // @[executor.scala 290:56]
  wire [7:0] _GEN_680 = 8'h3 < length_0 ? _GEN_584 : _GEN_488; // @[executor.scala 290:56]
  wire [7:0] _GEN_681 = 8'h3 < length_0 ? _GEN_585 : _GEN_489; // @[executor.scala 290:56]
  wire [7:0] _GEN_682 = 8'h3 < length_0 ? _GEN_586 : _GEN_490; // @[executor.scala 290:56]
  wire [7:0] _GEN_683 = 8'h3 < length_0 ? _GEN_587 : _GEN_491; // @[executor.scala 290:56]
  wire [7:0] _GEN_684 = 8'h3 < length_0 ? _GEN_588 : _GEN_492; // @[executor.scala 290:56]
  wire [7:0] _GEN_685 = 8'h3 < length_0 ? _GEN_589 : _GEN_493; // @[executor.scala 290:56]
  wire [7:0] _GEN_686 = 8'h3 < length_0 ? _GEN_590 : _GEN_494; // @[executor.scala 290:56]
  wire [7:0] _GEN_687 = 8'h3 < length_0 ? _GEN_591 : _GEN_495; // @[executor.scala 290:56]
  wire [7:0] _GEN_688 = 8'h3 < length_0 ? _GEN_592 : _GEN_496; // @[executor.scala 290:56]
  wire [7:0] _GEN_689 = 8'h3 < length_0 ? _GEN_593 : _GEN_497; // @[executor.scala 290:56]
  wire [7:0] _GEN_690 = 8'h3 < length_0 ? _GEN_594 : _GEN_498; // @[executor.scala 290:56]
  wire [7:0] _GEN_691 = 8'h3 < length_0 ? _GEN_595 : _GEN_499; // @[executor.scala 290:56]
  wire [7:0] _GEN_692 = 8'h3 < length_0 ? _GEN_596 : _GEN_500; // @[executor.scala 290:56]
  wire [7:0] _GEN_693 = 8'h3 < length_0 ? _GEN_597 : _GEN_501; // @[executor.scala 290:56]
  wire [7:0] _GEN_694 = 8'h3 < length_0 ? _GEN_598 : _GEN_502; // @[executor.scala 290:56]
  wire [7:0] _GEN_695 = 8'h3 < length_0 ? _GEN_599 : _GEN_503; // @[executor.scala 290:56]
  wire [7:0] _GEN_696 = 8'h3 < length_0 ? _GEN_600 : _GEN_504; // @[executor.scala 290:56]
  wire [7:0] _GEN_697 = 8'h3 < length_0 ? _GEN_601 : _GEN_505; // @[executor.scala 290:56]
  wire [7:0] _GEN_698 = 8'h3 < length_0 ? _GEN_602 : _GEN_506; // @[executor.scala 290:56]
  wire [7:0] _GEN_699 = 8'h3 < length_0 ? _GEN_603 : _GEN_507; // @[executor.scala 290:56]
  wire [7:0] _GEN_700 = 8'h3 < length_0 ? _GEN_604 : _GEN_508; // @[executor.scala 290:56]
  wire [7:0] _GEN_701 = 8'h3 < length_0 ? _GEN_605 : _GEN_509; // @[executor.scala 290:56]
  wire [7:0] _GEN_702 = 8'h3 < length_0 ? _GEN_606 : _GEN_510; // @[executor.scala 290:56]
  wire [7:0] _GEN_703 = 8'h3 < length_0 ? _GEN_607 : _GEN_511; // @[executor.scala 290:56]
  wire [7:0] _GEN_704 = 8'h3 < length_0 ? _GEN_608 : _GEN_512; // @[executor.scala 290:56]
  wire [7:0] _GEN_705 = 8'h3 < length_0 ? _GEN_609 : _GEN_513; // @[executor.scala 290:56]
  wire [7:0] _GEN_706 = 8'h3 < length_0 ? _GEN_610 : _GEN_514; // @[executor.scala 290:56]
  wire [7:0] _GEN_707 = 8'h3 < length_0 ? _GEN_611 : _GEN_515; // @[executor.scala 290:56]
  wire [7:0] _GEN_708 = 8'h3 < length_0 ? _GEN_612 : _GEN_516; // @[executor.scala 290:56]
  wire [7:0] _GEN_709 = 8'h3 < length_0 ? _GEN_613 : _GEN_517; // @[executor.scala 290:56]
  wire [7:0] _GEN_710 = 8'h3 < length_0 ? _GEN_614 : _GEN_518; // @[executor.scala 290:56]
  wire [7:0] _GEN_711 = 8'h3 < length_0 ? _GEN_615 : _GEN_519; // @[executor.scala 290:56]
  wire [7:0] _GEN_712 = 8'h3 < length_0 ? _GEN_616 : _GEN_520; // @[executor.scala 290:56]
  wire [7:0] _GEN_713 = 8'h3 < length_0 ? _GEN_617 : _GEN_521; // @[executor.scala 290:56]
  wire [7:0] _GEN_714 = 8'h3 < length_0 ? _GEN_618 : _GEN_522; // @[executor.scala 290:56]
  wire [7:0] _GEN_715 = 8'h3 < length_0 ? _GEN_619 : _GEN_523; // @[executor.scala 290:56]
  wire [7:0] _GEN_716 = 8'h3 < length_0 ? _GEN_620 : _GEN_524; // @[executor.scala 290:56]
  wire [7:0] _GEN_717 = 8'h3 < length_0 ? _GEN_621 : _GEN_525; // @[executor.scala 290:56]
  wire [7:0] _GEN_718 = 8'h3 < length_0 ? _GEN_622 : _GEN_526; // @[executor.scala 290:56]
  wire [7:0] _GEN_719 = 8'h3 < length_0 ? _GEN_623 : _GEN_527; // @[executor.scala 290:56]
  wire [7:0] _GEN_720 = 8'h3 < length_0 ? _GEN_624 : _GEN_528; // @[executor.scala 290:56]
  wire [7:0] _GEN_721 = 8'h3 < length_0 ? _GEN_625 : _GEN_529; // @[executor.scala 290:56]
  wire [7:0] _GEN_722 = 8'h3 < length_0 ? _GEN_626 : _GEN_530; // @[executor.scala 290:56]
  wire [7:0] _GEN_723 = 8'h3 < length_0 ? _GEN_627 : _GEN_531; // @[executor.scala 290:56]
  wire [7:0] _GEN_724 = 8'h3 < length_0 ? _GEN_628 : _GEN_532; // @[executor.scala 290:56]
  wire [7:0] _GEN_725 = 8'h3 < length_0 ? _GEN_629 : _GEN_533; // @[executor.scala 290:56]
  wire [7:0] _GEN_726 = 8'h3 < length_0 ? _GEN_630 : _GEN_534; // @[executor.scala 290:56]
  wire [7:0] _GEN_727 = 8'h3 < length_0 ? _GEN_631 : _GEN_535; // @[executor.scala 290:56]
  wire [7:0] _GEN_728 = 8'h3 < length_0 ? _GEN_632 : _GEN_536; // @[executor.scala 290:56]
  wire [7:0] _GEN_729 = 8'h3 < length_0 ? _GEN_633 : _GEN_537; // @[executor.scala 290:56]
  wire [7:0] _GEN_730 = 8'h3 < length_0 ? _GEN_634 : _GEN_538; // @[executor.scala 290:56]
  wire [7:0] _GEN_731 = 8'h3 < length_0 ? _GEN_635 : _GEN_539; // @[executor.scala 290:56]
  wire [7:0] _GEN_732 = 8'h3 < length_0 ? _GEN_636 : _GEN_540; // @[executor.scala 290:56]
  wire [7:0] _GEN_733 = 8'h3 < length_0 ? _GEN_637 : _GEN_541; // @[executor.scala 290:56]
  wire [7:0] _GEN_734 = 8'h3 < length_0 ? _GEN_638 : _GEN_542; // @[executor.scala 290:56]
  wire [7:0] _GEN_735 = 8'h3 < length_0 ? _GEN_639 : _GEN_543; // @[executor.scala 290:56]
  wire [7:0] _GEN_736 = 8'h3 < length_0 ? _GEN_640 : _GEN_544; // @[executor.scala 290:56]
  wire [7:0] _GEN_737 = 8'h3 < length_0 ? _GEN_641 : _GEN_545; // @[executor.scala 290:56]
  wire [7:0] _GEN_738 = 8'h3 < length_0 ? _GEN_642 : _GEN_546; // @[executor.scala 290:56]
  wire [7:0] _GEN_739 = 8'h3 < length_0 ? _GEN_643 : _GEN_547; // @[executor.scala 290:56]
  wire [7:0] _GEN_740 = 8'h3 < length_0 ? _GEN_644 : _GEN_548; // @[executor.scala 290:56]
  wire [7:0] _GEN_741 = 8'h3 < length_0 ? _GEN_645 : _GEN_549; // @[executor.scala 290:56]
  wire [7:0] _GEN_742 = 8'h3 < length_0 ? _GEN_646 : _GEN_550; // @[executor.scala 290:56]
  wire [7:0] _GEN_743 = 8'h3 < length_0 ? _GEN_647 : _GEN_551; // @[executor.scala 290:56]
  wire [7:0] _GEN_744 = 8'h3 < length_0 ? _GEN_648 : _GEN_552; // @[executor.scala 290:56]
  wire [7:0] _GEN_745 = 8'h3 < length_0 ? _GEN_649 : _GEN_553; // @[executor.scala 290:56]
  wire [7:0] _GEN_746 = 8'h3 < length_0 ? _GEN_650 : _GEN_554; // @[executor.scala 290:56]
  wire [7:0] _GEN_747 = 8'h3 < length_0 ? _GEN_651 : _GEN_555; // @[executor.scala 290:56]
  wire [7:0] _GEN_748 = 8'h3 < length_0 ? _GEN_652 : _GEN_556; // @[executor.scala 290:56]
  wire [7:0] _GEN_749 = 8'h3 < length_0 ? _GEN_653 : _GEN_557; // @[executor.scala 290:56]
  wire [7:0] _GEN_750 = 8'h3 < length_0 ? _GEN_654 : _GEN_558; // @[executor.scala 290:56]
  wire [7:0] _GEN_751 = 8'h3 < length_0 ? _GEN_655 : _GEN_559; // @[executor.scala 290:56]
  wire [7:0] _GEN_752 = 8'h3 < length_0 ? _GEN_656 : _GEN_560; // @[executor.scala 290:56]
  wire [7:0] _GEN_753 = 8'h3 < length_0 ? _GEN_657 : _GEN_561; // @[executor.scala 290:56]
  wire [7:0] _GEN_754 = 8'h3 < length_0 ? _GEN_658 : _GEN_562; // @[executor.scala 290:56]
  wire [7:0] _GEN_755 = 8'h3 < length_0 ? _GEN_659 : _GEN_563; // @[executor.scala 290:56]
  wire [7:0] _GEN_756 = 8'h3 < length_0 ? _GEN_660 : _GEN_564; // @[executor.scala 290:56]
  wire [7:0] _GEN_757 = 8'h3 < length_0 ? _GEN_661 : _GEN_565; // @[executor.scala 290:56]
  wire [7:0] _GEN_758 = 8'h3 < length_0 ? _GEN_662 : _GEN_566; // @[executor.scala 290:56]
  wire [7:0] _GEN_759 = 8'h3 < length_0 ? _GEN_663 : _GEN_567; // @[executor.scala 290:56]
  wire [7:0] _GEN_760 = 8'h3 < length_0 ? _GEN_664 : _GEN_568; // @[executor.scala 290:56]
  wire [7:0] _GEN_761 = 8'h3 < length_0 ? _GEN_665 : _GEN_569; // @[executor.scala 290:56]
  wire [7:0] _GEN_762 = 8'h3 < length_0 ? _GEN_666 : _GEN_570; // @[executor.scala 290:56]
  wire [7:0] _GEN_763 = 8'h3 < length_0 ? _GEN_667 : _GEN_571; // @[executor.scala 290:56]
  wire [7:0] _GEN_764 = 8'h3 < length_0 ? _GEN_668 : _GEN_572; // @[executor.scala 290:56]
  wire [7:0] _GEN_765 = 8'h3 < length_0 ? _GEN_669 : _GEN_573; // @[executor.scala 290:56]
  wire [7:0] _GEN_766 = 8'h3 < length_0 ? _GEN_670 : _GEN_574; // @[executor.scala 290:56]
  wire [7:0] _GEN_767 = 8'h3 < length_0 ? _GEN_671 : _GEN_575; // @[executor.scala 290:56]
  wire [7:0] field_byte_4 = field_0[31:24]; // @[executor.scala 287:53]
  wire [7:0] total_offset_4 = offset_0 + 8'h4; // @[executor.scala 289:53]
  wire [7:0] _GEN_768 = 7'h0 == total_offset_4[6:0] ? field_byte_4 : _GEN_672; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_769 = 7'h1 == total_offset_4[6:0] ? field_byte_4 : _GEN_673; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_770 = 7'h2 == total_offset_4[6:0] ? field_byte_4 : _GEN_674; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_771 = 7'h3 == total_offset_4[6:0] ? field_byte_4 : _GEN_675; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_772 = 7'h4 == total_offset_4[6:0] ? field_byte_4 : _GEN_676; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_773 = 7'h5 == total_offset_4[6:0] ? field_byte_4 : _GEN_677; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_774 = 7'h6 == total_offset_4[6:0] ? field_byte_4 : _GEN_678; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_775 = 7'h7 == total_offset_4[6:0] ? field_byte_4 : _GEN_679; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_776 = 7'h8 == total_offset_4[6:0] ? field_byte_4 : _GEN_680; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_777 = 7'h9 == total_offset_4[6:0] ? field_byte_4 : _GEN_681; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_778 = 7'ha == total_offset_4[6:0] ? field_byte_4 : _GEN_682; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_779 = 7'hb == total_offset_4[6:0] ? field_byte_4 : _GEN_683; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_780 = 7'hc == total_offset_4[6:0] ? field_byte_4 : _GEN_684; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_781 = 7'hd == total_offset_4[6:0] ? field_byte_4 : _GEN_685; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_782 = 7'he == total_offset_4[6:0] ? field_byte_4 : _GEN_686; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_783 = 7'hf == total_offset_4[6:0] ? field_byte_4 : _GEN_687; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_784 = 7'h10 == total_offset_4[6:0] ? field_byte_4 : _GEN_688; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_785 = 7'h11 == total_offset_4[6:0] ? field_byte_4 : _GEN_689; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_786 = 7'h12 == total_offset_4[6:0] ? field_byte_4 : _GEN_690; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_787 = 7'h13 == total_offset_4[6:0] ? field_byte_4 : _GEN_691; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_788 = 7'h14 == total_offset_4[6:0] ? field_byte_4 : _GEN_692; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_789 = 7'h15 == total_offset_4[6:0] ? field_byte_4 : _GEN_693; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_790 = 7'h16 == total_offset_4[6:0] ? field_byte_4 : _GEN_694; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_791 = 7'h17 == total_offset_4[6:0] ? field_byte_4 : _GEN_695; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_792 = 7'h18 == total_offset_4[6:0] ? field_byte_4 : _GEN_696; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_793 = 7'h19 == total_offset_4[6:0] ? field_byte_4 : _GEN_697; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_794 = 7'h1a == total_offset_4[6:0] ? field_byte_4 : _GEN_698; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_795 = 7'h1b == total_offset_4[6:0] ? field_byte_4 : _GEN_699; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_796 = 7'h1c == total_offset_4[6:0] ? field_byte_4 : _GEN_700; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_797 = 7'h1d == total_offset_4[6:0] ? field_byte_4 : _GEN_701; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_798 = 7'h1e == total_offset_4[6:0] ? field_byte_4 : _GEN_702; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_799 = 7'h1f == total_offset_4[6:0] ? field_byte_4 : _GEN_703; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_800 = 7'h20 == total_offset_4[6:0] ? field_byte_4 : _GEN_704; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_801 = 7'h21 == total_offset_4[6:0] ? field_byte_4 : _GEN_705; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_802 = 7'h22 == total_offset_4[6:0] ? field_byte_4 : _GEN_706; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_803 = 7'h23 == total_offset_4[6:0] ? field_byte_4 : _GEN_707; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_804 = 7'h24 == total_offset_4[6:0] ? field_byte_4 : _GEN_708; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_805 = 7'h25 == total_offset_4[6:0] ? field_byte_4 : _GEN_709; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_806 = 7'h26 == total_offset_4[6:0] ? field_byte_4 : _GEN_710; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_807 = 7'h27 == total_offset_4[6:0] ? field_byte_4 : _GEN_711; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_808 = 7'h28 == total_offset_4[6:0] ? field_byte_4 : _GEN_712; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_809 = 7'h29 == total_offset_4[6:0] ? field_byte_4 : _GEN_713; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_810 = 7'h2a == total_offset_4[6:0] ? field_byte_4 : _GEN_714; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_811 = 7'h2b == total_offset_4[6:0] ? field_byte_4 : _GEN_715; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_812 = 7'h2c == total_offset_4[6:0] ? field_byte_4 : _GEN_716; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_813 = 7'h2d == total_offset_4[6:0] ? field_byte_4 : _GEN_717; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_814 = 7'h2e == total_offset_4[6:0] ? field_byte_4 : _GEN_718; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_815 = 7'h2f == total_offset_4[6:0] ? field_byte_4 : _GEN_719; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_816 = 7'h30 == total_offset_4[6:0] ? field_byte_4 : _GEN_720; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_817 = 7'h31 == total_offset_4[6:0] ? field_byte_4 : _GEN_721; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_818 = 7'h32 == total_offset_4[6:0] ? field_byte_4 : _GEN_722; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_819 = 7'h33 == total_offset_4[6:0] ? field_byte_4 : _GEN_723; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_820 = 7'h34 == total_offset_4[6:0] ? field_byte_4 : _GEN_724; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_821 = 7'h35 == total_offset_4[6:0] ? field_byte_4 : _GEN_725; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_822 = 7'h36 == total_offset_4[6:0] ? field_byte_4 : _GEN_726; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_823 = 7'h37 == total_offset_4[6:0] ? field_byte_4 : _GEN_727; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_824 = 7'h38 == total_offset_4[6:0] ? field_byte_4 : _GEN_728; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_825 = 7'h39 == total_offset_4[6:0] ? field_byte_4 : _GEN_729; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_826 = 7'h3a == total_offset_4[6:0] ? field_byte_4 : _GEN_730; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_827 = 7'h3b == total_offset_4[6:0] ? field_byte_4 : _GEN_731; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_828 = 7'h3c == total_offset_4[6:0] ? field_byte_4 : _GEN_732; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_829 = 7'h3d == total_offset_4[6:0] ? field_byte_4 : _GEN_733; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_830 = 7'h3e == total_offset_4[6:0] ? field_byte_4 : _GEN_734; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_831 = 7'h3f == total_offset_4[6:0] ? field_byte_4 : _GEN_735; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_832 = 7'h40 == total_offset_4[6:0] ? field_byte_4 : _GEN_736; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_833 = 7'h41 == total_offset_4[6:0] ? field_byte_4 : _GEN_737; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_834 = 7'h42 == total_offset_4[6:0] ? field_byte_4 : _GEN_738; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_835 = 7'h43 == total_offset_4[6:0] ? field_byte_4 : _GEN_739; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_836 = 7'h44 == total_offset_4[6:0] ? field_byte_4 : _GEN_740; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_837 = 7'h45 == total_offset_4[6:0] ? field_byte_4 : _GEN_741; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_838 = 7'h46 == total_offset_4[6:0] ? field_byte_4 : _GEN_742; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_839 = 7'h47 == total_offset_4[6:0] ? field_byte_4 : _GEN_743; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_840 = 7'h48 == total_offset_4[6:0] ? field_byte_4 : _GEN_744; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_841 = 7'h49 == total_offset_4[6:0] ? field_byte_4 : _GEN_745; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_842 = 7'h4a == total_offset_4[6:0] ? field_byte_4 : _GEN_746; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_843 = 7'h4b == total_offset_4[6:0] ? field_byte_4 : _GEN_747; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_844 = 7'h4c == total_offset_4[6:0] ? field_byte_4 : _GEN_748; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_845 = 7'h4d == total_offset_4[6:0] ? field_byte_4 : _GEN_749; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_846 = 7'h4e == total_offset_4[6:0] ? field_byte_4 : _GEN_750; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_847 = 7'h4f == total_offset_4[6:0] ? field_byte_4 : _GEN_751; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_848 = 7'h50 == total_offset_4[6:0] ? field_byte_4 : _GEN_752; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_849 = 7'h51 == total_offset_4[6:0] ? field_byte_4 : _GEN_753; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_850 = 7'h52 == total_offset_4[6:0] ? field_byte_4 : _GEN_754; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_851 = 7'h53 == total_offset_4[6:0] ? field_byte_4 : _GEN_755; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_852 = 7'h54 == total_offset_4[6:0] ? field_byte_4 : _GEN_756; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_853 = 7'h55 == total_offset_4[6:0] ? field_byte_4 : _GEN_757; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_854 = 7'h56 == total_offset_4[6:0] ? field_byte_4 : _GEN_758; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_855 = 7'h57 == total_offset_4[6:0] ? field_byte_4 : _GEN_759; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_856 = 7'h58 == total_offset_4[6:0] ? field_byte_4 : _GEN_760; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_857 = 7'h59 == total_offset_4[6:0] ? field_byte_4 : _GEN_761; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_858 = 7'h5a == total_offset_4[6:0] ? field_byte_4 : _GEN_762; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_859 = 7'h5b == total_offset_4[6:0] ? field_byte_4 : _GEN_763; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_860 = 7'h5c == total_offset_4[6:0] ? field_byte_4 : _GEN_764; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_861 = 7'h5d == total_offset_4[6:0] ? field_byte_4 : _GEN_765; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_862 = 7'h5e == total_offset_4[6:0] ? field_byte_4 : _GEN_766; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_863 = 7'h5f == total_offset_4[6:0] ? field_byte_4 : _GEN_767; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_864 = 8'h4 < length_0 ? _GEN_768 : _GEN_672; // @[executor.scala 290:56]
  wire [7:0] _GEN_865 = 8'h4 < length_0 ? _GEN_769 : _GEN_673; // @[executor.scala 290:56]
  wire [7:0] _GEN_866 = 8'h4 < length_0 ? _GEN_770 : _GEN_674; // @[executor.scala 290:56]
  wire [7:0] _GEN_867 = 8'h4 < length_0 ? _GEN_771 : _GEN_675; // @[executor.scala 290:56]
  wire [7:0] _GEN_868 = 8'h4 < length_0 ? _GEN_772 : _GEN_676; // @[executor.scala 290:56]
  wire [7:0] _GEN_869 = 8'h4 < length_0 ? _GEN_773 : _GEN_677; // @[executor.scala 290:56]
  wire [7:0] _GEN_870 = 8'h4 < length_0 ? _GEN_774 : _GEN_678; // @[executor.scala 290:56]
  wire [7:0] _GEN_871 = 8'h4 < length_0 ? _GEN_775 : _GEN_679; // @[executor.scala 290:56]
  wire [7:0] _GEN_872 = 8'h4 < length_0 ? _GEN_776 : _GEN_680; // @[executor.scala 290:56]
  wire [7:0] _GEN_873 = 8'h4 < length_0 ? _GEN_777 : _GEN_681; // @[executor.scala 290:56]
  wire [7:0] _GEN_874 = 8'h4 < length_0 ? _GEN_778 : _GEN_682; // @[executor.scala 290:56]
  wire [7:0] _GEN_875 = 8'h4 < length_0 ? _GEN_779 : _GEN_683; // @[executor.scala 290:56]
  wire [7:0] _GEN_876 = 8'h4 < length_0 ? _GEN_780 : _GEN_684; // @[executor.scala 290:56]
  wire [7:0] _GEN_877 = 8'h4 < length_0 ? _GEN_781 : _GEN_685; // @[executor.scala 290:56]
  wire [7:0] _GEN_878 = 8'h4 < length_0 ? _GEN_782 : _GEN_686; // @[executor.scala 290:56]
  wire [7:0] _GEN_879 = 8'h4 < length_0 ? _GEN_783 : _GEN_687; // @[executor.scala 290:56]
  wire [7:0] _GEN_880 = 8'h4 < length_0 ? _GEN_784 : _GEN_688; // @[executor.scala 290:56]
  wire [7:0] _GEN_881 = 8'h4 < length_0 ? _GEN_785 : _GEN_689; // @[executor.scala 290:56]
  wire [7:0] _GEN_882 = 8'h4 < length_0 ? _GEN_786 : _GEN_690; // @[executor.scala 290:56]
  wire [7:0] _GEN_883 = 8'h4 < length_0 ? _GEN_787 : _GEN_691; // @[executor.scala 290:56]
  wire [7:0] _GEN_884 = 8'h4 < length_0 ? _GEN_788 : _GEN_692; // @[executor.scala 290:56]
  wire [7:0] _GEN_885 = 8'h4 < length_0 ? _GEN_789 : _GEN_693; // @[executor.scala 290:56]
  wire [7:0] _GEN_886 = 8'h4 < length_0 ? _GEN_790 : _GEN_694; // @[executor.scala 290:56]
  wire [7:0] _GEN_887 = 8'h4 < length_0 ? _GEN_791 : _GEN_695; // @[executor.scala 290:56]
  wire [7:0] _GEN_888 = 8'h4 < length_0 ? _GEN_792 : _GEN_696; // @[executor.scala 290:56]
  wire [7:0] _GEN_889 = 8'h4 < length_0 ? _GEN_793 : _GEN_697; // @[executor.scala 290:56]
  wire [7:0] _GEN_890 = 8'h4 < length_0 ? _GEN_794 : _GEN_698; // @[executor.scala 290:56]
  wire [7:0] _GEN_891 = 8'h4 < length_0 ? _GEN_795 : _GEN_699; // @[executor.scala 290:56]
  wire [7:0] _GEN_892 = 8'h4 < length_0 ? _GEN_796 : _GEN_700; // @[executor.scala 290:56]
  wire [7:0] _GEN_893 = 8'h4 < length_0 ? _GEN_797 : _GEN_701; // @[executor.scala 290:56]
  wire [7:0] _GEN_894 = 8'h4 < length_0 ? _GEN_798 : _GEN_702; // @[executor.scala 290:56]
  wire [7:0] _GEN_895 = 8'h4 < length_0 ? _GEN_799 : _GEN_703; // @[executor.scala 290:56]
  wire [7:0] _GEN_896 = 8'h4 < length_0 ? _GEN_800 : _GEN_704; // @[executor.scala 290:56]
  wire [7:0] _GEN_897 = 8'h4 < length_0 ? _GEN_801 : _GEN_705; // @[executor.scala 290:56]
  wire [7:0] _GEN_898 = 8'h4 < length_0 ? _GEN_802 : _GEN_706; // @[executor.scala 290:56]
  wire [7:0] _GEN_899 = 8'h4 < length_0 ? _GEN_803 : _GEN_707; // @[executor.scala 290:56]
  wire [7:0] _GEN_900 = 8'h4 < length_0 ? _GEN_804 : _GEN_708; // @[executor.scala 290:56]
  wire [7:0] _GEN_901 = 8'h4 < length_0 ? _GEN_805 : _GEN_709; // @[executor.scala 290:56]
  wire [7:0] _GEN_902 = 8'h4 < length_0 ? _GEN_806 : _GEN_710; // @[executor.scala 290:56]
  wire [7:0] _GEN_903 = 8'h4 < length_0 ? _GEN_807 : _GEN_711; // @[executor.scala 290:56]
  wire [7:0] _GEN_904 = 8'h4 < length_0 ? _GEN_808 : _GEN_712; // @[executor.scala 290:56]
  wire [7:0] _GEN_905 = 8'h4 < length_0 ? _GEN_809 : _GEN_713; // @[executor.scala 290:56]
  wire [7:0] _GEN_906 = 8'h4 < length_0 ? _GEN_810 : _GEN_714; // @[executor.scala 290:56]
  wire [7:0] _GEN_907 = 8'h4 < length_0 ? _GEN_811 : _GEN_715; // @[executor.scala 290:56]
  wire [7:0] _GEN_908 = 8'h4 < length_0 ? _GEN_812 : _GEN_716; // @[executor.scala 290:56]
  wire [7:0] _GEN_909 = 8'h4 < length_0 ? _GEN_813 : _GEN_717; // @[executor.scala 290:56]
  wire [7:0] _GEN_910 = 8'h4 < length_0 ? _GEN_814 : _GEN_718; // @[executor.scala 290:56]
  wire [7:0] _GEN_911 = 8'h4 < length_0 ? _GEN_815 : _GEN_719; // @[executor.scala 290:56]
  wire [7:0] _GEN_912 = 8'h4 < length_0 ? _GEN_816 : _GEN_720; // @[executor.scala 290:56]
  wire [7:0] _GEN_913 = 8'h4 < length_0 ? _GEN_817 : _GEN_721; // @[executor.scala 290:56]
  wire [7:0] _GEN_914 = 8'h4 < length_0 ? _GEN_818 : _GEN_722; // @[executor.scala 290:56]
  wire [7:0] _GEN_915 = 8'h4 < length_0 ? _GEN_819 : _GEN_723; // @[executor.scala 290:56]
  wire [7:0] _GEN_916 = 8'h4 < length_0 ? _GEN_820 : _GEN_724; // @[executor.scala 290:56]
  wire [7:0] _GEN_917 = 8'h4 < length_0 ? _GEN_821 : _GEN_725; // @[executor.scala 290:56]
  wire [7:0] _GEN_918 = 8'h4 < length_0 ? _GEN_822 : _GEN_726; // @[executor.scala 290:56]
  wire [7:0] _GEN_919 = 8'h4 < length_0 ? _GEN_823 : _GEN_727; // @[executor.scala 290:56]
  wire [7:0] _GEN_920 = 8'h4 < length_0 ? _GEN_824 : _GEN_728; // @[executor.scala 290:56]
  wire [7:0] _GEN_921 = 8'h4 < length_0 ? _GEN_825 : _GEN_729; // @[executor.scala 290:56]
  wire [7:0] _GEN_922 = 8'h4 < length_0 ? _GEN_826 : _GEN_730; // @[executor.scala 290:56]
  wire [7:0] _GEN_923 = 8'h4 < length_0 ? _GEN_827 : _GEN_731; // @[executor.scala 290:56]
  wire [7:0] _GEN_924 = 8'h4 < length_0 ? _GEN_828 : _GEN_732; // @[executor.scala 290:56]
  wire [7:0] _GEN_925 = 8'h4 < length_0 ? _GEN_829 : _GEN_733; // @[executor.scala 290:56]
  wire [7:0] _GEN_926 = 8'h4 < length_0 ? _GEN_830 : _GEN_734; // @[executor.scala 290:56]
  wire [7:0] _GEN_927 = 8'h4 < length_0 ? _GEN_831 : _GEN_735; // @[executor.scala 290:56]
  wire [7:0] _GEN_928 = 8'h4 < length_0 ? _GEN_832 : _GEN_736; // @[executor.scala 290:56]
  wire [7:0] _GEN_929 = 8'h4 < length_0 ? _GEN_833 : _GEN_737; // @[executor.scala 290:56]
  wire [7:0] _GEN_930 = 8'h4 < length_0 ? _GEN_834 : _GEN_738; // @[executor.scala 290:56]
  wire [7:0] _GEN_931 = 8'h4 < length_0 ? _GEN_835 : _GEN_739; // @[executor.scala 290:56]
  wire [7:0] _GEN_932 = 8'h4 < length_0 ? _GEN_836 : _GEN_740; // @[executor.scala 290:56]
  wire [7:0] _GEN_933 = 8'h4 < length_0 ? _GEN_837 : _GEN_741; // @[executor.scala 290:56]
  wire [7:0] _GEN_934 = 8'h4 < length_0 ? _GEN_838 : _GEN_742; // @[executor.scala 290:56]
  wire [7:0] _GEN_935 = 8'h4 < length_0 ? _GEN_839 : _GEN_743; // @[executor.scala 290:56]
  wire [7:0] _GEN_936 = 8'h4 < length_0 ? _GEN_840 : _GEN_744; // @[executor.scala 290:56]
  wire [7:0] _GEN_937 = 8'h4 < length_0 ? _GEN_841 : _GEN_745; // @[executor.scala 290:56]
  wire [7:0] _GEN_938 = 8'h4 < length_0 ? _GEN_842 : _GEN_746; // @[executor.scala 290:56]
  wire [7:0] _GEN_939 = 8'h4 < length_0 ? _GEN_843 : _GEN_747; // @[executor.scala 290:56]
  wire [7:0] _GEN_940 = 8'h4 < length_0 ? _GEN_844 : _GEN_748; // @[executor.scala 290:56]
  wire [7:0] _GEN_941 = 8'h4 < length_0 ? _GEN_845 : _GEN_749; // @[executor.scala 290:56]
  wire [7:0] _GEN_942 = 8'h4 < length_0 ? _GEN_846 : _GEN_750; // @[executor.scala 290:56]
  wire [7:0] _GEN_943 = 8'h4 < length_0 ? _GEN_847 : _GEN_751; // @[executor.scala 290:56]
  wire [7:0] _GEN_944 = 8'h4 < length_0 ? _GEN_848 : _GEN_752; // @[executor.scala 290:56]
  wire [7:0] _GEN_945 = 8'h4 < length_0 ? _GEN_849 : _GEN_753; // @[executor.scala 290:56]
  wire [7:0] _GEN_946 = 8'h4 < length_0 ? _GEN_850 : _GEN_754; // @[executor.scala 290:56]
  wire [7:0] _GEN_947 = 8'h4 < length_0 ? _GEN_851 : _GEN_755; // @[executor.scala 290:56]
  wire [7:0] _GEN_948 = 8'h4 < length_0 ? _GEN_852 : _GEN_756; // @[executor.scala 290:56]
  wire [7:0] _GEN_949 = 8'h4 < length_0 ? _GEN_853 : _GEN_757; // @[executor.scala 290:56]
  wire [7:0] _GEN_950 = 8'h4 < length_0 ? _GEN_854 : _GEN_758; // @[executor.scala 290:56]
  wire [7:0] _GEN_951 = 8'h4 < length_0 ? _GEN_855 : _GEN_759; // @[executor.scala 290:56]
  wire [7:0] _GEN_952 = 8'h4 < length_0 ? _GEN_856 : _GEN_760; // @[executor.scala 290:56]
  wire [7:0] _GEN_953 = 8'h4 < length_0 ? _GEN_857 : _GEN_761; // @[executor.scala 290:56]
  wire [7:0] _GEN_954 = 8'h4 < length_0 ? _GEN_858 : _GEN_762; // @[executor.scala 290:56]
  wire [7:0] _GEN_955 = 8'h4 < length_0 ? _GEN_859 : _GEN_763; // @[executor.scala 290:56]
  wire [7:0] _GEN_956 = 8'h4 < length_0 ? _GEN_860 : _GEN_764; // @[executor.scala 290:56]
  wire [7:0] _GEN_957 = 8'h4 < length_0 ? _GEN_861 : _GEN_765; // @[executor.scala 290:56]
  wire [7:0] _GEN_958 = 8'h4 < length_0 ? _GEN_862 : _GEN_766; // @[executor.scala 290:56]
  wire [7:0] _GEN_959 = 8'h4 < length_0 ? _GEN_863 : _GEN_767; // @[executor.scala 290:56]
  wire [7:0] field_byte_5 = field_0[23:16]; // @[executor.scala 287:53]
  wire [7:0] total_offset_5 = offset_0 + 8'h5; // @[executor.scala 289:53]
  wire [7:0] _GEN_960 = 7'h0 == total_offset_5[6:0] ? field_byte_5 : _GEN_864; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_961 = 7'h1 == total_offset_5[6:0] ? field_byte_5 : _GEN_865; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_962 = 7'h2 == total_offset_5[6:0] ? field_byte_5 : _GEN_866; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_963 = 7'h3 == total_offset_5[6:0] ? field_byte_5 : _GEN_867; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_964 = 7'h4 == total_offset_5[6:0] ? field_byte_5 : _GEN_868; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_965 = 7'h5 == total_offset_5[6:0] ? field_byte_5 : _GEN_869; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_966 = 7'h6 == total_offset_5[6:0] ? field_byte_5 : _GEN_870; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_967 = 7'h7 == total_offset_5[6:0] ? field_byte_5 : _GEN_871; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_968 = 7'h8 == total_offset_5[6:0] ? field_byte_5 : _GEN_872; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_969 = 7'h9 == total_offset_5[6:0] ? field_byte_5 : _GEN_873; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_970 = 7'ha == total_offset_5[6:0] ? field_byte_5 : _GEN_874; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_971 = 7'hb == total_offset_5[6:0] ? field_byte_5 : _GEN_875; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_972 = 7'hc == total_offset_5[6:0] ? field_byte_5 : _GEN_876; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_973 = 7'hd == total_offset_5[6:0] ? field_byte_5 : _GEN_877; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_974 = 7'he == total_offset_5[6:0] ? field_byte_5 : _GEN_878; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_975 = 7'hf == total_offset_5[6:0] ? field_byte_5 : _GEN_879; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_976 = 7'h10 == total_offset_5[6:0] ? field_byte_5 : _GEN_880; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_977 = 7'h11 == total_offset_5[6:0] ? field_byte_5 : _GEN_881; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_978 = 7'h12 == total_offset_5[6:0] ? field_byte_5 : _GEN_882; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_979 = 7'h13 == total_offset_5[6:0] ? field_byte_5 : _GEN_883; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_980 = 7'h14 == total_offset_5[6:0] ? field_byte_5 : _GEN_884; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_981 = 7'h15 == total_offset_5[6:0] ? field_byte_5 : _GEN_885; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_982 = 7'h16 == total_offset_5[6:0] ? field_byte_5 : _GEN_886; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_983 = 7'h17 == total_offset_5[6:0] ? field_byte_5 : _GEN_887; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_984 = 7'h18 == total_offset_5[6:0] ? field_byte_5 : _GEN_888; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_985 = 7'h19 == total_offset_5[6:0] ? field_byte_5 : _GEN_889; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_986 = 7'h1a == total_offset_5[6:0] ? field_byte_5 : _GEN_890; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_987 = 7'h1b == total_offset_5[6:0] ? field_byte_5 : _GEN_891; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_988 = 7'h1c == total_offset_5[6:0] ? field_byte_5 : _GEN_892; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_989 = 7'h1d == total_offset_5[6:0] ? field_byte_5 : _GEN_893; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_990 = 7'h1e == total_offset_5[6:0] ? field_byte_5 : _GEN_894; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_991 = 7'h1f == total_offset_5[6:0] ? field_byte_5 : _GEN_895; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_992 = 7'h20 == total_offset_5[6:0] ? field_byte_5 : _GEN_896; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_993 = 7'h21 == total_offset_5[6:0] ? field_byte_5 : _GEN_897; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_994 = 7'h22 == total_offset_5[6:0] ? field_byte_5 : _GEN_898; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_995 = 7'h23 == total_offset_5[6:0] ? field_byte_5 : _GEN_899; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_996 = 7'h24 == total_offset_5[6:0] ? field_byte_5 : _GEN_900; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_997 = 7'h25 == total_offset_5[6:0] ? field_byte_5 : _GEN_901; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_998 = 7'h26 == total_offset_5[6:0] ? field_byte_5 : _GEN_902; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_999 = 7'h27 == total_offset_5[6:0] ? field_byte_5 : _GEN_903; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1000 = 7'h28 == total_offset_5[6:0] ? field_byte_5 : _GEN_904; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1001 = 7'h29 == total_offset_5[6:0] ? field_byte_5 : _GEN_905; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1002 = 7'h2a == total_offset_5[6:0] ? field_byte_5 : _GEN_906; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1003 = 7'h2b == total_offset_5[6:0] ? field_byte_5 : _GEN_907; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1004 = 7'h2c == total_offset_5[6:0] ? field_byte_5 : _GEN_908; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1005 = 7'h2d == total_offset_5[6:0] ? field_byte_5 : _GEN_909; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1006 = 7'h2e == total_offset_5[6:0] ? field_byte_5 : _GEN_910; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1007 = 7'h2f == total_offset_5[6:0] ? field_byte_5 : _GEN_911; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1008 = 7'h30 == total_offset_5[6:0] ? field_byte_5 : _GEN_912; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1009 = 7'h31 == total_offset_5[6:0] ? field_byte_5 : _GEN_913; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1010 = 7'h32 == total_offset_5[6:0] ? field_byte_5 : _GEN_914; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1011 = 7'h33 == total_offset_5[6:0] ? field_byte_5 : _GEN_915; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1012 = 7'h34 == total_offset_5[6:0] ? field_byte_5 : _GEN_916; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1013 = 7'h35 == total_offset_5[6:0] ? field_byte_5 : _GEN_917; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1014 = 7'h36 == total_offset_5[6:0] ? field_byte_5 : _GEN_918; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1015 = 7'h37 == total_offset_5[6:0] ? field_byte_5 : _GEN_919; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1016 = 7'h38 == total_offset_5[6:0] ? field_byte_5 : _GEN_920; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1017 = 7'h39 == total_offset_5[6:0] ? field_byte_5 : _GEN_921; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1018 = 7'h3a == total_offset_5[6:0] ? field_byte_5 : _GEN_922; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1019 = 7'h3b == total_offset_5[6:0] ? field_byte_5 : _GEN_923; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1020 = 7'h3c == total_offset_5[6:0] ? field_byte_5 : _GEN_924; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1021 = 7'h3d == total_offset_5[6:0] ? field_byte_5 : _GEN_925; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1022 = 7'h3e == total_offset_5[6:0] ? field_byte_5 : _GEN_926; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1023 = 7'h3f == total_offset_5[6:0] ? field_byte_5 : _GEN_927; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1024 = 7'h40 == total_offset_5[6:0] ? field_byte_5 : _GEN_928; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1025 = 7'h41 == total_offset_5[6:0] ? field_byte_5 : _GEN_929; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1026 = 7'h42 == total_offset_5[6:0] ? field_byte_5 : _GEN_930; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1027 = 7'h43 == total_offset_5[6:0] ? field_byte_5 : _GEN_931; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1028 = 7'h44 == total_offset_5[6:0] ? field_byte_5 : _GEN_932; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1029 = 7'h45 == total_offset_5[6:0] ? field_byte_5 : _GEN_933; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1030 = 7'h46 == total_offset_5[6:0] ? field_byte_5 : _GEN_934; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1031 = 7'h47 == total_offset_5[6:0] ? field_byte_5 : _GEN_935; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1032 = 7'h48 == total_offset_5[6:0] ? field_byte_5 : _GEN_936; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1033 = 7'h49 == total_offset_5[6:0] ? field_byte_5 : _GEN_937; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1034 = 7'h4a == total_offset_5[6:0] ? field_byte_5 : _GEN_938; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1035 = 7'h4b == total_offset_5[6:0] ? field_byte_5 : _GEN_939; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1036 = 7'h4c == total_offset_5[6:0] ? field_byte_5 : _GEN_940; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1037 = 7'h4d == total_offset_5[6:0] ? field_byte_5 : _GEN_941; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1038 = 7'h4e == total_offset_5[6:0] ? field_byte_5 : _GEN_942; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1039 = 7'h4f == total_offset_5[6:0] ? field_byte_5 : _GEN_943; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1040 = 7'h50 == total_offset_5[6:0] ? field_byte_5 : _GEN_944; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1041 = 7'h51 == total_offset_5[6:0] ? field_byte_5 : _GEN_945; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1042 = 7'h52 == total_offset_5[6:0] ? field_byte_5 : _GEN_946; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1043 = 7'h53 == total_offset_5[6:0] ? field_byte_5 : _GEN_947; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1044 = 7'h54 == total_offset_5[6:0] ? field_byte_5 : _GEN_948; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1045 = 7'h55 == total_offset_5[6:0] ? field_byte_5 : _GEN_949; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1046 = 7'h56 == total_offset_5[6:0] ? field_byte_5 : _GEN_950; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1047 = 7'h57 == total_offset_5[6:0] ? field_byte_5 : _GEN_951; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1048 = 7'h58 == total_offset_5[6:0] ? field_byte_5 : _GEN_952; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1049 = 7'h59 == total_offset_5[6:0] ? field_byte_5 : _GEN_953; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1050 = 7'h5a == total_offset_5[6:0] ? field_byte_5 : _GEN_954; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1051 = 7'h5b == total_offset_5[6:0] ? field_byte_5 : _GEN_955; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1052 = 7'h5c == total_offset_5[6:0] ? field_byte_5 : _GEN_956; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1053 = 7'h5d == total_offset_5[6:0] ? field_byte_5 : _GEN_957; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1054 = 7'h5e == total_offset_5[6:0] ? field_byte_5 : _GEN_958; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1055 = 7'h5f == total_offset_5[6:0] ? field_byte_5 : _GEN_959; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1056 = 8'h5 < length_0 ? _GEN_960 : _GEN_864; // @[executor.scala 290:56]
  wire [7:0] _GEN_1057 = 8'h5 < length_0 ? _GEN_961 : _GEN_865; // @[executor.scala 290:56]
  wire [7:0] _GEN_1058 = 8'h5 < length_0 ? _GEN_962 : _GEN_866; // @[executor.scala 290:56]
  wire [7:0] _GEN_1059 = 8'h5 < length_0 ? _GEN_963 : _GEN_867; // @[executor.scala 290:56]
  wire [7:0] _GEN_1060 = 8'h5 < length_0 ? _GEN_964 : _GEN_868; // @[executor.scala 290:56]
  wire [7:0] _GEN_1061 = 8'h5 < length_0 ? _GEN_965 : _GEN_869; // @[executor.scala 290:56]
  wire [7:0] _GEN_1062 = 8'h5 < length_0 ? _GEN_966 : _GEN_870; // @[executor.scala 290:56]
  wire [7:0] _GEN_1063 = 8'h5 < length_0 ? _GEN_967 : _GEN_871; // @[executor.scala 290:56]
  wire [7:0] _GEN_1064 = 8'h5 < length_0 ? _GEN_968 : _GEN_872; // @[executor.scala 290:56]
  wire [7:0] _GEN_1065 = 8'h5 < length_0 ? _GEN_969 : _GEN_873; // @[executor.scala 290:56]
  wire [7:0] _GEN_1066 = 8'h5 < length_0 ? _GEN_970 : _GEN_874; // @[executor.scala 290:56]
  wire [7:0] _GEN_1067 = 8'h5 < length_0 ? _GEN_971 : _GEN_875; // @[executor.scala 290:56]
  wire [7:0] _GEN_1068 = 8'h5 < length_0 ? _GEN_972 : _GEN_876; // @[executor.scala 290:56]
  wire [7:0] _GEN_1069 = 8'h5 < length_0 ? _GEN_973 : _GEN_877; // @[executor.scala 290:56]
  wire [7:0] _GEN_1070 = 8'h5 < length_0 ? _GEN_974 : _GEN_878; // @[executor.scala 290:56]
  wire [7:0] _GEN_1071 = 8'h5 < length_0 ? _GEN_975 : _GEN_879; // @[executor.scala 290:56]
  wire [7:0] _GEN_1072 = 8'h5 < length_0 ? _GEN_976 : _GEN_880; // @[executor.scala 290:56]
  wire [7:0] _GEN_1073 = 8'h5 < length_0 ? _GEN_977 : _GEN_881; // @[executor.scala 290:56]
  wire [7:0] _GEN_1074 = 8'h5 < length_0 ? _GEN_978 : _GEN_882; // @[executor.scala 290:56]
  wire [7:0] _GEN_1075 = 8'h5 < length_0 ? _GEN_979 : _GEN_883; // @[executor.scala 290:56]
  wire [7:0] _GEN_1076 = 8'h5 < length_0 ? _GEN_980 : _GEN_884; // @[executor.scala 290:56]
  wire [7:0] _GEN_1077 = 8'h5 < length_0 ? _GEN_981 : _GEN_885; // @[executor.scala 290:56]
  wire [7:0] _GEN_1078 = 8'h5 < length_0 ? _GEN_982 : _GEN_886; // @[executor.scala 290:56]
  wire [7:0] _GEN_1079 = 8'h5 < length_0 ? _GEN_983 : _GEN_887; // @[executor.scala 290:56]
  wire [7:0] _GEN_1080 = 8'h5 < length_0 ? _GEN_984 : _GEN_888; // @[executor.scala 290:56]
  wire [7:0] _GEN_1081 = 8'h5 < length_0 ? _GEN_985 : _GEN_889; // @[executor.scala 290:56]
  wire [7:0] _GEN_1082 = 8'h5 < length_0 ? _GEN_986 : _GEN_890; // @[executor.scala 290:56]
  wire [7:0] _GEN_1083 = 8'h5 < length_0 ? _GEN_987 : _GEN_891; // @[executor.scala 290:56]
  wire [7:0] _GEN_1084 = 8'h5 < length_0 ? _GEN_988 : _GEN_892; // @[executor.scala 290:56]
  wire [7:0] _GEN_1085 = 8'h5 < length_0 ? _GEN_989 : _GEN_893; // @[executor.scala 290:56]
  wire [7:0] _GEN_1086 = 8'h5 < length_0 ? _GEN_990 : _GEN_894; // @[executor.scala 290:56]
  wire [7:0] _GEN_1087 = 8'h5 < length_0 ? _GEN_991 : _GEN_895; // @[executor.scala 290:56]
  wire [7:0] _GEN_1088 = 8'h5 < length_0 ? _GEN_992 : _GEN_896; // @[executor.scala 290:56]
  wire [7:0] _GEN_1089 = 8'h5 < length_0 ? _GEN_993 : _GEN_897; // @[executor.scala 290:56]
  wire [7:0] _GEN_1090 = 8'h5 < length_0 ? _GEN_994 : _GEN_898; // @[executor.scala 290:56]
  wire [7:0] _GEN_1091 = 8'h5 < length_0 ? _GEN_995 : _GEN_899; // @[executor.scala 290:56]
  wire [7:0] _GEN_1092 = 8'h5 < length_0 ? _GEN_996 : _GEN_900; // @[executor.scala 290:56]
  wire [7:0] _GEN_1093 = 8'h5 < length_0 ? _GEN_997 : _GEN_901; // @[executor.scala 290:56]
  wire [7:0] _GEN_1094 = 8'h5 < length_0 ? _GEN_998 : _GEN_902; // @[executor.scala 290:56]
  wire [7:0] _GEN_1095 = 8'h5 < length_0 ? _GEN_999 : _GEN_903; // @[executor.scala 290:56]
  wire [7:0] _GEN_1096 = 8'h5 < length_0 ? _GEN_1000 : _GEN_904; // @[executor.scala 290:56]
  wire [7:0] _GEN_1097 = 8'h5 < length_0 ? _GEN_1001 : _GEN_905; // @[executor.scala 290:56]
  wire [7:0] _GEN_1098 = 8'h5 < length_0 ? _GEN_1002 : _GEN_906; // @[executor.scala 290:56]
  wire [7:0] _GEN_1099 = 8'h5 < length_0 ? _GEN_1003 : _GEN_907; // @[executor.scala 290:56]
  wire [7:0] _GEN_1100 = 8'h5 < length_0 ? _GEN_1004 : _GEN_908; // @[executor.scala 290:56]
  wire [7:0] _GEN_1101 = 8'h5 < length_0 ? _GEN_1005 : _GEN_909; // @[executor.scala 290:56]
  wire [7:0] _GEN_1102 = 8'h5 < length_0 ? _GEN_1006 : _GEN_910; // @[executor.scala 290:56]
  wire [7:0] _GEN_1103 = 8'h5 < length_0 ? _GEN_1007 : _GEN_911; // @[executor.scala 290:56]
  wire [7:0] _GEN_1104 = 8'h5 < length_0 ? _GEN_1008 : _GEN_912; // @[executor.scala 290:56]
  wire [7:0] _GEN_1105 = 8'h5 < length_0 ? _GEN_1009 : _GEN_913; // @[executor.scala 290:56]
  wire [7:0] _GEN_1106 = 8'h5 < length_0 ? _GEN_1010 : _GEN_914; // @[executor.scala 290:56]
  wire [7:0] _GEN_1107 = 8'h5 < length_0 ? _GEN_1011 : _GEN_915; // @[executor.scala 290:56]
  wire [7:0] _GEN_1108 = 8'h5 < length_0 ? _GEN_1012 : _GEN_916; // @[executor.scala 290:56]
  wire [7:0] _GEN_1109 = 8'h5 < length_0 ? _GEN_1013 : _GEN_917; // @[executor.scala 290:56]
  wire [7:0] _GEN_1110 = 8'h5 < length_0 ? _GEN_1014 : _GEN_918; // @[executor.scala 290:56]
  wire [7:0] _GEN_1111 = 8'h5 < length_0 ? _GEN_1015 : _GEN_919; // @[executor.scala 290:56]
  wire [7:0] _GEN_1112 = 8'h5 < length_0 ? _GEN_1016 : _GEN_920; // @[executor.scala 290:56]
  wire [7:0] _GEN_1113 = 8'h5 < length_0 ? _GEN_1017 : _GEN_921; // @[executor.scala 290:56]
  wire [7:0] _GEN_1114 = 8'h5 < length_0 ? _GEN_1018 : _GEN_922; // @[executor.scala 290:56]
  wire [7:0] _GEN_1115 = 8'h5 < length_0 ? _GEN_1019 : _GEN_923; // @[executor.scala 290:56]
  wire [7:0] _GEN_1116 = 8'h5 < length_0 ? _GEN_1020 : _GEN_924; // @[executor.scala 290:56]
  wire [7:0] _GEN_1117 = 8'h5 < length_0 ? _GEN_1021 : _GEN_925; // @[executor.scala 290:56]
  wire [7:0] _GEN_1118 = 8'h5 < length_0 ? _GEN_1022 : _GEN_926; // @[executor.scala 290:56]
  wire [7:0] _GEN_1119 = 8'h5 < length_0 ? _GEN_1023 : _GEN_927; // @[executor.scala 290:56]
  wire [7:0] _GEN_1120 = 8'h5 < length_0 ? _GEN_1024 : _GEN_928; // @[executor.scala 290:56]
  wire [7:0] _GEN_1121 = 8'h5 < length_0 ? _GEN_1025 : _GEN_929; // @[executor.scala 290:56]
  wire [7:0] _GEN_1122 = 8'h5 < length_0 ? _GEN_1026 : _GEN_930; // @[executor.scala 290:56]
  wire [7:0] _GEN_1123 = 8'h5 < length_0 ? _GEN_1027 : _GEN_931; // @[executor.scala 290:56]
  wire [7:0] _GEN_1124 = 8'h5 < length_0 ? _GEN_1028 : _GEN_932; // @[executor.scala 290:56]
  wire [7:0] _GEN_1125 = 8'h5 < length_0 ? _GEN_1029 : _GEN_933; // @[executor.scala 290:56]
  wire [7:0] _GEN_1126 = 8'h5 < length_0 ? _GEN_1030 : _GEN_934; // @[executor.scala 290:56]
  wire [7:0] _GEN_1127 = 8'h5 < length_0 ? _GEN_1031 : _GEN_935; // @[executor.scala 290:56]
  wire [7:0] _GEN_1128 = 8'h5 < length_0 ? _GEN_1032 : _GEN_936; // @[executor.scala 290:56]
  wire [7:0] _GEN_1129 = 8'h5 < length_0 ? _GEN_1033 : _GEN_937; // @[executor.scala 290:56]
  wire [7:0] _GEN_1130 = 8'h5 < length_0 ? _GEN_1034 : _GEN_938; // @[executor.scala 290:56]
  wire [7:0] _GEN_1131 = 8'h5 < length_0 ? _GEN_1035 : _GEN_939; // @[executor.scala 290:56]
  wire [7:0] _GEN_1132 = 8'h5 < length_0 ? _GEN_1036 : _GEN_940; // @[executor.scala 290:56]
  wire [7:0] _GEN_1133 = 8'h5 < length_0 ? _GEN_1037 : _GEN_941; // @[executor.scala 290:56]
  wire [7:0] _GEN_1134 = 8'h5 < length_0 ? _GEN_1038 : _GEN_942; // @[executor.scala 290:56]
  wire [7:0] _GEN_1135 = 8'h5 < length_0 ? _GEN_1039 : _GEN_943; // @[executor.scala 290:56]
  wire [7:0] _GEN_1136 = 8'h5 < length_0 ? _GEN_1040 : _GEN_944; // @[executor.scala 290:56]
  wire [7:0] _GEN_1137 = 8'h5 < length_0 ? _GEN_1041 : _GEN_945; // @[executor.scala 290:56]
  wire [7:0] _GEN_1138 = 8'h5 < length_0 ? _GEN_1042 : _GEN_946; // @[executor.scala 290:56]
  wire [7:0] _GEN_1139 = 8'h5 < length_0 ? _GEN_1043 : _GEN_947; // @[executor.scala 290:56]
  wire [7:0] _GEN_1140 = 8'h5 < length_0 ? _GEN_1044 : _GEN_948; // @[executor.scala 290:56]
  wire [7:0] _GEN_1141 = 8'h5 < length_0 ? _GEN_1045 : _GEN_949; // @[executor.scala 290:56]
  wire [7:0] _GEN_1142 = 8'h5 < length_0 ? _GEN_1046 : _GEN_950; // @[executor.scala 290:56]
  wire [7:0] _GEN_1143 = 8'h5 < length_0 ? _GEN_1047 : _GEN_951; // @[executor.scala 290:56]
  wire [7:0] _GEN_1144 = 8'h5 < length_0 ? _GEN_1048 : _GEN_952; // @[executor.scala 290:56]
  wire [7:0] _GEN_1145 = 8'h5 < length_0 ? _GEN_1049 : _GEN_953; // @[executor.scala 290:56]
  wire [7:0] _GEN_1146 = 8'h5 < length_0 ? _GEN_1050 : _GEN_954; // @[executor.scala 290:56]
  wire [7:0] _GEN_1147 = 8'h5 < length_0 ? _GEN_1051 : _GEN_955; // @[executor.scala 290:56]
  wire [7:0] _GEN_1148 = 8'h5 < length_0 ? _GEN_1052 : _GEN_956; // @[executor.scala 290:56]
  wire [7:0] _GEN_1149 = 8'h5 < length_0 ? _GEN_1053 : _GEN_957; // @[executor.scala 290:56]
  wire [7:0] _GEN_1150 = 8'h5 < length_0 ? _GEN_1054 : _GEN_958; // @[executor.scala 290:56]
  wire [7:0] _GEN_1151 = 8'h5 < length_0 ? _GEN_1055 : _GEN_959; // @[executor.scala 290:56]
  wire [7:0] field_byte_6 = field_0[15:8]; // @[executor.scala 287:53]
  wire [7:0] total_offset_6 = offset_0 + 8'h6; // @[executor.scala 289:53]
  wire [7:0] _GEN_1152 = 7'h0 == total_offset_6[6:0] ? field_byte_6 : _GEN_1056; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1153 = 7'h1 == total_offset_6[6:0] ? field_byte_6 : _GEN_1057; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1154 = 7'h2 == total_offset_6[6:0] ? field_byte_6 : _GEN_1058; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1155 = 7'h3 == total_offset_6[6:0] ? field_byte_6 : _GEN_1059; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1156 = 7'h4 == total_offset_6[6:0] ? field_byte_6 : _GEN_1060; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1157 = 7'h5 == total_offset_6[6:0] ? field_byte_6 : _GEN_1061; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1158 = 7'h6 == total_offset_6[6:0] ? field_byte_6 : _GEN_1062; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1159 = 7'h7 == total_offset_6[6:0] ? field_byte_6 : _GEN_1063; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1160 = 7'h8 == total_offset_6[6:0] ? field_byte_6 : _GEN_1064; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1161 = 7'h9 == total_offset_6[6:0] ? field_byte_6 : _GEN_1065; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1162 = 7'ha == total_offset_6[6:0] ? field_byte_6 : _GEN_1066; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1163 = 7'hb == total_offset_6[6:0] ? field_byte_6 : _GEN_1067; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1164 = 7'hc == total_offset_6[6:0] ? field_byte_6 : _GEN_1068; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1165 = 7'hd == total_offset_6[6:0] ? field_byte_6 : _GEN_1069; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1166 = 7'he == total_offset_6[6:0] ? field_byte_6 : _GEN_1070; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1167 = 7'hf == total_offset_6[6:0] ? field_byte_6 : _GEN_1071; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1168 = 7'h10 == total_offset_6[6:0] ? field_byte_6 : _GEN_1072; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1169 = 7'h11 == total_offset_6[6:0] ? field_byte_6 : _GEN_1073; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1170 = 7'h12 == total_offset_6[6:0] ? field_byte_6 : _GEN_1074; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1171 = 7'h13 == total_offset_6[6:0] ? field_byte_6 : _GEN_1075; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1172 = 7'h14 == total_offset_6[6:0] ? field_byte_6 : _GEN_1076; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1173 = 7'h15 == total_offset_6[6:0] ? field_byte_6 : _GEN_1077; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1174 = 7'h16 == total_offset_6[6:0] ? field_byte_6 : _GEN_1078; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1175 = 7'h17 == total_offset_6[6:0] ? field_byte_6 : _GEN_1079; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1176 = 7'h18 == total_offset_6[6:0] ? field_byte_6 : _GEN_1080; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1177 = 7'h19 == total_offset_6[6:0] ? field_byte_6 : _GEN_1081; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1178 = 7'h1a == total_offset_6[6:0] ? field_byte_6 : _GEN_1082; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1179 = 7'h1b == total_offset_6[6:0] ? field_byte_6 : _GEN_1083; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1180 = 7'h1c == total_offset_6[6:0] ? field_byte_6 : _GEN_1084; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1181 = 7'h1d == total_offset_6[6:0] ? field_byte_6 : _GEN_1085; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1182 = 7'h1e == total_offset_6[6:0] ? field_byte_6 : _GEN_1086; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1183 = 7'h1f == total_offset_6[6:0] ? field_byte_6 : _GEN_1087; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1184 = 7'h20 == total_offset_6[6:0] ? field_byte_6 : _GEN_1088; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1185 = 7'h21 == total_offset_6[6:0] ? field_byte_6 : _GEN_1089; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1186 = 7'h22 == total_offset_6[6:0] ? field_byte_6 : _GEN_1090; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1187 = 7'h23 == total_offset_6[6:0] ? field_byte_6 : _GEN_1091; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1188 = 7'h24 == total_offset_6[6:0] ? field_byte_6 : _GEN_1092; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1189 = 7'h25 == total_offset_6[6:0] ? field_byte_6 : _GEN_1093; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1190 = 7'h26 == total_offset_6[6:0] ? field_byte_6 : _GEN_1094; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1191 = 7'h27 == total_offset_6[6:0] ? field_byte_6 : _GEN_1095; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1192 = 7'h28 == total_offset_6[6:0] ? field_byte_6 : _GEN_1096; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1193 = 7'h29 == total_offset_6[6:0] ? field_byte_6 : _GEN_1097; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1194 = 7'h2a == total_offset_6[6:0] ? field_byte_6 : _GEN_1098; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1195 = 7'h2b == total_offset_6[6:0] ? field_byte_6 : _GEN_1099; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1196 = 7'h2c == total_offset_6[6:0] ? field_byte_6 : _GEN_1100; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1197 = 7'h2d == total_offset_6[6:0] ? field_byte_6 : _GEN_1101; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1198 = 7'h2e == total_offset_6[6:0] ? field_byte_6 : _GEN_1102; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1199 = 7'h2f == total_offset_6[6:0] ? field_byte_6 : _GEN_1103; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1200 = 7'h30 == total_offset_6[6:0] ? field_byte_6 : _GEN_1104; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1201 = 7'h31 == total_offset_6[6:0] ? field_byte_6 : _GEN_1105; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1202 = 7'h32 == total_offset_6[6:0] ? field_byte_6 : _GEN_1106; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1203 = 7'h33 == total_offset_6[6:0] ? field_byte_6 : _GEN_1107; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1204 = 7'h34 == total_offset_6[6:0] ? field_byte_6 : _GEN_1108; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1205 = 7'h35 == total_offset_6[6:0] ? field_byte_6 : _GEN_1109; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1206 = 7'h36 == total_offset_6[6:0] ? field_byte_6 : _GEN_1110; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1207 = 7'h37 == total_offset_6[6:0] ? field_byte_6 : _GEN_1111; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1208 = 7'h38 == total_offset_6[6:0] ? field_byte_6 : _GEN_1112; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1209 = 7'h39 == total_offset_6[6:0] ? field_byte_6 : _GEN_1113; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1210 = 7'h3a == total_offset_6[6:0] ? field_byte_6 : _GEN_1114; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1211 = 7'h3b == total_offset_6[6:0] ? field_byte_6 : _GEN_1115; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1212 = 7'h3c == total_offset_6[6:0] ? field_byte_6 : _GEN_1116; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1213 = 7'h3d == total_offset_6[6:0] ? field_byte_6 : _GEN_1117; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1214 = 7'h3e == total_offset_6[6:0] ? field_byte_6 : _GEN_1118; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1215 = 7'h3f == total_offset_6[6:0] ? field_byte_6 : _GEN_1119; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1216 = 7'h40 == total_offset_6[6:0] ? field_byte_6 : _GEN_1120; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1217 = 7'h41 == total_offset_6[6:0] ? field_byte_6 : _GEN_1121; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1218 = 7'h42 == total_offset_6[6:0] ? field_byte_6 : _GEN_1122; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1219 = 7'h43 == total_offset_6[6:0] ? field_byte_6 : _GEN_1123; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1220 = 7'h44 == total_offset_6[6:0] ? field_byte_6 : _GEN_1124; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1221 = 7'h45 == total_offset_6[6:0] ? field_byte_6 : _GEN_1125; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1222 = 7'h46 == total_offset_6[6:0] ? field_byte_6 : _GEN_1126; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1223 = 7'h47 == total_offset_6[6:0] ? field_byte_6 : _GEN_1127; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1224 = 7'h48 == total_offset_6[6:0] ? field_byte_6 : _GEN_1128; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1225 = 7'h49 == total_offset_6[6:0] ? field_byte_6 : _GEN_1129; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1226 = 7'h4a == total_offset_6[6:0] ? field_byte_6 : _GEN_1130; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1227 = 7'h4b == total_offset_6[6:0] ? field_byte_6 : _GEN_1131; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1228 = 7'h4c == total_offset_6[6:0] ? field_byte_6 : _GEN_1132; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1229 = 7'h4d == total_offset_6[6:0] ? field_byte_6 : _GEN_1133; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1230 = 7'h4e == total_offset_6[6:0] ? field_byte_6 : _GEN_1134; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1231 = 7'h4f == total_offset_6[6:0] ? field_byte_6 : _GEN_1135; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1232 = 7'h50 == total_offset_6[6:0] ? field_byte_6 : _GEN_1136; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1233 = 7'h51 == total_offset_6[6:0] ? field_byte_6 : _GEN_1137; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1234 = 7'h52 == total_offset_6[6:0] ? field_byte_6 : _GEN_1138; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1235 = 7'h53 == total_offset_6[6:0] ? field_byte_6 : _GEN_1139; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1236 = 7'h54 == total_offset_6[6:0] ? field_byte_6 : _GEN_1140; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1237 = 7'h55 == total_offset_6[6:0] ? field_byte_6 : _GEN_1141; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1238 = 7'h56 == total_offset_6[6:0] ? field_byte_6 : _GEN_1142; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1239 = 7'h57 == total_offset_6[6:0] ? field_byte_6 : _GEN_1143; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1240 = 7'h58 == total_offset_6[6:0] ? field_byte_6 : _GEN_1144; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1241 = 7'h59 == total_offset_6[6:0] ? field_byte_6 : _GEN_1145; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1242 = 7'h5a == total_offset_6[6:0] ? field_byte_6 : _GEN_1146; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1243 = 7'h5b == total_offset_6[6:0] ? field_byte_6 : _GEN_1147; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1244 = 7'h5c == total_offset_6[6:0] ? field_byte_6 : _GEN_1148; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1245 = 7'h5d == total_offset_6[6:0] ? field_byte_6 : _GEN_1149; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1246 = 7'h5e == total_offset_6[6:0] ? field_byte_6 : _GEN_1150; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1247 = 7'h5f == total_offset_6[6:0] ? field_byte_6 : _GEN_1151; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1248 = 8'h6 < length_0 ? _GEN_1152 : _GEN_1056; // @[executor.scala 290:56]
  wire [7:0] _GEN_1249 = 8'h6 < length_0 ? _GEN_1153 : _GEN_1057; // @[executor.scala 290:56]
  wire [7:0] _GEN_1250 = 8'h6 < length_0 ? _GEN_1154 : _GEN_1058; // @[executor.scala 290:56]
  wire [7:0] _GEN_1251 = 8'h6 < length_0 ? _GEN_1155 : _GEN_1059; // @[executor.scala 290:56]
  wire [7:0] _GEN_1252 = 8'h6 < length_0 ? _GEN_1156 : _GEN_1060; // @[executor.scala 290:56]
  wire [7:0] _GEN_1253 = 8'h6 < length_0 ? _GEN_1157 : _GEN_1061; // @[executor.scala 290:56]
  wire [7:0] _GEN_1254 = 8'h6 < length_0 ? _GEN_1158 : _GEN_1062; // @[executor.scala 290:56]
  wire [7:0] _GEN_1255 = 8'h6 < length_0 ? _GEN_1159 : _GEN_1063; // @[executor.scala 290:56]
  wire [7:0] _GEN_1256 = 8'h6 < length_0 ? _GEN_1160 : _GEN_1064; // @[executor.scala 290:56]
  wire [7:0] _GEN_1257 = 8'h6 < length_0 ? _GEN_1161 : _GEN_1065; // @[executor.scala 290:56]
  wire [7:0] _GEN_1258 = 8'h6 < length_0 ? _GEN_1162 : _GEN_1066; // @[executor.scala 290:56]
  wire [7:0] _GEN_1259 = 8'h6 < length_0 ? _GEN_1163 : _GEN_1067; // @[executor.scala 290:56]
  wire [7:0] _GEN_1260 = 8'h6 < length_0 ? _GEN_1164 : _GEN_1068; // @[executor.scala 290:56]
  wire [7:0] _GEN_1261 = 8'h6 < length_0 ? _GEN_1165 : _GEN_1069; // @[executor.scala 290:56]
  wire [7:0] _GEN_1262 = 8'h6 < length_0 ? _GEN_1166 : _GEN_1070; // @[executor.scala 290:56]
  wire [7:0] _GEN_1263 = 8'h6 < length_0 ? _GEN_1167 : _GEN_1071; // @[executor.scala 290:56]
  wire [7:0] _GEN_1264 = 8'h6 < length_0 ? _GEN_1168 : _GEN_1072; // @[executor.scala 290:56]
  wire [7:0] _GEN_1265 = 8'h6 < length_0 ? _GEN_1169 : _GEN_1073; // @[executor.scala 290:56]
  wire [7:0] _GEN_1266 = 8'h6 < length_0 ? _GEN_1170 : _GEN_1074; // @[executor.scala 290:56]
  wire [7:0] _GEN_1267 = 8'h6 < length_0 ? _GEN_1171 : _GEN_1075; // @[executor.scala 290:56]
  wire [7:0] _GEN_1268 = 8'h6 < length_0 ? _GEN_1172 : _GEN_1076; // @[executor.scala 290:56]
  wire [7:0] _GEN_1269 = 8'h6 < length_0 ? _GEN_1173 : _GEN_1077; // @[executor.scala 290:56]
  wire [7:0] _GEN_1270 = 8'h6 < length_0 ? _GEN_1174 : _GEN_1078; // @[executor.scala 290:56]
  wire [7:0] _GEN_1271 = 8'h6 < length_0 ? _GEN_1175 : _GEN_1079; // @[executor.scala 290:56]
  wire [7:0] _GEN_1272 = 8'h6 < length_0 ? _GEN_1176 : _GEN_1080; // @[executor.scala 290:56]
  wire [7:0] _GEN_1273 = 8'h6 < length_0 ? _GEN_1177 : _GEN_1081; // @[executor.scala 290:56]
  wire [7:0] _GEN_1274 = 8'h6 < length_0 ? _GEN_1178 : _GEN_1082; // @[executor.scala 290:56]
  wire [7:0] _GEN_1275 = 8'h6 < length_0 ? _GEN_1179 : _GEN_1083; // @[executor.scala 290:56]
  wire [7:0] _GEN_1276 = 8'h6 < length_0 ? _GEN_1180 : _GEN_1084; // @[executor.scala 290:56]
  wire [7:0] _GEN_1277 = 8'h6 < length_0 ? _GEN_1181 : _GEN_1085; // @[executor.scala 290:56]
  wire [7:0] _GEN_1278 = 8'h6 < length_0 ? _GEN_1182 : _GEN_1086; // @[executor.scala 290:56]
  wire [7:0] _GEN_1279 = 8'h6 < length_0 ? _GEN_1183 : _GEN_1087; // @[executor.scala 290:56]
  wire [7:0] _GEN_1280 = 8'h6 < length_0 ? _GEN_1184 : _GEN_1088; // @[executor.scala 290:56]
  wire [7:0] _GEN_1281 = 8'h6 < length_0 ? _GEN_1185 : _GEN_1089; // @[executor.scala 290:56]
  wire [7:0] _GEN_1282 = 8'h6 < length_0 ? _GEN_1186 : _GEN_1090; // @[executor.scala 290:56]
  wire [7:0] _GEN_1283 = 8'h6 < length_0 ? _GEN_1187 : _GEN_1091; // @[executor.scala 290:56]
  wire [7:0] _GEN_1284 = 8'h6 < length_0 ? _GEN_1188 : _GEN_1092; // @[executor.scala 290:56]
  wire [7:0] _GEN_1285 = 8'h6 < length_0 ? _GEN_1189 : _GEN_1093; // @[executor.scala 290:56]
  wire [7:0] _GEN_1286 = 8'h6 < length_0 ? _GEN_1190 : _GEN_1094; // @[executor.scala 290:56]
  wire [7:0] _GEN_1287 = 8'h6 < length_0 ? _GEN_1191 : _GEN_1095; // @[executor.scala 290:56]
  wire [7:0] _GEN_1288 = 8'h6 < length_0 ? _GEN_1192 : _GEN_1096; // @[executor.scala 290:56]
  wire [7:0] _GEN_1289 = 8'h6 < length_0 ? _GEN_1193 : _GEN_1097; // @[executor.scala 290:56]
  wire [7:0] _GEN_1290 = 8'h6 < length_0 ? _GEN_1194 : _GEN_1098; // @[executor.scala 290:56]
  wire [7:0] _GEN_1291 = 8'h6 < length_0 ? _GEN_1195 : _GEN_1099; // @[executor.scala 290:56]
  wire [7:0] _GEN_1292 = 8'h6 < length_0 ? _GEN_1196 : _GEN_1100; // @[executor.scala 290:56]
  wire [7:0] _GEN_1293 = 8'h6 < length_0 ? _GEN_1197 : _GEN_1101; // @[executor.scala 290:56]
  wire [7:0] _GEN_1294 = 8'h6 < length_0 ? _GEN_1198 : _GEN_1102; // @[executor.scala 290:56]
  wire [7:0] _GEN_1295 = 8'h6 < length_0 ? _GEN_1199 : _GEN_1103; // @[executor.scala 290:56]
  wire [7:0] _GEN_1296 = 8'h6 < length_0 ? _GEN_1200 : _GEN_1104; // @[executor.scala 290:56]
  wire [7:0] _GEN_1297 = 8'h6 < length_0 ? _GEN_1201 : _GEN_1105; // @[executor.scala 290:56]
  wire [7:0] _GEN_1298 = 8'h6 < length_0 ? _GEN_1202 : _GEN_1106; // @[executor.scala 290:56]
  wire [7:0] _GEN_1299 = 8'h6 < length_0 ? _GEN_1203 : _GEN_1107; // @[executor.scala 290:56]
  wire [7:0] _GEN_1300 = 8'h6 < length_0 ? _GEN_1204 : _GEN_1108; // @[executor.scala 290:56]
  wire [7:0] _GEN_1301 = 8'h6 < length_0 ? _GEN_1205 : _GEN_1109; // @[executor.scala 290:56]
  wire [7:0] _GEN_1302 = 8'h6 < length_0 ? _GEN_1206 : _GEN_1110; // @[executor.scala 290:56]
  wire [7:0] _GEN_1303 = 8'h6 < length_0 ? _GEN_1207 : _GEN_1111; // @[executor.scala 290:56]
  wire [7:0] _GEN_1304 = 8'h6 < length_0 ? _GEN_1208 : _GEN_1112; // @[executor.scala 290:56]
  wire [7:0] _GEN_1305 = 8'h6 < length_0 ? _GEN_1209 : _GEN_1113; // @[executor.scala 290:56]
  wire [7:0] _GEN_1306 = 8'h6 < length_0 ? _GEN_1210 : _GEN_1114; // @[executor.scala 290:56]
  wire [7:0] _GEN_1307 = 8'h6 < length_0 ? _GEN_1211 : _GEN_1115; // @[executor.scala 290:56]
  wire [7:0] _GEN_1308 = 8'h6 < length_0 ? _GEN_1212 : _GEN_1116; // @[executor.scala 290:56]
  wire [7:0] _GEN_1309 = 8'h6 < length_0 ? _GEN_1213 : _GEN_1117; // @[executor.scala 290:56]
  wire [7:0] _GEN_1310 = 8'h6 < length_0 ? _GEN_1214 : _GEN_1118; // @[executor.scala 290:56]
  wire [7:0] _GEN_1311 = 8'h6 < length_0 ? _GEN_1215 : _GEN_1119; // @[executor.scala 290:56]
  wire [7:0] _GEN_1312 = 8'h6 < length_0 ? _GEN_1216 : _GEN_1120; // @[executor.scala 290:56]
  wire [7:0] _GEN_1313 = 8'h6 < length_0 ? _GEN_1217 : _GEN_1121; // @[executor.scala 290:56]
  wire [7:0] _GEN_1314 = 8'h6 < length_0 ? _GEN_1218 : _GEN_1122; // @[executor.scala 290:56]
  wire [7:0] _GEN_1315 = 8'h6 < length_0 ? _GEN_1219 : _GEN_1123; // @[executor.scala 290:56]
  wire [7:0] _GEN_1316 = 8'h6 < length_0 ? _GEN_1220 : _GEN_1124; // @[executor.scala 290:56]
  wire [7:0] _GEN_1317 = 8'h6 < length_0 ? _GEN_1221 : _GEN_1125; // @[executor.scala 290:56]
  wire [7:0] _GEN_1318 = 8'h6 < length_0 ? _GEN_1222 : _GEN_1126; // @[executor.scala 290:56]
  wire [7:0] _GEN_1319 = 8'h6 < length_0 ? _GEN_1223 : _GEN_1127; // @[executor.scala 290:56]
  wire [7:0] _GEN_1320 = 8'h6 < length_0 ? _GEN_1224 : _GEN_1128; // @[executor.scala 290:56]
  wire [7:0] _GEN_1321 = 8'h6 < length_0 ? _GEN_1225 : _GEN_1129; // @[executor.scala 290:56]
  wire [7:0] _GEN_1322 = 8'h6 < length_0 ? _GEN_1226 : _GEN_1130; // @[executor.scala 290:56]
  wire [7:0] _GEN_1323 = 8'h6 < length_0 ? _GEN_1227 : _GEN_1131; // @[executor.scala 290:56]
  wire [7:0] _GEN_1324 = 8'h6 < length_0 ? _GEN_1228 : _GEN_1132; // @[executor.scala 290:56]
  wire [7:0] _GEN_1325 = 8'h6 < length_0 ? _GEN_1229 : _GEN_1133; // @[executor.scala 290:56]
  wire [7:0] _GEN_1326 = 8'h6 < length_0 ? _GEN_1230 : _GEN_1134; // @[executor.scala 290:56]
  wire [7:0] _GEN_1327 = 8'h6 < length_0 ? _GEN_1231 : _GEN_1135; // @[executor.scala 290:56]
  wire [7:0] _GEN_1328 = 8'h6 < length_0 ? _GEN_1232 : _GEN_1136; // @[executor.scala 290:56]
  wire [7:0] _GEN_1329 = 8'h6 < length_0 ? _GEN_1233 : _GEN_1137; // @[executor.scala 290:56]
  wire [7:0] _GEN_1330 = 8'h6 < length_0 ? _GEN_1234 : _GEN_1138; // @[executor.scala 290:56]
  wire [7:0] _GEN_1331 = 8'h6 < length_0 ? _GEN_1235 : _GEN_1139; // @[executor.scala 290:56]
  wire [7:0] _GEN_1332 = 8'h6 < length_0 ? _GEN_1236 : _GEN_1140; // @[executor.scala 290:56]
  wire [7:0] _GEN_1333 = 8'h6 < length_0 ? _GEN_1237 : _GEN_1141; // @[executor.scala 290:56]
  wire [7:0] _GEN_1334 = 8'h6 < length_0 ? _GEN_1238 : _GEN_1142; // @[executor.scala 290:56]
  wire [7:0] _GEN_1335 = 8'h6 < length_0 ? _GEN_1239 : _GEN_1143; // @[executor.scala 290:56]
  wire [7:0] _GEN_1336 = 8'h6 < length_0 ? _GEN_1240 : _GEN_1144; // @[executor.scala 290:56]
  wire [7:0] _GEN_1337 = 8'h6 < length_0 ? _GEN_1241 : _GEN_1145; // @[executor.scala 290:56]
  wire [7:0] _GEN_1338 = 8'h6 < length_0 ? _GEN_1242 : _GEN_1146; // @[executor.scala 290:56]
  wire [7:0] _GEN_1339 = 8'h6 < length_0 ? _GEN_1243 : _GEN_1147; // @[executor.scala 290:56]
  wire [7:0] _GEN_1340 = 8'h6 < length_0 ? _GEN_1244 : _GEN_1148; // @[executor.scala 290:56]
  wire [7:0] _GEN_1341 = 8'h6 < length_0 ? _GEN_1245 : _GEN_1149; // @[executor.scala 290:56]
  wire [7:0] _GEN_1342 = 8'h6 < length_0 ? _GEN_1246 : _GEN_1150; // @[executor.scala 290:56]
  wire [7:0] _GEN_1343 = 8'h6 < length_0 ? _GEN_1247 : _GEN_1151; // @[executor.scala 290:56]
  wire [7:0] field_byte_7 = field_0[7:0]; // @[executor.scala 287:53]
  wire [7:0] total_offset_7 = offset_0 + 8'h7; // @[executor.scala 289:53]
  wire [7:0] _GEN_1344 = 7'h0 == total_offset_7[6:0] ? field_byte_7 : _GEN_1248; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1345 = 7'h1 == total_offset_7[6:0] ? field_byte_7 : _GEN_1249; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1346 = 7'h2 == total_offset_7[6:0] ? field_byte_7 : _GEN_1250; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1347 = 7'h3 == total_offset_7[6:0] ? field_byte_7 : _GEN_1251; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1348 = 7'h4 == total_offset_7[6:0] ? field_byte_7 : _GEN_1252; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1349 = 7'h5 == total_offset_7[6:0] ? field_byte_7 : _GEN_1253; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1350 = 7'h6 == total_offset_7[6:0] ? field_byte_7 : _GEN_1254; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1351 = 7'h7 == total_offset_7[6:0] ? field_byte_7 : _GEN_1255; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1352 = 7'h8 == total_offset_7[6:0] ? field_byte_7 : _GEN_1256; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1353 = 7'h9 == total_offset_7[6:0] ? field_byte_7 : _GEN_1257; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1354 = 7'ha == total_offset_7[6:0] ? field_byte_7 : _GEN_1258; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1355 = 7'hb == total_offset_7[6:0] ? field_byte_7 : _GEN_1259; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1356 = 7'hc == total_offset_7[6:0] ? field_byte_7 : _GEN_1260; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1357 = 7'hd == total_offset_7[6:0] ? field_byte_7 : _GEN_1261; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1358 = 7'he == total_offset_7[6:0] ? field_byte_7 : _GEN_1262; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1359 = 7'hf == total_offset_7[6:0] ? field_byte_7 : _GEN_1263; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1360 = 7'h10 == total_offset_7[6:0] ? field_byte_7 : _GEN_1264; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1361 = 7'h11 == total_offset_7[6:0] ? field_byte_7 : _GEN_1265; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1362 = 7'h12 == total_offset_7[6:0] ? field_byte_7 : _GEN_1266; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1363 = 7'h13 == total_offset_7[6:0] ? field_byte_7 : _GEN_1267; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1364 = 7'h14 == total_offset_7[6:0] ? field_byte_7 : _GEN_1268; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1365 = 7'h15 == total_offset_7[6:0] ? field_byte_7 : _GEN_1269; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1366 = 7'h16 == total_offset_7[6:0] ? field_byte_7 : _GEN_1270; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1367 = 7'h17 == total_offset_7[6:0] ? field_byte_7 : _GEN_1271; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1368 = 7'h18 == total_offset_7[6:0] ? field_byte_7 : _GEN_1272; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1369 = 7'h19 == total_offset_7[6:0] ? field_byte_7 : _GEN_1273; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1370 = 7'h1a == total_offset_7[6:0] ? field_byte_7 : _GEN_1274; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1371 = 7'h1b == total_offset_7[6:0] ? field_byte_7 : _GEN_1275; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1372 = 7'h1c == total_offset_7[6:0] ? field_byte_7 : _GEN_1276; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1373 = 7'h1d == total_offset_7[6:0] ? field_byte_7 : _GEN_1277; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1374 = 7'h1e == total_offset_7[6:0] ? field_byte_7 : _GEN_1278; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1375 = 7'h1f == total_offset_7[6:0] ? field_byte_7 : _GEN_1279; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1376 = 7'h20 == total_offset_7[6:0] ? field_byte_7 : _GEN_1280; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1377 = 7'h21 == total_offset_7[6:0] ? field_byte_7 : _GEN_1281; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1378 = 7'h22 == total_offset_7[6:0] ? field_byte_7 : _GEN_1282; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1379 = 7'h23 == total_offset_7[6:0] ? field_byte_7 : _GEN_1283; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1380 = 7'h24 == total_offset_7[6:0] ? field_byte_7 : _GEN_1284; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1381 = 7'h25 == total_offset_7[6:0] ? field_byte_7 : _GEN_1285; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1382 = 7'h26 == total_offset_7[6:0] ? field_byte_7 : _GEN_1286; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1383 = 7'h27 == total_offset_7[6:0] ? field_byte_7 : _GEN_1287; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1384 = 7'h28 == total_offset_7[6:0] ? field_byte_7 : _GEN_1288; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1385 = 7'h29 == total_offset_7[6:0] ? field_byte_7 : _GEN_1289; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1386 = 7'h2a == total_offset_7[6:0] ? field_byte_7 : _GEN_1290; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1387 = 7'h2b == total_offset_7[6:0] ? field_byte_7 : _GEN_1291; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1388 = 7'h2c == total_offset_7[6:0] ? field_byte_7 : _GEN_1292; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1389 = 7'h2d == total_offset_7[6:0] ? field_byte_7 : _GEN_1293; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1390 = 7'h2e == total_offset_7[6:0] ? field_byte_7 : _GEN_1294; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1391 = 7'h2f == total_offset_7[6:0] ? field_byte_7 : _GEN_1295; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1392 = 7'h30 == total_offset_7[6:0] ? field_byte_7 : _GEN_1296; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1393 = 7'h31 == total_offset_7[6:0] ? field_byte_7 : _GEN_1297; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1394 = 7'h32 == total_offset_7[6:0] ? field_byte_7 : _GEN_1298; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1395 = 7'h33 == total_offset_7[6:0] ? field_byte_7 : _GEN_1299; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1396 = 7'h34 == total_offset_7[6:0] ? field_byte_7 : _GEN_1300; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1397 = 7'h35 == total_offset_7[6:0] ? field_byte_7 : _GEN_1301; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1398 = 7'h36 == total_offset_7[6:0] ? field_byte_7 : _GEN_1302; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1399 = 7'h37 == total_offset_7[6:0] ? field_byte_7 : _GEN_1303; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1400 = 7'h38 == total_offset_7[6:0] ? field_byte_7 : _GEN_1304; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1401 = 7'h39 == total_offset_7[6:0] ? field_byte_7 : _GEN_1305; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1402 = 7'h3a == total_offset_7[6:0] ? field_byte_7 : _GEN_1306; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1403 = 7'h3b == total_offset_7[6:0] ? field_byte_7 : _GEN_1307; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1404 = 7'h3c == total_offset_7[6:0] ? field_byte_7 : _GEN_1308; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1405 = 7'h3d == total_offset_7[6:0] ? field_byte_7 : _GEN_1309; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1406 = 7'h3e == total_offset_7[6:0] ? field_byte_7 : _GEN_1310; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1407 = 7'h3f == total_offset_7[6:0] ? field_byte_7 : _GEN_1311; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1408 = 7'h40 == total_offset_7[6:0] ? field_byte_7 : _GEN_1312; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1409 = 7'h41 == total_offset_7[6:0] ? field_byte_7 : _GEN_1313; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1410 = 7'h42 == total_offset_7[6:0] ? field_byte_7 : _GEN_1314; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1411 = 7'h43 == total_offset_7[6:0] ? field_byte_7 : _GEN_1315; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1412 = 7'h44 == total_offset_7[6:0] ? field_byte_7 : _GEN_1316; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1413 = 7'h45 == total_offset_7[6:0] ? field_byte_7 : _GEN_1317; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1414 = 7'h46 == total_offset_7[6:0] ? field_byte_7 : _GEN_1318; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1415 = 7'h47 == total_offset_7[6:0] ? field_byte_7 : _GEN_1319; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1416 = 7'h48 == total_offset_7[6:0] ? field_byte_7 : _GEN_1320; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1417 = 7'h49 == total_offset_7[6:0] ? field_byte_7 : _GEN_1321; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1418 = 7'h4a == total_offset_7[6:0] ? field_byte_7 : _GEN_1322; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1419 = 7'h4b == total_offset_7[6:0] ? field_byte_7 : _GEN_1323; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1420 = 7'h4c == total_offset_7[6:0] ? field_byte_7 : _GEN_1324; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1421 = 7'h4d == total_offset_7[6:0] ? field_byte_7 : _GEN_1325; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1422 = 7'h4e == total_offset_7[6:0] ? field_byte_7 : _GEN_1326; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1423 = 7'h4f == total_offset_7[6:0] ? field_byte_7 : _GEN_1327; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1424 = 7'h50 == total_offset_7[6:0] ? field_byte_7 : _GEN_1328; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1425 = 7'h51 == total_offset_7[6:0] ? field_byte_7 : _GEN_1329; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1426 = 7'h52 == total_offset_7[6:0] ? field_byte_7 : _GEN_1330; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1427 = 7'h53 == total_offset_7[6:0] ? field_byte_7 : _GEN_1331; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1428 = 7'h54 == total_offset_7[6:0] ? field_byte_7 : _GEN_1332; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1429 = 7'h55 == total_offset_7[6:0] ? field_byte_7 : _GEN_1333; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1430 = 7'h56 == total_offset_7[6:0] ? field_byte_7 : _GEN_1334; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1431 = 7'h57 == total_offset_7[6:0] ? field_byte_7 : _GEN_1335; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1432 = 7'h58 == total_offset_7[6:0] ? field_byte_7 : _GEN_1336; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1433 = 7'h59 == total_offset_7[6:0] ? field_byte_7 : _GEN_1337; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1434 = 7'h5a == total_offset_7[6:0] ? field_byte_7 : _GEN_1338; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1435 = 7'h5b == total_offset_7[6:0] ? field_byte_7 : _GEN_1339; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1436 = 7'h5c == total_offset_7[6:0] ? field_byte_7 : _GEN_1340; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1437 = 7'h5d == total_offset_7[6:0] ? field_byte_7 : _GEN_1341; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1438 = 7'h5e == total_offset_7[6:0] ? field_byte_7 : _GEN_1342; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1439 = 7'h5f == total_offset_7[6:0] ? field_byte_7 : _GEN_1343; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1440 = 8'h7 < length_0 ? _GEN_1344 : _GEN_1248; // @[executor.scala 290:56]
  wire [7:0] _GEN_1441 = 8'h7 < length_0 ? _GEN_1345 : _GEN_1249; // @[executor.scala 290:56]
  wire [7:0] _GEN_1442 = 8'h7 < length_0 ? _GEN_1346 : _GEN_1250; // @[executor.scala 290:56]
  wire [7:0] _GEN_1443 = 8'h7 < length_0 ? _GEN_1347 : _GEN_1251; // @[executor.scala 290:56]
  wire [7:0] _GEN_1444 = 8'h7 < length_0 ? _GEN_1348 : _GEN_1252; // @[executor.scala 290:56]
  wire [7:0] _GEN_1445 = 8'h7 < length_0 ? _GEN_1349 : _GEN_1253; // @[executor.scala 290:56]
  wire [7:0] _GEN_1446 = 8'h7 < length_0 ? _GEN_1350 : _GEN_1254; // @[executor.scala 290:56]
  wire [7:0] _GEN_1447 = 8'h7 < length_0 ? _GEN_1351 : _GEN_1255; // @[executor.scala 290:56]
  wire [7:0] _GEN_1448 = 8'h7 < length_0 ? _GEN_1352 : _GEN_1256; // @[executor.scala 290:56]
  wire [7:0] _GEN_1449 = 8'h7 < length_0 ? _GEN_1353 : _GEN_1257; // @[executor.scala 290:56]
  wire [7:0] _GEN_1450 = 8'h7 < length_0 ? _GEN_1354 : _GEN_1258; // @[executor.scala 290:56]
  wire [7:0] _GEN_1451 = 8'h7 < length_0 ? _GEN_1355 : _GEN_1259; // @[executor.scala 290:56]
  wire [7:0] _GEN_1452 = 8'h7 < length_0 ? _GEN_1356 : _GEN_1260; // @[executor.scala 290:56]
  wire [7:0] _GEN_1453 = 8'h7 < length_0 ? _GEN_1357 : _GEN_1261; // @[executor.scala 290:56]
  wire [7:0] _GEN_1454 = 8'h7 < length_0 ? _GEN_1358 : _GEN_1262; // @[executor.scala 290:56]
  wire [7:0] _GEN_1455 = 8'h7 < length_0 ? _GEN_1359 : _GEN_1263; // @[executor.scala 290:56]
  wire [7:0] _GEN_1456 = 8'h7 < length_0 ? _GEN_1360 : _GEN_1264; // @[executor.scala 290:56]
  wire [7:0] _GEN_1457 = 8'h7 < length_0 ? _GEN_1361 : _GEN_1265; // @[executor.scala 290:56]
  wire [7:0] _GEN_1458 = 8'h7 < length_0 ? _GEN_1362 : _GEN_1266; // @[executor.scala 290:56]
  wire [7:0] _GEN_1459 = 8'h7 < length_0 ? _GEN_1363 : _GEN_1267; // @[executor.scala 290:56]
  wire [7:0] _GEN_1460 = 8'h7 < length_0 ? _GEN_1364 : _GEN_1268; // @[executor.scala 290:56]
  wire [7:0] _GEN_1461 = 8'h7 < length_0 ? _GEN_1365 : _GEN_1269; // @[executor.scala 290:56]
  wire [7:0] _GEN_1462 = 8'h7 < length_0 ? _GEN_1366 : _GEN_1270; // @[executor.scala 290:56]
  wire [7:0] _GEN_1463 = 8'h7 < length_0 ? _GEN_1367 : _GEN_1271; // @[executor.scala 290:56]
  wire [7:0] _GEN_1464 = 8'h7 < length_0 ? _GEN_1368 : _GEN_1272; // @[executor.scala 290:56]
  wire [7:0] _GEN_1465 = 8'h7 < length_0 ? _GEN_1369 : _GEN_1273; // @[executor.scala 290:56]
  wire [7:0] _GEN_1466 = 8'h7 < length_0 ? _GEN_1370 : _GEN_1274; // @[executor.scala 290:56]
  wire [7:0] _GEN_1467 = 8'h7 < length_0 ? _GEN_1371 : _GEN_1275; // @[executor.scala 290:56]
  wire [7:0] _GEN_1468 = 8'h7 < length_0 ? _GEN_1372 : _GEN_1276; // @[executor.scala 290:56]
  wire [7:0] _GEN_1469 = 8'h7 < length_0 ? _GEN_1373 : _GEN_1277; // @[executor.scala 290:56]
  wire [7:0] _GEN_1470 = 8'h7 < length_0 ? _GEN_1374 : _GEN_1278; // @[executor.scala 290:56]
  wire [7:0] _GEN_1471 = 8'h7 < length_0 ? _GEN_1375 : _GEN_1279; // @[executor.scala 290:56]
  wire [7:0] _GEN_1472 = 8'h7 < length_0 ? _GEN_1376 : _GEN_1280; // @[executor.scala 290:56]
  wire [7:0] _GEN_1473 = 8'h7 < length_0 ? _GEN_1377 : _GEN_1281; // @[executor.scala 290:56]
  wire [7:0] _GEN_1474 = 8'h7 < length_0 ? _GEN_1378 : _GEN_1282; // @[executor.scala 290:56]
  wire [7:0] _GEN_1475 = 8'h7 < length_0 ? _GEN_1379 : _GEN_1283; // @[executor.scala 290:56]
  wire [7:0] _GEN_1476 = 8'h7 < length_0 ? _GEN_1380 : _GEN_1284; // @[executor.scala 290:56]
  wire [7:0] _GEN_1477 = 8'h7 < length_0 ? _GEN_1381 : _GEN_1285; // @[executor.scala 290:56]
  wire [7:0] _GEN_1478 = 8'h7 < length_0 ? _GEN_1382 : _GEN_1286; // @[executor.scala 290:56]
  wire [7:0] _GEN_1479 = 8'h7 < length_0 ? _GEN_1383 : _GEN_1287; // @[executor.scala 290:56]
  wire [7:0] _GEN_1480 = 8'h7 < length_0 ? _GEN_1384 : _GEN_1288; // @[executor.scala 290:56]
  wire [7:0] _GEN_1481 = 8'h7 < length_0 ? _GEN_1385 : _GEN_1289; // @[executor.scala 290:56]
  wire [7:0] _GEN_1482 = 8'h7 < length_0 ? _GEN_1386 : _GEN_1290; // @[executor.scala 290:56]
  wire [7:0] _GEN_1483 = 8'h7 < length_0 ? _GEN_1387 : _GEN_1291; // @[executor.scala 290:56]
  wire [7:0] _GEN_1484 = 8'h7 < length_0 ? _GEN_1388 : _GEN_1292; // @[executor.scala 290:56]
  wire [7:0] _GEN_1485 = 8'h7 < length_0 ? _GEN_1389 : _GEN_1293; // @[executor.scala 290:56]
  wire [7:0] _GEN_1486 = 8'h7 < length_0 ? _GEN_1390 : _GEN_1294; // @[executor.scala 290:56]
  wire [7:0] _GEN_1487 = 8'h7 < length_0 ? _GEN_1391 : _GEN_1295; // @[executor.scala 290:56]
  wire [7:0] _GEN_1488 = 8'h7 < length_0 ? _GEN_1392 : _GEN_1296; // @[executor.scala 290:56]
  wire [7:0] _GEN_1489 = 8'h7 < length_0 ? _GEN_1393 : _GEN_1297; // @[executor.scala 290:56]
  wire [7:0] _GEN_1490 = 8'h7 < length_0 ? _GEN_1394 : _GEN_1298; // @[executor.scala 290:56]
  wire [7:0] _GEN_1491 = 8'h7 < length_0 ? _GEN_1395 : _GEN_1299; // @[executor.scala 290:56]
  wire [7:0] _GEN_1492 = 8'h7 < length_0 ? _GEN_1396 : _GEN_1300; // @[executor.scala 290:56]
  wire [7:0] _GEN_1493 = 8'h7 < length_0 ? _GEN_1397 : _GEN_1301; // @[executor.scala 290:56]
  wire [7:0] _GEN_1494 = 8'h7 < length_0 ? _GEN_1398 : _GEN_1302; // @[executor.scala 290:56]
  wire [7:0] _GEN_1495 = 8'h7 < length_0 ? _GEN_1399 : _GEN_1303; // @[executor.scala 290:56]
  wire [7:0] _GEN_1496 = 8'h7 < length_0 ? _GEN_1400 : _GEN_1304; // @[executor.scala 290:56]
  wire [7:0] _GEN_1497 = 8'h7 < length_0 ? _GEN_1401 : _GEN_1305; // @[executor.scala 290:56]
  wire [7:0] _GEN_1498 = 8'h7 < length_0 ? _GEN_1402 : _GEN_1306; // @[executor.scala 290:56]
  wire [7:0] _GEN_1499 = 8'h7 < length_0 ? _GEN_1403 : _GEN_1307; // @[executor.scala 290:56]
  wire [7:0] _GEN_1500 = 8'h7 < length_0 ? _GEN_1404 : _GEN_1308; // @[executor.scala 290:56]
  wire [7:0] _GEN_1501 = 8'h7 < length_0 ? _GEN_1405 : _GEN_1309; // @[executor.scala 290:56]
  wire [7:0] _GEN_1502 = 8'h7 < length_0 ? _GEN_1406 : _GEN_1310; // @[executor.scala 290:56]
  wire [7:0] _GEN_1503 = 8'h7 < length_0 ? _GEN_1407 : _GEN_1311; // @[executor.scala 290:56]
  wire [7:0] _GEN_1504 = 8'h7 < length_0 ? _GEN_1408 : _GEN_1312; // @[executor.scala 290:56]
  wire [7:0] _GEN_1505 = 8'h7 < length_0 ? _GEN_1409 : _GEN_1313; // @[executor.scala 290:56]
  wire [7:0] _GEN_1506 = 8'h7 < length_0 ? _GEN_1410 : _GEN_1314; // @[executor.scala 290:56]
  wire [7:0] _GEN_1507 = 8'h7 < length_0 ? _GEN_1411 : _GEN_1315; // @[executor.scala 290:56]
  wire [7:0] _GEN_1508 = 8'h7 < length_0 ? _GEN_1412 : _GEN_1316; // @[executor.scala 290:56]
  wire [7:0] _GEN_1509 = 8'h7 < length_0 ? _GEN_1413 : _GEN_1317; // @[executor.scala 290:56]
  wire [7:0] _GEN_1510 = 8'h7 < length_0 ? _GEN_1414 : _GEN_1318; // @[executor.scala 290:56]
  wire [7:0] _GEN_1511 = 8'h7 < length_0 ? _GEN_1415 : _GEN_1319; // @[executor.scala 290:56]
  wire [7:0] _GEN_1512 = 8'h7 < length_0 ? _GEN_1416 : _GEN_1320; // @[executor.scala 290:56]
  wire [7:0] _GEN_1513 = 8'h7 < length_0 ? _GEN_1417 : _GEN_1321; // @[executor.scala 290:56]
  wire [7:0] _GEN_1514 = 8'h7 < length_0 ? _GEN_1418 : _GEN_1322; // @[executor.scala 290:56]
  wire [7:0] _GEN_1515 = 8'h7 < length_0 ? _GEN_1419 : _GEN_1323; // @[executor.scala 290:56]
  wire [7:0] _GEN_1516 = 8'h7 < length_0 ? _GEN_1420 : _GEN_1324; // @[executor.scala 290:56]
  wire [7:0] _GEN_1517 = 8'h7 < length_0 ? _GEN_1421 : _GEN_1325; // @[executor.scala 290:56]
  wire [7:0] _GEN_1518 = 8'h7 < length_0 ? _GEN_1422 : _GEN_1326; // @[executor.scala 290:56]
  wire [7:0] _GEN_1519 = 8'h7 < length_0 ? _GEN_1423 : _GEN_1327; // @[executor.scala 290:56]
  wire [7:0] _GEN_1520 = 8'h7 < length_0 ? _GEN_1424 : _GEN_1328; // @[executor.scala 290:56]
  wire [7:0] _GEN_1521 = 8'h7 < length_0 ? _GEN_1425 : _GEN_1329; // @[executor.scala 290:56]
  wire [7:0] _GEN_1522 = 8'h7 < length_0 ? _GEN_1426 : _GEN_1330; // @[executor.scala 290:56]
  wire [7:0] _GEN_1523 = 8'h7 < length_0 ? _GEN_1427 : _GEN_1331; // @[executor.scala 290:56]
  wire [7:0] _GEN_1524 = 8'h7 < length_0 ? _GEN_1428 : _GEN_1332; // @[executor.scala 290:56]
  wire [7:0] _GEN_1525 = 8'h7 < length_0 ? _GEN_1429 : _GEN_1333; // @[executor.scala 290:56]
  wire [7:0] _GEN_1526 = 8'h7 < length_0 ? _GEN_1430 : _GEN_1334; // @[executor.scala 290:56]
  wire [7:0] _GEN_1527 = 8'h7 < length_0 ? _GEN_1431 : _GEN_1335; // @[executor.scala 290:56]
  wire [7:0] _GEN_1528 = 8'h7 < length_0 ? _GEN_1432 : _GEN_1336; // @[executor.scala 290:56]
  wire [7:0] _GEN_1529 = 8'h7 < length_0 ? _GEN_1433 : _GEN_1337; // @[executor.scala 290:56]
  wire [7:0] _GEN_1530 = 8'h7 < length_0 ? _GEN_1434 : _GEN_1338; // @[executor.scala 290:56]
  wire [7:0] _GEN_1531 = 8'h7 < length_0 ? _GEN_1435 : _GEN_1339; // @[executor.scala 290:56]
  wire [7:0] _GEN_1532 = 8'h7 < length_0 ? _GEN_1436 : _GEN_1340; // @[executor.scala 290:56]
  wire [7:0] _GEN_1533 = 8'h7 < length_0 ? _GEN_1437 : _GEN_1341; // @[executor.scala 290:56]
  wire [7:0] _GEN_1534 = 8'h7 < length_0 ? _GEN_1438 : _GEN_1342; // @[executor.scala 290:56]
  wire [7:0] _GEN_1535 = 8'h7 < length_0 ? _GEN_1439 : _GEN_1343; // @[executor.scala 290:56]
  wire [63:0] _GEN_1536 = length_0 == 8'h0 ? field_0 : {{62'd0}, phv_next_processor_id}; // @[executor.scala 283:67 executor.scala 284:51 executor.scala 270:25]
  wire [7:0] _GEN_1537 = length_0 == 8'h0 ? phv_data_0 : _GEN_1440; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1538 = length_0 == 8'h0 ? phv_data_1 : _GEN_1441; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1539 = length_0 == 8'h0 ? phv_data_2 : _GEN_1442; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1540 = length_0 == 8'h0 ? phv_data_3 : _GEN_1443; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1541 = length_0 == 8'h0 ? phv_data_4 : _GEN_1444; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1542 = length_0 == 8'h0 ? phv_data_5 : _GEN_1445; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1543 = length_0 == 8'h0 ? phv_data_6 : _GEN_1446; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1544 = length_0 == 8'h0 ? phv_data_7 : _GEN_1447; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1545 = length_0 == 8'h0 ? phv_data_8 : _GEN_1448; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1546 = length_0 == 8'h0 ? phv_data_9 : _GEN_1449; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1547 = length_0 == 8'h0 ? phv_data_10 : _GEN_1450; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1548 = length_0 == 8'h0 ? phv_data_11 : _GEN_1451; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1549 = length_0 == 8'h0 ? phv_data_12 : _GEN_1452; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1550 = length_0 == 8'h0 ? phv_data_13 : _GEN_1453; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1551 = length_0 == 8'h0 ? phv_data_14 : _GEN_1454; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1552 = length_0 == 8'h0 ? phv_data_15 : _GEN_1455; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1553 = length_0 == 8'h0 ? phv_data_16 : _GEN_1456; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1554 = length_0 == 8'h0 ? phv_data_17 : _GEN_1457; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1555 = length_0 == 8'h0 ? phv_data_18 : _GEN_1458; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1556 = length_0 == 8'h0 ? phv_data_19 : _GEN_1459; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1557 = length_0 == 8'h0 ? phv_data_20 : _GEN_1460; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1558 = length_0 == 8'h0 ? phv_data_21 : _GEN_1461; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1559 = length_0 == 8'h0 ? phv_data_22 : _GEN_1462; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1560 = length_0 == 8'h0 ? phv_data_23 : _GEN_1463; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1561 = length_0 == 8'h0 ? phv_data_24 : _GEN_1464; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1562 = length_0 == 8'h0 ? phv_data_25 : _GEN_1465; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1563 = length_0 == 8'h0 ? phv_data_26 : _GEN_1466; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1564 = length_0 == 8'h0 ? phv_data_27 : _GEN_1467; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1565 = length_0 == 8'h0 ? phv_data_28 : _GEN_1468; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1566 = length_0 == 8'h0 ? phv_data_29 : _GEN_1469; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1567 = length_0 == 8'h0 ? phv_data_30 : _GEN_1470; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1568 = length_0 == 8'h0 ? phv_data_31 : _GEN_1471; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1569 = length_0 == 8'h0 ? phv_data_32 : _GEN_1472; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1570 = length_0 == 8'h0 ? phv_data_33 : _GEN_1473; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1571 = length_0 == 8'h0 ? phv_data_34 : _GEN_1474; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1572 = length_0 == 8'h0 ? phv_data_35 : _GEN_1475; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1573 = length_0 == 8'h0 ? phv_data_36 : _GEN_1476; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1574 = length_0 == 8'h0 ? phv_data_37 : _GEN_1477; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1575 = length_0 == 8'h0 ? phv_data_38 : _GEN_1478; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1576 = length_0 == 8'h0 ? phv_data_39 : _GEN_1479; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1577 = length_0 == 8'h0 ? phv_data_40 : _GEN_1480; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1578 = length_0 == 8'h0 ? phv_data_41 : _GEN_1481; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1579 = length_0 == 8'h0 ? phv_data_42 : _GEN_1482; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1580 = length_0 == 8'h0 ? phv_data_43 : _GEN_1483; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1581 = length_0 == 8'h0 ? phv_data_44 : _GEN_1484; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1582 = length_0 == 8'h0 ? phv_data_45 : _GEN_1485; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1583 = length_0 == 8'h0 ? phv_data_46 : _GEN_1486; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1584 = length_0 == 8'h0 ? phv_data_47 : _GEN_1487; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1585 = length_0 == 8'h0 ? phv_data_48 : _GEN_1488; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1586 = length_0 == 8'h0 ? phv_data_49 : _GEN_1489; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1587 = length_0 == 8'h0 ? phv_data_50 : _GEN_1490; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1588 = length_0 == 8'h0 ? phv_data_51 : _GEN_1491; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1589 = length_0 == 8'h0 ? phv_data_52 : _GEN_1492; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1590 = length_0 == 8'h0 ? phv_data_53 : _GEN_1493; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1591 = length_0 == 8'h0 ? phv_data_54 : _GEN_1494; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1592 = length_0 == 8'h0 ? phv_data_55 : _GEN_1495; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1593 = length_0 == 8'h0 ? phv_data_56 : _GEN_1496; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1594 = length_0 == 8'h0 ? phv_data_57 : _GEN_1497; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1595 = length_0 == 8'h0 ? phv_data_58 : _GEN_1498; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1596 = length_0 == 8'h0 ? phv_data_59 : _GEN_1499; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1597 = length_0 == 8'h0 ? phv_data_60 : _GEN_1500; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1598 = length_0 == 8'h0 ? phv_data_61 : _GEN_1501; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1599 = length_0 == 8'h0 ? phv_data_62 : _GEN_1502; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1600 = length_0 == 8'h0 ? phv_data_63 : _GEN_1503; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1601 = length_0 == 8'h0 ? phv_data_64 : _GEN_1504; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1602 = length_0 == 8'h0 ? phv_data_65 : _GEN_1505; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1603 = length_0 == 8'h0 ? phv_data_66 : _GEN_1506; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1604 = length_0 == 8'h0 ? phv_data_67 : _GEN_1507; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1605 = length_0 == 8'h0 ? phv_data_68 : _GEN_1508; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1606 = length_0 == 8'h0 ? phv_data_69 : _GEN_1509; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1607 = length_0 == 8'h0 ? phv_data_70 : _GEN_1510; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1608 = length_0 == 8'h0 ? phv_data_71 : _GEN_1511; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1609 = length_0 == 8'h0 ? phv_data_72 : _GEN_1512; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1610 = length_0 == 8'h0 ? phv_data_73 : _GEN_1513; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1611 = length_0 == 8'h0 ? phv_data_74 : _GEN_1514; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1612 = length_0 == 8'h0 ? phv_data_75 : _GEN_1515; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1613 = length_0 == 8'h0 ? phv_data_76 : _GEN_1516; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1614 = length_0 == 8'h0 ? phv_data_77 : _GEN_1517; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1615 = length_0 == 8'h0 ? phv_data_78 : _GEN_1518; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1616 = length_0 == 8'h0 ? phv_data_79 : _GEN_1519; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1617 = length_0 == 8'h0 ? phv_data_80 : _GEN_1520; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1618 = length_0 == 8'h0 ? phv_data_81 : _GEN_1521; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1619 = length_0 == 8'h0 ? phv_data_82 : _GEN_1522; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1620 = length_0 == 8'h0 ? phv_data_83 : _GEN_1523; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1621 = length_0 == 8'h0 ? phv_data_84 : _GEN_1524; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1622 = length_0 == 8'h0 ? phv_data_85 : _GEN_1525; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1623 = length_0 == 8'h0 ? phv_data_86 : _GEN_1526; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1624 = length_0 == 8'h0 ? phv_data_87 : _GEN_1527; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1625 = length_0 == 8'h0 ? phv_data_88 : _GEN_1528; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1626 = length_0 == 8'h0 ? phv_data_89 : _GEN_1529; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1627 = length_0 == 8'h0 ? phv_data_90 : _GEN_1530; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1628 = length_0 == 8'h0 ? phv_data_91 : _GEN_1531; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1629 = length_0 == 8'h0 ? phv_data_92 : _GEN_1532; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1630 = length_0 == 8'h0 ? phv_data_93 : _GEN_1533; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1631 = length_0 == 8'h0 ? phv_data_94 : _GEN_1534; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] _GEN_1632 = length_0 == 8'h0 ? phv_data_95 : _GEN_1535; // @[executor.scala 283:67 executor.scala 270:25]
  wire [7:0] field_byte_8 = field_1[63:56]; // @[executor.scala 287:53]
  wire [8:0] _total_offset_T_8 = {{1'd0}, offset_1}; // @[executor.scala 289:53]
  wire [7:0] total_offset_8 = _total_offset_T_8[7:0]; // @[executor.scala 289:53]
  wire [7:0] _GEN_1633 = 7'h0 == total_offset_8[6:0] ? field_byte_8 : _GEN_1537; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1634 = 7'h1 == total_offset_8[6:0] ? field_byte_8 : _GEN_1538; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1635 = 7'h2 == total_offset_8[6:0] ? field_byte_8 : _GEN_1539; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1636 = 7'h3 == total_offset_8[6:0] ? field_byte_8 : _GEN_1540; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1637 = 7'h4 == total_offset_8[6:0] ? field_byte_8 : _GEN_1541; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1638 = 7'h5 == total_offset_8[6:0] ? field_byte_8 : _GEN_1542; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1639 = 7'h6 == total_offset_8[6:0] ? field_byte_8 : _GEN_1543; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1640 = 7'h7 == total_offset_8[6:0] ? field_byte_8 : _GEN_1544; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1641 = 7'h8 == total_offset_8[6:0] ? field_byte_8 : _GEN_1545; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1642 = 7'h9 == total_offset_8[6:0] ? field_byte_8 : _GEN_1546; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1643 = 7'ha == total_offset_8[6:0] ? field_byte_8 : _GEN_1547; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1644 = 7'hb == total_offset_8[6:0] ? field_byte_8 : _GEN_1548; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1645 = 7'hc == total_offset_8[6:0] ? field_byte_8 : _GEN_1549; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1646 = 7'hd == total_offset_8[6:0] ? field_byte_8 : _GEN_1550; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1647 = 7'he == total_offset_8[6:0] ? field_byte_8 : _GEN_1551; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1648 = 7'hf == total_offset_8[6:0] ? field_byte_8 : _GEN_1552; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1649 = 7'h10 == total_offset_8[6:0] ? field_byte_8 : _GEN_1553; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1650 = 7'h11 == total_offset_8[6:0] ? field_byte_8 : _GEN_1554; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1651 = 7'h12 == total_offset_8[6:0] ? field_byte_8 : _GEN_1555; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1652 = 7'h13 == total_offset_8[6:0] ? field_byte_8 : _GEN_1556; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1653 = 7'h14 == total_offset_8[6:0] ? field_byte_8 : _GEN_1557; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1654 = 7'h15 == total_offset_8[6:0] ? field_byte_8 : _GEN_1558; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1655 = 7'h16 == total_offset_8[6:0] ? field_byte_8 : _GEN_1559; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1656 = 7'h17 == total_offset_8[6:0] ? field_byte_8 : _GEN_1560; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1657 = 7'h18 == total_offset_8[6:0] ? field_byte_8 : _GEN_1561; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1658 = 7'h19 == total_offset_8[6:0] ? field_byte_8 : _GEN_1562; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1659 = 7'h1a == total_offset_8[6:0] ? field_byte_8 : _GEN_1563; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1660 = 7'h1b == total_offset_8[6:0] ? field_byte_8 : _GEN_1564; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1661 = 7'h1c == total_offset_8[6:0] ? field_byte_8 : _GEN_1565; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1662 = 7'h1d == total_offset_8[6:0] ? field_byte_8 : _GEN_1566; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1663 = 7'h1e == total_offset_8[6:0] ? field_byte_8 : _GEN_1567; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1664 = 7'h1f == total_offset_8[6:0] ? field_byte_8 : _GEN_1568; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1665 = 7'h20 == total_offset_8[6:0] ? field_byte_8 : _GEN_1569; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1666 = 7'h21 == total_offset_8[6:0] ? field_byte_8 : _GEN_1570; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1667 = 7'h22 == total_offset_8[6:0] ? field_byte_8 : _GEN_1571; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1668 = 7'h23 == total_offset_8[6:0] ? field_byte_8 : _GEN_1572; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1669 = 7'h24 == total_offset_8[6:0] ? field_byte_8 : _GEN_1573; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1670 = 7'h25 == total_offset_8[6:0] ? field_byte_8 : _GEN_1574; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1671 = 7'h26 == total_offset_8[6:0] ? field_byte_8 : _GEN_1575; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1672 = 7'h27 == total_offset_8[6:0] ? field_byte_8 : _GEN_1576; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1673 = 7'h28 == total_offset_8[6:0] ? field_byte_8 : _GEN_1577; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1674 = 7'h29 == total_offset_8[6:0] ? field_byte_8 : _GEN_1578; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1675 = 7'h2a == total_offset_8[6:0] ? field_byte_8 : _GEN_1579; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1676 = 7'h2b == total_offset_8[6:0] ? field_byte_8 : _GEN_1580; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1677 = 7'h2c == total_offset_8[6:0] ? field_byte_8 : _GEN_1581; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1678 = 7'h2d == total_offset_8[6:0] ? field_byte_8 : _GEN_1582; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1679 = 7'h2e == total_offset_8[6:0] ? field_byte_8 : _GEN_1583; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1680 = 7'h2f == total_offset_8[6:0] ? field_byte_8 : _GEN_1584; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1681 = 7'h30 == total_offset_8[6:0] ? field_byte_8 : _GEN_1585; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1682 = 7'h31 == total_offset_8[6:0] ? field_byte_8 : _GEN_1586; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1683 = 7'h32 == total_offset_8[6:0] ? field_byte_8 : _GEN_1587; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1684 = 7'h33 == total_offset_8[6:0] ? field_byte_8 : _GEN_1588; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1685 = 7'h34 == total_offset_8[6:0] ? field_byte_8 : _GEN_1589; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1686 = 7'h35 == total_offset_8[6:0] ? field_byte_8 : _GEN_1590; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1687 = 7'h36 == total_offset_8[6:0] ? field_byte_8 : _GEN_1591; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1688 = 7'h37 == total_offset_8[6:0] ? field_byte_8 : _GEN_1592; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1689 = 7'h38 == total_offset_8[6:0] ? field_byte_8 : _GEN_1593; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1690 = 7'h39 == total_offset_8[6:0] ? field_byte_8 : _GEN_1594; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1691 = 7'h3a == total_offset_8[6:0] ? field_byte_8 : _GEN_1595; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1692 = 7'h3b == total_offset_8[6:0] ? field_byte_8 : _GEN_1596; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1693 = 7'h3c == total_offset_8[6:0] ? field_byte_8 : _GEN_1597; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1694 = 7'h3d == total_offset_8[6:0] ? field_byte_8 : _GEN_1598; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1695 = 7'h3e == total_offset_8[6:0] ? field_byte_8 : _GEN_1599; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1696 = 7'h3f == total_offset_8[6:0] ? field_byte_8 : _GEN_1600; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1697 = 7'h40 == total_offset_8[6:0] ? field_byte_8 : _GEN_1601; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1698 = 7'h41 == total_offset_8[6:0] ? field_byte_8 : _GEN_1602; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1699 = 7'h42 == total_offset_8[6:0] ? field_byte_8 : _GEN_1603; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1700 = 7'h43 == total_offset_8[6:0] ? field_byte_8 : _GEN_1604; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1701 = 7'h44 == total_offset_8[6:0] ? field_byte_8 : _GEN_1605; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1702 = 7'h45 == total_offset_8[6:0] ? field_byte_8 : _GEN_1606; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1703 = 7'h46 == total_offset_8[6:0] ? field_byte_8 : _GEN_1607; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1704 = 7'h47 == total_offset_8[6:0] ? field_byte_8 : _GEN_1608; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1705 = 7'h48 == total_offset_8[6:0] ? field_byte_8 : _GEN_1609; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1706 = 7'h49 == total_offset_8[6:0] ? field_byte_8 : _GEN_1610; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1707 = 7'h4a == total_offset_8[6:0] ? field_byte_8 : _GEN_1611; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1708 = 7'h4b == total_offset_8[6:0] ? field_byte_8 : _GEN_1612; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1709 = 7'h4c == total_offset_8[6:0] ? field_byte_8 : _GEN_1613; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1710 = 7'h4d == total_offset_8[6:0] ? field_byte_8 : _GEN_1614; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1711 = 7'h4e == total_offset_8[6:0] ? field_byte_8 : _GEN_1615; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1712 = 7'h4f == total_offset_8[6:0] ? field_byte_8 : _GEN_1616; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1713 = 7'h50 == total_offset_8[6:0] ? field_byte_8 : _GEN_1617; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1714 = 7'h51 == total_offset_8[6:0] ? field_byte_8 : _GEN_1618; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1715 = 7'h52 == total_offset_8[6:0] ? field_byte_8 : _GEN_1619; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1716 = 7'h53 == total_offset_8[6:0] ? field_byte_8 : _GEN_1620; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1717 = 7'h54 == total_offset_8[6:0] ? field_byte_8 : _GEN_1621; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1718 = 7'h55 == total_offset_8[6:0] ? field_byte_8 : _GEN_1622; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1719 = 7'h56 == total_offset_8[6:0] ? field_byte_8 : _GEN_1623; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1720 = 7'h57 == total_offset_8[6:0] ? field_byte_8 : _GEN_1624; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1721 = 7'h58 == total_offset_8[6:0] ? field_byte_8 : _GEN_1625; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1722 = 7'h59 == total_offset_8[6:0] ? field_byte_8 : _GEN_1626; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1723 = 7'h5a == total_offset_8[6:0] ? field_byte_8 : _GEN_1627; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1724 = 7'h5b == total_offset_8[6:0] ? field_byte_8 : _GEN_1628; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1725 = 7'h5c == total_offset_8[6:0] ? field_byte_8 : _GEN_1629; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1726 = 7'h5d == total_offset_8[6:0] ? field_byte_8 : _GEN_1630; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1727 = 7'h5e == total_offset_8[6:0] ? field_byte_8 : _GEN_1631; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1728 = 7'h5f == total_offset_8[6:0] ? field_byte_8 : _GEN_1632; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1729 = 8'h0 < length_1 ? _GEN_1633 : _GEN_1537; // @[executor.scala 290:56]
  wire [7:0] _GEN_1730 = 8'h0 < length_1 ? _GEN_1634 : _GEN_1538; // @[executor.scala 290:56]
  wire [7:0] _GEN_1731 = 8'h0 < length_1 ? _GEN_1635 : _GEN_1539; // @[executor.scala 290:56]
  wire [7:0] _GEN_1732 = 8'h0 < length_1 ? _GEN_1636 : _GEN_1540; // @[executor.scala 290:56]
  wire [7:0] _GEN_1733 = 8'h0 < length_1 ? _GEN_1637 : _GEN_1541; // @[executor.scala 290:56]
  wire [7:0] _GEN_1734 = 8'h0 < length_1 ? _GEN_1638 : _GEN_1542; // @[executor.scala 290:56]
  wire [7:0] _GEN_1735 = 8'h0 < length_1 ? _GEN_1639 : _GEN_1543; // @[executor.scala 290:56]
  wire [7:0] _GEN_1736 = 8'h0 < length_1 ? _GEN_1640 : _GEN_1544; // @[executor.scala 290:56]
  wire [7:0] _GEN_1737 = 8'h0 < length_1 ? _GEN_1641 : _GEN_1545; // @[executor.scala 290:56]
  wire [7:0] _GEN_1738 = 8'h0 < length_1 ? _GEN_1642 : _GEN_1546; // @[executor.scala 290:56]
  wire [7:0] _GEN_1739 = 8'h0 < length_1 ? _GEN_1643 : _GEN_1547; // @[executor.scala 290:56]
  wire [7:0] _GEN_1740 = 8'h0 < length_1 ? _GEN_1644 : _GEN_1548; // @[executor.scala 290:56]
  wire [7:0] _GEN_1741 = 8'h0 < length_1 ? _GEN_1645 : _GEN_1549; // @[executor.scala 290:56]
  wire [7:0] _GEN_1742 = 8'h0 < length_1 ? _GEN_1646 : _GEN_1550; // @[executor.scala 290:56]
  wire [7:0] _GEN_1743 = 8'h0 < length_1 ? _GEN_1647 : _GEN_1551; // @[executor.scala 290:56]
  wire [7:0] _GEN_1744 = 8'h0 < length_1 ? _GEN_1648 : _GEN_1552; // @[executor.scala 290:56]
  wire [7:0] _GEN_1745 = 8'h0 < length_1 ? _GEN_1649 : _GEN_1553; // @[executor.scala 290:56]
  wire [7:0] _GEN_1746 = 8'h0 < length_1 ? _GEN_1650 : _GEN_1554; // @[executor.scala 290:56]
  wire [7:0] _GEN_1747 = 8'h0 < length_1 ? _GEN_1651 : _GEN_1555; // @[executor.scala 290:56]
  wire [7:0] _GEN_1748 = 8'h0 < length_1 ? _GEN_1652 : _GEN_1556; // @[executor.scala 290:56]
  wire [7:0] _GEN_1749 = 8'h0 < length_1 ? _GEN_1653 : _GEN_1557; // @[executor.scala 290:56]
  wire [7:0] _GEN_1750 = 8'h0 < length_1 ? _GEN_1654 : _GEN_1558; // @[executor.scala 290:56]
  wire [7:0] _GEN_1751 = 8'h0 < length_1 ? _GEN_1655 : _GEN_1559; // @[executor.scala 290:56]
  wire [7:0] _GEN_1752 = 8'h0 < length_1 ? _GEN_1656 : _GEN_1560; // @[executor.scala 290:56]
  wire [7:0] _GEN_1753 = 8'h0 < length_1 ? _GEN_1657 : _GEN_1561; // @[executor.scala 290:56]
  wire [7:0] _GEN_1754 = 8'h0 < length_1 ? _GEN_1658 : _GEN_1562; // @[executor.scala 290:56]
  wire [7:0] _GEN_1755 = 8'h0 < length_1 ? _GEN_1659 : _GEN_1563; // @[executor.scala 290:56]
  wire [7:0] _GEN_1756 = 8'h0 < length_1 ? _GEN_1660 : _GEN_1564; // @[executor.scala 290:56]
  wire [7:0] _GEN_1757 = 8'h0 < length_1 ? _GEN_1661 : _GEN_1565; // @[executor.scala 290:56]
  wire [7:0] _GEN_1758 = 8'h0 < length_1 ? _GEN_1662 : _GEN_1566; // @[executor.scala 290:56]
  wire [7:0] _GEN_1759 = 8'h0 < length_1 ? _GEN_1663 : _GEN_1567; // @[executor.scala 290:56]
  wire [7:0] _GEN_1760 = 8'h0 < length_1 ? _GEN_1664 : _GEN_1568; // @[executor.scala 290:56]
  wire [7:0] _GEN_1761 = 8'h0 < length_1 ? _GEN_1665 : _GEN_1569; // @[executor.scala 290:56]
  wire [7:0] _GEN_1762 = 8'h0 < length_1 ? _GEN_1666 : _GEN_1570; // @[executor.scala 290:56]
  wire [7:0] _GEN_1763 = 8'h0 < length_1 ? _GEN_1667 : _GEN_1571; // @[executor.scala 290:56]
  wire [7:0] _GEN_1764 = 8'h0 < length_1 ? _GEN_1668 : _GEN_1572; // @[executor.scala 290:56]
  wire [7:0] _GEN_1765 = 8'h0 < length_1 ? _GEN_1669 : _GEN_1573; // @[executor.scala 290:56]
  wire [7:0] _GEN_1766 = 8'h0 < length_1 ? _GEN_1670 : _GEN_1574; // @[executor.scala 290:56]
  wire [7:0] _GEN_1767 = 8'h0 < length_1 ? _GEN_1671 : _GEN_1575; // @[executor.scala 290:56]
  wire [7:0] _GEN_1768 = 8'h0 < length_1 ? _GEN_1672 : _GEN_1576; // @[executor.scala 290:56]
  wire [7:0] _GEN_1769 = 8'h0 < length_1 ? _GEN_1673 : _GEN_1577; // @[executor.scala 290:56]
  wire [7:0] _GEN_1770 = 8'h0 < length_1 ? _GEN_1674 : _GEN_1578; // @[executor.scala 290:56]
  wire [7:0] _GEN_1771 = 8'h0 < length_1 ? _GEN_1675 : _GEN_1579; // @[executor.scala 290:56]
  wire [7:0] _GEN_1772 = 8'h0 < length_1 ? _GEN_1676 : _GEN_1580; // @[executor.scala 290:56]
  wire [7:0] _GEN_1773 = 8'h0 < length_1 ? _GEN_1677 : _GEN_1581; // @[executor.scala 290:56]
  wire [7:0] _GEN_1774 = 8'h0 < length_1 ? _GEN_1678 : _GEN_1582; // @[executor.scala 290:56]
  wire [7:0] _GEN_1775 = 8'h0 < length_1 ? _GEN_1679 : _GEN_1583; // @[executor.scala 290:56]
  wire [7:0] _GEN_1776 = 8'h0 < length_1 ? _GEN_1680 : _GEN_1584; // @[executor.scala 290:56]
  wire [7:0] _GEN_1777 = 8'h0 < length_1 ? _GEN_1681 : _GEN_1585; // @[executor.scala 290:56]
  wire [7:0] _GEN_1778 = 8'h0 < length_1 ? _GEN_1682 : _GEN_1586; // @[executor.scala 290:56]
  wire [7:0] _GEN_1779 = 8'h0 < length_1 ? _GEN_1683 : _GEN_1587; // @[executor.scala 290:56]
  wire [7:0] _GEN_1780 = 8'h0 < length_1 ? _GEN_1684 : _GEN_1588; // @[executor.scala 290:56]
  wire [7:0] _GEN_1781 = 8'h0 < length_1 ? _GEN_1685 : _GEN_1589; // @[executor.scala 290:56]
  wire [7:0] _GEN_1782 = 8'h0 < length_1 ? _GEN_1686 : _GEN_1590; // @[executor.scala 290:56]
  wire [7:0] _GEN_1783 = 8'h0 < length_1 ? _GEN_1687 : _GEN_1591; // @[executor.scala 290:56]
  wire [7:0] _GEN_1784 = 8'h0 < length_1 ? _GEN_1688 : _GEN_1592; // @[executor.scala 290:56]
  wire [7:0] _GEN_1785 = 8'h0 < length_1 ? _GEN_1689 : _GEN_1593; // @[executor.scala 290:56]
  wire [7:0] _GEN_1786 = 8'h0 < length_1 ? _GEN_1690 : _GEN_1594; // @[executor.scala 290:56]
  wire [7:0] _GEN_1787 = 8'h0 < length_1 ? _GEN_1691 : _GEN_1595; // @[executor.scala 290:56]
  wire [7:0] _GEN_1788 = 8'h0 < length_1 ? _GEN_1692 : _GEN_1596; // @[executor.scala 290:56]
  wire [7:0] _GEN_1789 = 8'h0 < length_1 ? _GEN_1693 : _GEN_1597; // @[executor.scala 290:56]
  wire [7:0] _GEN_1790 = 8'h0 < length_1 ? _GEN_1694 : _GEN_1598; // @[executor.scala 290:56]
  wire [7:0] _GEN_1791 = 8'h0 < length_1 ? _GEN_1695 : _GEN_1599; // @[executor.scala 290:56]
  wire [7:0] _GEN_1792 = 8'h0 < length_1 ? _GEN_1696 : _GEN_1600; // @[executor.scala 290:56]
  wire [7:0] _GEN_1793 = 8'h0 < length_1 ? _GEN_1697 : _GEN_1601; // @[executor.scala 290:56]
  wire [7:0] _GEN_1794 = 8'h0 < length_1 ? _GEN_1698 : _GEN_1602; // @[executor.scala 290:56]
  wire [7:0] _GEN_1795 = 8'h0 < length_1 ? _GEN_1699 : _GEN_1603; // @[executor.scala 290:56]
  wire [7:0] _GEN_1796 = 8'h0 < length_1 ? _GEN_1700 : _GEN_1604; // @[executor.scala 290:56]
  wire [7:0] _GEN_1797 = 8'h0 < length_1 ? _GEN_1701 : _GEN_1605; // @[executor.scala 290:56]
  wire [7:0] _GEN_1798 = 8'h0 < length_1 ? _GEN_1702 : _GEN_1606; // @[executor.scala 290:56]
  wire [7:0] _GEN_1799 = 8'h0 < length_1 ? _GEN_1703 : _GEN_1607; // @[executor.scala 290:56]
  wire [7:0] _GEN_1800 = 8'h0 < length_1 ? _GEN_1704 : _GEN_1608; // @[executor.scala 290:56]
  wire [7:0] _GEN_1801 = 8'h0 < length_1 ? _GEN_1705 : _GEN_1609; // @[executor.scala 290:56]
  wire [7:0] _GEN_1802 = 8'h0 < length_1 ? _GEN_1706 : _GEN_1610; // @[executor.scala 290:56]
  wire [7:0] _GEN_1803 = 8'h0 < length_1 ? _GEN_1707 : _GEN_1611; // @[executor.scala 290:56]
  wire [7:0] _GEN_1804 = 8'h0 < length_1 ? _GEN_1708 : _GEN_1612; // @[executor.scala 290:56]
  wire [7:0] _GEN_1805 = 8'h0 < length_1 ? _GEN_1709 : _GEN_1613; // @[executor.scala 290:56]
  wire [7:0] _GEN_1806 = 8'h0 < length_1 ? _GEN_1710 : _GEN_1614; // @[executor.scala 290:56]
  wire [7:0] _GEN_1807 = 8'h0 < length_1 ? _GEN_1711 : _GEN_1615; // @[executor.scala 290:56]
  wire [7:0] _GEN_1808 = 8'h0 < length_1 ? _GEN_1712 : _GEN_1616; // @[executor.scala 290:56]
  wire [7:0] _GEN_1809 = 8'h0 < length_1 ? _GEN_1713 : _GEN_1617; // @[executor.scala 290:56]
  wire [7:0] _GEN_1810 = 8'h0 < length_1 ? _GEN_1714 : _GEN_1618; // @[executor.scala 290:56]
  wire [7:0] _GEN_1811 = 8'h0 < length_1 ? _GEN_1715 : _GEN_1619; // @[executor.scala 290:56]
  wire [7:0] _GEN_1812 = 8'h0 < length_1 ? _GEN_1716 : _GEN_1620; // @[executor.scala 290:56]
  wire [7:0] _GEN_1813 = 8'h0 < length_1 ? _GEN_1717 : _GEN_1621; // @[executor.scala 290:56]
  wire [7:0] _GEN_1814 = 8'h0 < length_1 ? _GEN_1718 : _GEN_1622; // @[executor.scala 290:56]
  wire [7:0] _GEN_1815 = 8'h0 < length_1 ? _GEN_1719 : _GEN_1623; // @[executor.scala 290:56]
  wire [7:0] _GEN_1816 = 8'h0 < length_1 ? _GEN_1720 : _GEN_1624; // @[executor.scala 290:56]
  wire [7:0] _GEN_1817 = 8'h0 < length_1 ? _GEN_1721 : _GEN_1625; // @[executor.scala 290:56]
  wire [7:0] _GEN_1818 = 8'h0 < length_1 ? _GEN_1722 : _GEN_1626; // @[executor.scala 290:56]
  wire [7:0] _GEN_1819 = 8'h0 < length_1 ? _GEN_1723 : _GEN_1627; // @[executor.scala 290:56]
  wire [7:0] _GEN_1820 = 8'h0 < length_1 ? _GEN_1724 : _GEN_1628; // @[executor.scala 290:56]
  wire [7:0] _GEN_1821 = 8'h0 < length_1 ? _GEN_1725 : _GEN_1629; // @[executor.scala 290:56]
  wire [7:0] _GEN_1822 = 8'h0 < length_1 ? _GEN_1726 : _GEN_1630; // @[executor.scala 290:56]
  wire [7:0] _GEN_1823 = 8'h0 < length_1 ? _GEN_1727 : _GEN_1631; // @[executor.scala 290:56]
  wire [7:0] _GEN_1824 = 8'h0 < length_1 ? _GEN_1728 : _GEN_1632; // @[executor.scala 290:56]
  wire [7:0] field_byte_9 = field_1[55:48]; // @[executor.scala 287:53]
  wire [7:0] total_offset_9 = offset_1 + 8'h1; // @[executor.scala 289:53]
  wire [7:0] _GEN_1825 = 7'h0 == total_offset_9[6:0] ? field_byte_9 : _GEN_1729; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1826 = 7'h1 == total_offset_9[6:0] ? field_byte_9 : _GEN_1730; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1827 = 7'h2 == total_offset_9[6:0] ? field_byte_9 : _GEN_1731; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1828 = 7'h3 == total_offset_9[6:0] ? field_byte_9 : _GEN_1732; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1829 = 7'h4 == total_offset_9[6:0] ? field_byte_9 : _GEN_1733; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1830 = 7'h5 == total_offset_9[6:0] ? field_byte_9 : _GEN_1734; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1831 = 7'h6 == total_offset_9[6:0] ? field_byte_9 : _GEN_1735; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1832 = 7'h7 == total_offset_9[6:0] ? field_byte_9 : _GEN_1736; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1833 = 7'h8 == total_offset_9[6:0] ? field_byte_9 : _GEN_1737; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1834 = 7'h9 == total_offset_9[6:0] ? field_byte_9 : _GEN_1738; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1835 = 7'ha == total_offset_9[6:0] ? field_byte_9 : _GEN_1739; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1836 = 7'hb == total_offset_9[6:0] ? field_byte_9 : _GEN_1740; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1837 = 7'hc == total_offset_9[6:0] ? field_byte_9 : _GEN_1741; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1838 = 7'hd == total_offset_9[6:0] ? field_byte_9 : _GEN_1742; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1839 = 7'he == total_offset_9[6:0] ? field_byte_9 : _GEN_1743; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1840 = 7'hf == total_offset_9[6:0] ? field_byte_9 : _GEN_1744; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1841 = 7'h10 == total_offset_9[6:0] ? field_byte_9 : _GEN_1745; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1842 = 7'h11 == total_offset_9[6:0] ? field_byte_9 : _GEN_1746; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1843 = 7'h12 == total_offset_9[6:0] ? field_byte_9 : _GEN_1747; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1844 = 7'h13 == total_offset_9[6:0] ? field_byte_9 : _GEN_1748; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1845 = 7'h14 == total_offset_9[6:0] ? field_byte_9 : _GEN_1749; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1846 = 7'h15 == total_offset_9[6:0] ? field_byte_9 : _GEN_1750; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1847 = 7'h16 == total_offset_9[6:0] ? field_byte_9 : _GEN_1751; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1848 = 7'h17 == total_offset_9[6:0] ? field_byte_9 : _GEN_1752; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1849 = 7'h18 == total_offset_9[6:0] ? field_byte_9 : _GEN_1753; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1850 = 7'h19 == total_offset_9[6:0] ? field_byte_9 : _GEN_1754; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1851 = 7'h1a == total_offset_9[6:0] ? field_byte_9 : _GEN_1755; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1852 = 7'h1b == total_offset_9[6:0] ? field_byte_9 : _GEN_1756; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1853 = 7'h1c == total_offset_9[6:0] ? field_byte_9 : _GEN_1757; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1854 = 7'h1d == total_offset_9[6:0] ? field_byte_9 : _GEN_1758; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1855 = 7'h1e == total_offset_9[6:0] ? field_byte_9 : _GEN_1759; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1856 = 7'h1f == total_offset_9[6:0] ? field_byte_9 : _GEN_1760; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1857 = 7'h20 == total_offset_9[6:0] ? field_byte_9 : _GEN_1761; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1858 = 7'h21 == total_offset_9[6:0] ? field_byte_9 : _GEN_1762; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1859 = 7'h22 == total_offset_9[6:0] ? field_byte_9 : _GEN_1763; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1860 = 7'h23 == total_offset_9[6:0] ? field_byte_9 : _GEN_1764; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1861 = 7'h24 == total_offset_9[6:0] ? field_byte_9 : _GEN_1765; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1862 = 7'h25 == total_offset_9[6:0] ? field_byte_9 : _GEN_1766; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1863 = 7'h26 == total_offset_9[6:0] ? field_byte_9 : _GEN_1767; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1864 = 7'h27 == total_offset_9[6:0] ? field_byte_9 : _GEN_1768; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1865 = 7'h28 == total_offset_9[6:0] ? field_byte_9 : _GEN_1769; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1866 = 7'h29 == total_offset_9[6:0] ? field_byte_9 : _GEN_1770; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1867 = 7'h2a == total_offset_9[6:0] ? field_byte_9 : _GEN_1771; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1868 = 7'h2b == total_offset_9[6:0] ? field_byte_9 : _GEN_1772; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1869 = 7'h2c == total_offset_9[6:0] ? field_byte_9 : _GEN_1773; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1870 = 7'h2d == total_offset_9[6:0] ? field_byte_9 : _GEN_1774; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1871 = 7'h2e == total_offset_9[6:0] ? field_byte_9 : _GEN_1775; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1872 = 7'h2f == total_offset_9[6:0] ? field_byte_9 : _GEN_1776; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1873 = 7'h30 == total_offset_9[6:0] ? field_byte_9 : _GEN_1777; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1874 = 7'h31 == total_offset_9[6:0] ? field_byte_9 : _GEN_1778; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1875 = 7'h32 == total_offset_9[6:0] ? field_byte_9 : _GEN_1779; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1876 = 7'h33 == total_offset_9[6:0] ? field_byte_9 : _GEN_1780; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1877 = 7'h34 == total_offset_9[6:0] ? field_byte_9 : _GEN_1781; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1878 = 7'h35 == total_offset_9[6:0] ? field_byte_9 : _GEN_1782; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1879 = 7'h36 == total_offset_9[6:0] ? field_byte_9 : _GEN_1783; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1880 = 7'h37 == total_offset_9[6:0] ? field_byte_9 : _GEN_1784; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1881 = 7'h38 == total_offset_9[6:0] ? field_byte_9 : _GEN_1785; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1882 = 7'h39 == total_offset_9[6:0] ? field_byte_9 : _GEN_1786; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1883 = 7'h3a == total_offset_9[6:0] ? field_byte_9 : _GEN_1787; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1884 = 7'h3b == total_offset_9[6:0] ? field_byte_9 : _GEN_1788; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1885 = 7'h3c == total_offset_9[6:0] ? field_byte_9 : _GEN_1789; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1886 = 7'h3d == total_offset_9[6:0] ? field_byte_9 : _GEN_1790; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1887 = 7'h3e == total_offset_9[6:0] ? field_byte_9 : _GEN_1791; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1888 = 7'h3f == total_offset_9[6:0] ? field_byte_9 : _GEN_1792; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1889 = 7'h40 == total_offset_9[6:0] ? field_byte_9 : _GEN_1793; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1890 = 7'h41 == total_offset_9[6:0] ? field_byte_9 : _GEN_1794; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1891 = 7'h42 == total_offset_9[6:0] ? field_byte_9 : _GEN_1795; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1892 = 7'h43 == total_offset_9[6:0] ? field_byte_9 : _GEN_1796; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1893 = 7'h44 == total_offset_9[6:0] ? field_byte_9 : _GEN_1797; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1894 = 7'h45 == total_offset_9[6:0] ? field_byte_9 : _GEN_1798; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1895 = 7'h46 == total_offset_9[6:0] ? field_byte_9 : _GEN_1799; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1896 = 7'h47 == total_offset_9[6:0] ? field_byte_9 : _GEN_1800; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1897 = 7'h48 == total_offset_9[6:0] ? field_byte_9 : _GEN_1801; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1898 = 7'h49 == total_offset_9[6:0] ? field_byte_9 : _GEN_1802; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1899 = 7'h4a == total_offset_9[6:0] ? field_byte_9 : _GEN_1803; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1900 = 7'h4b == total_offset_9[6:0] ? field_byte_9 : _GEN_1804; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1901 = 7'h4c == total_offset_9[6:0] ? field_byte_9 : _GEN_1805; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1902 = 7'h4d == total_offset_9[6:0] ? field_byte_9 : _GEN_1806; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1903 = 7'h4e == total_offset_9[6:0] ? field_byte_9 : _GEN_1807; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1904 = 7'h4f == total_offset_9[6:0] ? field_byte_9 : _GEN_1808; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1905 = 7'h50 == total_offset_9[6:0] ? field_byte_9 : _GEN_1809; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1906 = 7'h51 == total_offset_9[6:0] ? field_byte_9 : _GEN_1810; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1907 = 7'h52 == total_offset_9[6:0] ? field_byte_9 : _GEN_1811; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1908 = 7'h53 == total_offset_9[6:0] ? field_byte_9 : _GEN_1812; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1909 = 7'h54 == total_offset_9[6:0] ? field_byte_9 : _GEN_1813; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1910 = 7'h55 == total_offset_9[6:0] ? field_byte_9 : _GEN_1814; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1911 = 7'h56 == total_offset_9[6:0] ? field_byte_9 : _GEN_1815; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1912 = 7'h57 == total_offset_9[6:0] ? field_byte_9 : _GEN_1816; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1913 = 7'h58 == total_offset_9[6:0] ? field_byte_9 : _GEN_1817; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1914 = 7'h59 == total_offset_9[6:0] ? field_byte_9 : _GEN_1818; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1915 = 7'h5a == total_offset_9[6:0] ? field_byte_9 : _GEN_1819; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1916 = 7'h5b == total_offset_9[6:0] ? field_byte_9 : _GEN_1820; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1917 = 7'h5c == total_offset_9[6:0] ? field_byte_9 : _GEN_1821; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1918 = 7'h5d == total_offset_9[6:0] ? field_byte_9 : _GEN_1822; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1919 = 7'h5e == total_offset_9[6:0] ? field_byte_9 : _GEN_1823; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1920 = 7'h5f == total_offset_9[6:0] ? field_byte_9 : _GEN_1824; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_1921 = 8'h1 < length_1 ? _GEN_1825 : _GEN_1729; // @[executor.scala 290:56]
  wire [7:0] _GEN_1922 = 8'h1 < length_1 ? _GEN_1826 : _GEN_1730; // @[executor.scala 290:56]
  wire [7:0] _GEN_1923 = 8'h1 < length_1 ? _GEN_1827 : _GEN_1731; // @[executor.scala 290:56]
  wire [7:0] _GEN_1924 = 8'h1 < length_1 ? _GEN_1828 : _GEN_1732; // @[executor.scala 290:56]
  wire [7:0] _GEN_1925 = 8'h1 < length_1 ? _GEN_1829 : _GEN_1733; // @[executor.scala 290:56]
  wire [7:0] _GEN_1926 = 8'h1 < length_1 ? _GEN_1830 : _GEN_1734; // @[executor.scala 290:56]
  wire [7:0] _GEN_1927 = 8'h1 < length_1 ? _GEN_1831 : _GEN_1735; // @[executor.scala 290:56]
  wire [7:0] _GEN_1928 = 8'h1 < length_1 ? _GEN_1832 : _GEN_1736; // @[executor.scala 290:56]
  wire [7:0] _GEN_1929 = 8'h1 < length_1 ? _GEN_1833 : _GEN_1737; // @[executor.scala 290:56]
  wire [7:0] _GEN_1930 = 8'h1 < length_1 ? _GEN_1834 : _GEN_1738; // @[executor.scala 290:56]
  wire [7:0] _GEN_1931 = 8'h1 < length_1 ? _GEN_1835 : _GEN_1739; // @[executor.scala 290:56]
  wire [7:0] _GEN_1932 = 8'h1 < length_1 ? _GEN_1836 : _GEN_1740; // @[executor.scala 290:56]
  wire [7:0] _GEN_1933 = 8'h1 < length_1 ? _GEN_1837 : _GEN_1741; // @[executor.scala 290:56]
  wire [7:0] _GEN_1934 = 8'h1 < length_1 ? _GEN_1838 : _GEN_1742; // @[executor.scala 290:56]
  wire [7:0] _GEN_1935 = 8'h1 < length_1 ? _GEN_1839 : _GEN_1743; // @[executor.scala 290:56]
  wire [7:0] _GEN_1936 = 8'h1 < length_1 ? _GEN_1840 : _GEN_1744; // @[executor.scala 290:56]
  wire [7:0] _GEN_1937 = 8'h1 < length_1 ? _GEN_1841 : _GEN_1745; // @[executor.scala 290:56]
  wire [7:0] _GEN_1938 = 8'h1 < length_1 ? _GEN_1842 : _GEN_1746; // @[executor.scala 290:56]
  wire [7:0] _GEN_1939 = 8'h1 < length_1 ? _GEN_1843 : _GEN_1747; // @[executor.scala 290:56]
  wire [7:0] _GEN_1940 = 8'h1 < length_1 ? _GEN_1844 : _GEN_1748; // @[executor.scala 290:56]
  wire [7:0] _GEN_1941 = 8'h1 < length_1 ? _GEN_1845 : _GEN_1749; // @[executor.scala 290:56]
  wire [7:0] _GEN_1942 = 8'h1 < length_1 ? _GEN_1846 : _GEN_1750; // @[executor.scala 290:56]
  wire [7:0] _GEN_1943 = 8'h1 < length_1 ? _GEN_1847 : _GEN_1751; // @[executor.scala 290:56]
  wire [7:0] _GEN_1944 = 8'h1 < length_1 ? _GEN_1848 : _GEN_1752; // @[executor.scala 290:56]
  wire [7:0] _GEN_1945 = 8'h1 < length_1 ? _GEN_1849 : _GEN_1753; // @[executor.scala 290:56]
  wire [7:0] _GEN_1946 = 8'h1 < length_1 ? _GEN_1850 : _GEN_1754; // @[executor.scala 290:56]
  wire [7:0] _GEN_1947 = 8'h1 < length_1 ? _GEN_1851 : _GEN_1755; // @[executor.scala 290:56]
  wire [7:0] _GEN_1948 = 8'h1 < length_1 ? _GEN_1852 : _GEN_1756; // @[executor.scala 290:56]
  wire [7:0] _GEN_1949 = 8'h1 < length_1 ? _GEN_1853 : _GEN_1757; // @[executor.scala 290:56]
  wire [7:0] _GEN_1950 = 8'h1 < length_1 ? _GEN_1854 : _GEN_1758; // @[executor.scala 290:56]
  wire [7:0] _GEN_1951 = 8'h1 < length_1 ? _GEN_1855 : _GEN_1759; // @[executor.scala 290:56]
  wire [7:0] _GEN_1952 = 8'h1 < length_1 ? _GEN_1856 : _GEN_1760; // @[executor.scala 290:56]
  wire [7:0] _GEN_1953 = 8'h1 < length_1 ? _GEN_1857 : _GEN_1761; // @[executor.scala 290:56]
  wire [7:0] _GEN_1954 = 8'h1 < length_1 ? _GEN_1858 : _GEN_1762; // @[executor.scala 290:56]
  wire [7:0] _GEN_1955 = 8'h1 < length_1 ? _GEN_1859 : _GEN_1763; // @[executor.scala 290:56]
  wire [7:0] _GEN_1956 = 8'h1 < length_1 ? _GEN_1860 : _GEN_1764; // @[executor.scala 290:56]
  wire [7:0] _GEN_1957 = 8'h1 < length_1 ? _GEN_1861 : _GEN_1765; // @[executor.scala 290:56]
  wire [7:0] _GEN_1958 = 8'h1 < length_1 ? _GEN_1862 : _GEN_1766; // @[executor.scala 290:56]
  wire [7:0] _GEN_1959 = 8'h1 < length_1 ? _GEN_1863 : _GEN_1767; // @[executor.scala 290:56]
  wire [7:0] _GEN_1960 = 8'h1 < length_1 ? _GEN_1864 : _GEN_1768; // @[executor.scala 290:56]
  wire [7:0] _GEN_1961 = 8'h1 < length_1 ? _GEN_1865 : _GEN_1769; // @[executor.scala 290:56]
  wire [7:0] _GEN_1962 = 8'h1 < length_1 ? _GEN_1866 : _GEN_1770; // @[executor.scala 290:56]
  wire [7:0] _GEN_1963 = 8'h1 < length_1 ? _GEN_1867 : _GEN_1771; // @[executor.scala 290:56]
  wire [7:0] _GEN_1964 = 8'h1 < length_1 ? _GEN_1868 : _GEN_1772; // @[executor.scala 290:56]
  wire [7:0] _GEN_1965 = 8'h1 < length_1 ? _GEN_1869 : _GEN_1773; // @[executor.scala 290:56]
  wire [7:0] _GEN_1966 = 8'h1 < length_1 ? _GEN_1870 : _GEN_1774; // @[executor.scala 290:56]
  wire [7:0] _GEN_1967 = 8'h1 < length_1 ? _GEN_1871 : _GEN_1775; // @[executor.scala 290:56]
  wire [7:0] _GEN_1968 = 8'h1 < length_1 ? _GEN_1872 : _GEN_1776; // @[executor.scala 290:56]
  wire [7:0] _GEN_1969 = 8'h1 < length_1 ? _GEN_1873 : _GEN_1777; // @[executor.scala 290:56]
  wire [7:0] _GEN_1970 = 8'h1 < length_1 ? _GEN_1874 : _GEN_1778; // @[executor.scala 290:56]
  wire [7:0] _GEN_1971 = 8'h1 < length_1 ? _GEN_1875 : _GEN_1779; // @[executor.scala 290:56]
  wire [7:0] _GEN_1972 = 8'h1 < length_1 ? _GEN_1876 : _GEN_1780; // @[executor.scala 290:56]
  wire [7:0] _GEN_1973 = 8'h1 < length_1 ? _GEN_1877 : _GEN_1781; // @[executor.scala 290:56]
  wire [7:0] _GEN_1974 = 8'h1 < length_1 ? _GEN_1878 : _GEN_1782; // @[executor.scala 290:56]
  wire [7:0] _GEN_1975 = 8'h1 < length_1 ? _GEN_1879 : _GEN_1783; // @[executor.scala 290:56]
  wire [7:0] _GEN_1976 = 8'h1 < length_1 ? _GEN_1880 : _GEN_1784; // @[executor.scala 290:56]
  wire [7:0] _GEN_1977 = 8'h1 < length_1 ? _GEN_1881 : _GEN_1785; // @[executor.scala 290:56]
  wire [7:0] _GEN_1978 = 8'h1 < length_1 ? _GEN_1882 : _GEN_1786; // @[executor.scala 290:56]
  wire [7:0] _GEN_1979 = 8'h1 < length_1 ? _GEN_1883 : _GEN_1787; // @[executor.scala 290:56]
  wire [7:0] _GEN_1980 = 8'h1 < length_1 ? _GEN_1884 : _GEN_1788; // @[executor.scala 290:56]
  wire [7:0] _GEN_1981 = 8'h1 < length_1 ? _GEN_1885 : _GEN_1789; // @[executor.scala 290:56]
  wire [7:0] _GEN_1982 = 8'h1 < length_1 ? _GEN_1886 : _GEN_1790; // @[executor.scala 290:56]
  wire [7:0] _GEN_1983 = 8'h1 < length_1 ? _GEN_1887 : _GEN_1791; // @[executor.scala 290:56]
  wire [7:0] _GEN_1984 = 8'h1 < length_1 ? _GEN_1888 : _GEN_1792; // @[executor.scala 290:56]
  wire [7:0] _GEN_1985 = 8'h1 < length_1 ? _GEN_1889 : _GEN_1793; // @[executor.scala 290:56]
  wire [7:0] _GEN_1986 = 8'h1 < length_1 ? _GEN_1890 : _GEN_1794; // @[executor.scala 290:56]
  wire [7:0] _GEN_1987 = 8'h1 < length_1 ? _GEN_1891 : _GEN_1795; // @[executor.scala 290:56]
  wire [7:0] _GEN_1988 = 8'h1 < length_1 ? _GEN_1892 : _GEN_1796; // @[executor.scala 290:56]
  wire [7:0] _GEN_1989 = 8'h1 < length_1 ? _GEN_1893 : _GEN_1797; // @[executor.scala 290:56]
  wire [7:0] _GEN_1990 = 8'h1 < length_1 ? _GEN_1894 : _GEN_1798; // @[executor.scala 290:56]
  wire [7:0] _GEN_1991 = 8'h1 < length_1 ? _GEN_1895 : _GEN_1799; // @[executor.scala 290:56]
  wire [7:0] _GEN_1992 = 8'h1 < length_1 ? _GEN_1896 : _GEN_1800; // @[executor.scala 290:56]
  wire [7:0] _GEN_1993 = 8'h1 < length_1 ? _GEN_1897 : _GEN_1801; // @[executor.scala 290:56]
  wire [7:0] _GEN_1994 = 8'h1 < length_1 ? _GEN_1898 : _GEN_1802; // @[executor.scala 290:56]
  wire [7:0] _GEN_1995 = 8'h1 < length_1 ? _GEN_1899 : _GEN_1803; // @[executor.scala 290:56]
  wire [7:0] _GEN_1996 = 8'h1 < length_1 ? _GEN_1900 : _GEN_1804; // @[executor.scala 290:56]
  wire [7:0] _GEN_1997 = 8'h1 < length_1 ? _GEN_1901 : _GEN_1805; // @[executor.scala 290:56]
  wire [7:0] _GEN_1998 = 8'h1 < length_1 ? _GEN_1902 : _GEN_1806; // @[executor.scala 290:56]
  wire [7:0] _GEN_1999 = 8'h1 < length_1 ? _GEN_1903 : _GEN_1807; // @[executor.scala 290:56]
  wire [7:0] _GEN_2000 = 8'h1 < length_1 ? _GEN_1904 : _GEN_1808; // @[executor.scala 290:56]
  wire [7:0] _GEN_2001 = 8'h1 < length_1 ? _GEN_1905 : _GEN_1809; // @[executor.scala 290:56]
  wire [7:0] _GEN_2002 = 8'h1 < length_1 ? _GEN_1906 : _GEN_1810; // @[executor.scala 290:56]
  wire [7:0] _GEN_2003 = 8'h1 < length_1 ? _GEN_1907 : _GEN_1811; // @[executor.scala 290:56]
  wire [7:0] _GEN_2004 = 8'h1 < length_1 ? _GEN_1908 : _GEN_1812; // @[executor.scala 290:56]
  wire [7:0] _GEN_2005 = 8'h1 < length_1 ? _GEN_1909 : _GEN_1813; // @[executor.scala 290:56]
  wire [7:0] _GEN_2006 = 8'h1 < length_1 ? _GEN_1910 : _GEN_1814; // @[executor.scala 290:56]
  wire [7:0] _GEN_2007 = 8'h1 < length_1 ? _GEN_1911 : _GEN_1815; // @[executor.scala 290:56]
  wire [7:0] _GEN_2008 = 8'h1 < length_1 ? _GEN_1912 : _GEN_1816; // @[executor.scala 290:56]
  wire [7:0] _GEN_2009 = 8'h1 < length_1 ? _GEN_1913 : _GEN_1817; // @[executor.scala 290:56]
  wire [7:0] _GEN_2010 = 8'h1 < length_1 ? _GEN_1914 : _GEN_1818; // @[executor.scala 290:56]
  wire [7:0] _GEN_2011 = 8'h1 < length_1 ? _GEN_1915 : _GEN_1819; // @[executor.scala 290:56]
  wire [7:0] _GEN_2012 = 8'h1 < length_1 ? _GEN_1916 : _GEN_1820; // @[executor.scala 290:56]
  wire [7:0] _GEN_2013 = 8'h1 < length_1 ? _GEN_1917 : _GEN_1821; // @[executor.scala 290:56]
  wire [7:0] _GEN_2014 = 8'h1 < length_1 ? _GEN_1918 : _GEN_1822; // @[executor.scala 290:56]
  wire [7:0] _GEN_2015 = 8'h1 < length_1 ? _GEN_1919 : _GEN_1823; // @[executor.scala 290:56]
  wire [7:0] _GEN_2016 = 8'h1 < length_1 ? _GEN_1920 : _GEN_1824; // @[executor.scala 290:56]
  wire [7:0] field_byte_10 = field_1[47:40]; // @[executor.scala 287:53]
  wire [7:0] total_offset_10 = offset_1 + 8'h2; // @[executor.scala 289:53]
  wire [7:0] _GEN_2017 = 7'h0 == total_offset_10[6:0] ? field_byte_10 : _GEN_1921; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2018 = 7'h1 == total_offset_10[6:0] ? field_byte_10 : _GEN_1922; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2019 = 7'h2 == total_offset_10[6:0] ? field_byte_10 : _GEN_1923; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2020 = 7'h3 == total_offset_10[6:0] ? field_byte_10 : _GEN_1924; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2021 = 7'h4 == total_offset_10[6:0] ? field_byte_10 : _GEN_1925; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2022 = 7'h5 == total_offset_10[6:0] ? field_byte_10 : _GEN_1926; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2023 = 7'h6 == total_offset_10[6:0] ? field_byte_10 : _GEN_1927; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2024 = 7'h7 == total_offset_10[6:0] ? field_byte_10 : _GEN_1928; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2025 = 7'h8 == total_offset_10[6:0] ? field_byte_10 : _GEN_1929; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2026 = 7'h9 == total_offset_10[6:0] ? field_byte_10 : _GEN_1930; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2027 = 7'ha == total_offset_10[6:0] ? field_byte_10 : _GEN_1931; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2028 = 7'hb == total_offset_10[6:0] ? field_byte_10 : _GEN_1932; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2029 = 7'hc == total_offset_10[6:0] ? field_byte_10 : _GEN_1933; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2030 = 7'hd == total_offset_10[6:0] ? field_byte_10 : _GEN_1934; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2031 = 7'he == total_offset_10[6:0] ? field_byte_10 : _GEN_1935; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2032 = 7'hf == total_offset_10[6:0] ? field_byte_10 : _GEN_1936; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2033 = 7'h10 == total_offset_10[6:0] ? field_byte_10 : _GEN_1937; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2034 = 7'h11 == total_offset_10[6:0] ? field_byte_10 : _GEN_1938; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2035 = 7'h12 == total_offset_10[6:0] ? field_byte_10 : _GEN_1939; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2036 = 7'h13 == total_offset_10[6:0] ? field_byte_10 : _GEN_1940; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2037 = 7'h14 == total_offset_10[6:0] ? field_byte_10 : _GEN_1941; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2038 = 7'h15 == total_offset_10[6:0] ? field_byte_10 : _GEN_1942; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2039 = 7'h16 == total_offset_10[6:0] ? field_byte_10 : _GEN_1943; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2040 = 7'h17 == total_offset_10[6:0] ? field_byte_10 : _GEN_1944; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2041 = 7'h18 == total_offset_10[6:0] ? field_byte_10 : _GEN_1945; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2042 = 7'h19 == total_offset_10[6:0] ? field_byte_10 : _GEN_1946; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2043 = 7'h1a == total_offset_10[6:0] ? field_byte_10 : _GEN_1947; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2044 = 7'h1b == total_offset_10[6:0] ? field_byte_10 : _GEN_1948; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2045 = 7'h1c == total_offset_10[6:0] ? field_byte_10 : _GEN_1949; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2046 = 7'h1d == total_offset_10[6:0] ? field_byte_10 : _GEN_1950; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2047 = 7'h1e == total_offset_10[6:0] ? field_byte_10 : _GEN_1951; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2048 = 7'h1f == total_offset_10[6:0] ? field_byte_10 : _GEN_1952; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2049 = 7'h20 == total_offset_10[6:0] ? field_byte_10 : _GEN_1953; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2050 = 7'h21 == total_offset_10[6:0] ? field_byte_10 : _GEN_1954; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2051 = 7'h22 == total_offset_10[6:0] ? field_byte_10 : _GEN_1955; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2052 = 7'h23 == total_offset_10[6:0] ? field_byte_10 : _GEN_1956; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2053 = 7'h24 == total_offset_10[6:0] ? field_byte_10 : _GEN_1957; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2054 = 7'h25 == total_offset_10[6:0] ? field_byte_10 : _GEN_1958; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2055 = 7'h26 == total_offset_10[6:0] ? field_byte_10 : _GEN_1959; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2056 = 7'h27 == total_offset_10[6:0] ? field_byte_10 : _GEN_1960; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2057 = 7'h28 == total_offset_10[6:0] ? field_byte_10 : _GEN_1961; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2058 = 7'h29 == total_offset_10[6:0] ? field_byte_10 : _GEN_1962; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2059 = 7'h2a == total_offset_10[6:0] ? field_byte_10 : _GEN_1963; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2060 = 7'h2b == total_offset_10[6:0] ? field_byte_10 : _GEN_1964; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2061 = 7'h2c == total_offset_10[6:0] ? field_byte_10 : _GEN_1965; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2062 = 7'h2d == total_offset_10[6:0] ? field_byte_10 : _GEN_1966; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2063 = 7'h2e == total_offset_10[6:0] ? field_byte_10 : _GEN_1967; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2064 = 7'h2f == total_offset_10[6:0] ? field_byte_10 : _GEN_1968; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2065 = 7'h30 == total_offset_10[6:0] ? field_byte_10 : _GEN_1969; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2066 = 7'h31 == total_offset_10[6:0] ? field_byte_10 : _GEN_1970; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2067 = 7'h32 == total_offset_10[6:0] ? field_byte_10 : _GEN_1971; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2068 = 7'h33 == total_offset_10[6:0] ? field_byte_10 : _GEN_1972; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2069 = 7'h34 == total_offset_10[6:0] ? field_byte_10 : _GEN_1973; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2070 = 7'h35 == total_offset_10[6:0] ? field_byte_10 : _GEN_1974; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2071 = 7'h36 == total_offset_10[6:0] ? field_byte_10 : _GEN_1975; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2072 = 7'h37 == total_offset_10[6:0] ? field_byte_10 : _GEN_1976; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2073 = 7'h38 == total_offset_10[6:0] ? field_byte_10 : _GEN_1977; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2074 = 7'h39 == total_offset_10[6:0] ? field_byte_10 : _GEN_1978; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2075 = 7'h3a == total_offset_10[6:0] ? field_byte_10 : _GEN_1979; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2076 = 7'h3b == total_offset_10[6:0] ? field_byte_10 : _GEN_1980; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2077 = 7'h3c == total_offset_10[6:0] ? field_byte_10 : _GEN_1981; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2078 = 7'h3d == total_offset_10[6:0] ? field_byte_10 : _GEN_1982; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2079 = 7'h3e == total_offset_10[6:0] ? field_byte_10 : _GEN_1983; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2080 = 7'h3f == total_offset_10[6:0] ? field_byte_10 : _GEN_1984; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2081 = 7'h40 == total_offset_10[6:0] ? field_byte_10 : _GEN_1985; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2082 = 7'h41 == total_offset_10[6:0] ? field_byte_10 : _GEN_1986; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2083 = 7'h42 == total_offset_10[6:0] ? field_byte_10 : _GEN_1987; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2084 = 7'h43 == total_offset_10[6:0] ? field_byte_10 : _GEN_1988; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2085 = 7'h44 == total_offset_10[6:0] ? field_byte_10 : _GEN_1989; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2086 = 7'h45 == total_offset_10[6:0] ? field_byte_10 : _GEN_1990; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2087 = 7'h46 == total_offset_10[6:0] ? field_byte_10 : _GEN_1991; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2088 = 7'h47 == total_offset_10[6:0] ? field_byte_10 : _GEN_1992; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2089 = 7'h48 == total_offset_10[6:0] ? field_byte_10 : _GEN_1993; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2090 = 7'h49 == total_offset_10[6:0] ? field_byte_10 : _GEN_1994; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2091 = 7'h4a == total_offset_10[6:0] ? field_byte_10 : _GEN_1995; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2092 = 7'h4b == total_offset_10[6:0] ? field_byte_10 : _GEN_1996; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2093 = 7'h4c == total_offset_10[6:0] ? field_byte_10 : _GEN_1997; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2094 = 7'h4d == total_offset_10[6:0] ? field_byte_10 : _GEN_1998; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2095 = 7'h4e == total_offset_10[6:0] ? field_byte_10 : _GEN_1999; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2096 = 7'h4f == total_offset_10[6:0] ? field_byte_10 : _GEN_2000; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2097 = 7'h50 == total_offset_10[6:0] ? field_byte_10 : _GEN_2001; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2098 = 7'h51 == total_offset_10[6:0] ? field_byte_10 : _GEN_2002; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2099 = 7'h52 == total_offset_10[6:0] ? field_byte_10 : _GEN_2003; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2100 = 7'h53 == total_offset_10[6:0] ? field_byte_10 : _GEN_2004; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2101 = 7'h54 == total_offset_10[6:0] ? field_byte_10 : _GEN_2005; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2102 = 7'h55 == total_offset_10[6:0] ? field_byte_10 : _GEN_2006; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2103 = 7'h56 == total_offset_10[6:0] ? field_byte_10 : _GEN_2007; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2104 = 7'h57 == total_offset_10[6:0] ? field_byte_10 : _GEN_2008; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2105 = 7'h58 == total_offset_10[6:0] ? field_byte_10 : _GEN_2009; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2106 = 7'h59 == total_offset_10[6:0] ? field_byte_10 : _GEN_2010; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2107 = 7'h5a == total_offset_10[6:0] ? field_byte_10 : _GEN_2011; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2108 = 7'h5b == total_offset_10[6:0] ? field_byte_10 : _GEN_2012; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2109 = 7'h5c == total_offset_10[6:0] ? field_byte_10 : _GEN_2013; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2110 = 7'h5d == total_offset_10[6:0] ? field_byte_10 : _GEN_2014; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2111 = 7'h5e == total_offset_10[6:0] ? field_byte_10 : _GEN_2015; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2112 = 7'h5f == total_offset_10[6:0] ? field_byte_10 : _GEN_2016; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2113 = 8'h2 < length_1 ? _GEN_2017 : _GEN_1921; // @[executor.scala 290:56]
  wire [7:0] _GEN_2114 = 8'h2 < length_1 ? _GEN_2018 : _GEN_1922; // @[executor.scala 290:56]
  wire [7:0] _GEN_2115 = 8'h2 < length_1 ? _GEN_2019 : _GEN_1923; // @[executor.scala 290:56]
  wire [7:0] _GEN_2116 = 8'h2 < length_1 ? _GEN_2020 : _GEN_1924; // @[executor.scala 290:56]
  wire [7:0] _GEN_2117 = 8'h2 < length_1 ? _GEN_2021 : _GEN_1925; // @[executor.scala 290:56]
  wire [7:0] _GEN_2118 = 8'h2 < length_1 ? _GEN_2022 : _GEN_1926; // @[executor.scala 290:56]
  wire [7:0] _GEN_2119 = 8'h2 < length_1 ? _GEN_2023 : _GEN_1927; // @[executor.scala 290:56]
  wire [7:0] _GEN_2120 = 8'h2 < length_1 ? _GEN_2024 : _GEN_1928; // @[executor.scala 290:56]
  wire [7:0] _GEN_2121 = 8'h2 < length_1 ? _GEN_2025 : _GEN_1929; // @[executor.scala 290:56]
  wire [7:0] _GEN_2122 = 8'h2 < length_1 ? _GEN_2026 : _GEN_1930; // @[executor.scala 290:56]
  wire [7:0] _GEN_2123 = 8'h2 < length_1 ? _GEN_2027 : _GEN_1931; // @[executor.scala 290:56]
  wire [7:0] _GEN_2124 = 8'h2 < length_1 ? _GEN_2028 : _GEN_1932; // @[executor.scala 290:56]
  wire [7:0] _GEN_2125 = 8'h2 < length_1 ? _GEN_2029 : _GEN_1933; // @[executor.scala 290:56]
  wire [7:0] _GEN_2126 = 8'h2 < length_1 ? _GEN_2030 : _GEN_1934; // @[executor.scala 290:56]
  wire [7:0] _GEN_2127 = 8'h2 < length_1 ? _GEN_2031 : _GEN_1935; // @[executor.scala 290:56]
  wire [7:0] _GEN_2128 = 8'h2 < length_1 ? _GEN_2032 : _GEN_1936; // @[executor.scala 290:56]
  wire [7:0] _GEN_2129 = 8'h2 < length_1 ? _GEN_2033 : _GEN_1937; // @[executor.scala 290:56]
  wire [7:0] _GEN_2130 = 8'h2 < length_1 ? _GEN_2034 : _GEN_1938; // @[executor.scala 290:56]
  wire [7:0] _GEN_2131 = 8'h2 < length_1 ? _GEN_2035 : _GEN_1939; // @[executor.scala 290:56]
  wire [7:0] _GEN_2132 = 8'h2 < length_1 ? _GEN_2036 : _GEN_1940; // @[executor.scala 290:56]
  wire [7:0] _GEN_2133 = 8'h2 < length_1 ? _GEN_2037 : _GEN_1941; // @[executor.scala 290:56]
  wire [7:0] _GEN_2134 = 8'h2 < length_1 ? _GEN_2038 : _GEN_1942; // @[executor.scala 290:56]
  wire [7:0] _GEN_2135 = 8'h2 < length_1 ? _GEN_2039 : _GEN_1943; // @[executor.scala 290:56]
  wire [7:0] _GEN_2136 = 8'h2 < length_1 ? _GEN_2040 : _GEN_1944; // @[executor.scala 290:56]
  wire [7:0] _GEN_2137 = 8'h2 < length_1 ? _GEN_2041 : _GEN_1945; // @[executor.scala 290:56]
  wire [7:0] _GEN_2138 = 8'h2 < length_1 ? _GEN_2042 : _GEN_1946; // @[executor.scala 290:56]
  wire [7:0] _GEN_2139 = 8'h2 < length_1 ? _GEN_2043 : _GEN_1947; // @[executor.scala 290:56]
  wire [7:0] _GEN_2140 = 8'h2 < length_1 ? _GEN_2044 : _GEN_1948; // @[executor.scala 290:56]
  wire [7:0] _GEN_2141 = 8'h2 < length_1 ? _GEN_2045 : _GEN_1949; // @[executor.scala 290:56]
  wire [7:0] _GEN_2142 = 8'h2 < length_1 ? _GEN_2046 : _GEN_1950; // @[executor.scala 290:56]
  wire [7:0] _GEN_2143 = 8'h2 < length_1 ? _GEN_2047 : _GEN_1951; // @[executor.scala 290:56]
  wire [7:0] _GEN_2144 = 8'h2 < length_1 ? _GEN_2048 : _GEN_1952; // @[executor.scala 290:56]
  wire [7:0] _GEN_2145 = 8'h2 < length_1 ? _GEN_2049 : _GEN_1953; // @[executor.scala 290:56]
  wire [7:0] _GEN_2146 = 8'h2 < length_1 ? _GEN_2050 : _GEN_1954; // @[executor.scala 290:56]
  wire [7:0] _GEN_2147 = 8'h2 < length_1 ? _GEN_2051 : _GEN_1955; // @[executor.scala 290:56]
  wire [7:0] _GEN_2148 = 8'h2 < length_1 ? _GEN_2052 : _GEN_1956; // @[executor.scala 290:56]
  wire [7:0] _GEN_2149 = 8'h2 < length_1 ? _GEN_2053 : _GEN_1957; // @[executor.scala 290:56]
  wire [7:0] _GEN_2150 = 8'h2 < length_1 ? _GEN_2054 : _GEN_1958; // @[executor.scala 290:56]
  wire [7:0] _GEN_2151 = 8'h2 < length_1 ? _GEN_2055 : _GEN_1959; // @[executor.scala 290:56]
  wire [7:0] _GEN_2152 = 8'h2 < length_1 ? _GEN_2056 : _GEN_1960; // @[executor.scala 290:56]
  wire [7:0] _GEN_2153 = 8'h2 < length_1 ? _GEN_2057 : _GEN_1961; // @[executor.scala 290:56]
  wire [7:0] _GEN_2154 = 8'h2 < length_1 ? _GEN_2058 : _GEN_1962; // @[executor.scala 290:56]
  wire [7:0] _GEN_2155 = 8'h2 < length_1 ? _GEN_2059 : _GEN_1963; // @[executor.scala 290:56]
  wire [7:0] _GEN_2156 = 8'h2 < length_1 ? _GEN_2060 : _GEN_1964; // @[executor.scala 290:56]
  wire [7:0] _GEN_2157 = 8'h2 < length_1 ? _GEN_2061 : _GEN_1965; // @[executor.scala 290:56]
  wire [7:0] _GEN_2158 = 8'h2 < length_1 ? _GEN_2062 : _GEN_1966; // @[executor.scala 290:56]
  wire [7:0] _GEN_2159 = 8'h2 < length_1 ? _GEN_2063 : _GEN_1967; // @[executor.scala 290:56]
  wire [7:0] _GEN_2160 = 8'h2 < length_1 ? _GEN_2064 : _GEN_1968; // @[executor.scala 290:56]
  wire [7:0] _GEN_2161 = 8'h2 < length_1 ? _GEN_2065 : _GEN_1969; // @[executor.scala 290:56]
  wire [7:0] _GEN_2162 = 8'h2 < length_1 ? _GEN_2066 : _GEN_1970; // @[executor.scala 290:56]
  wire [7:0] _GEN_2163 = 8'h2 < length_1 ? _GEN_2067 : _GEN_1971; // @[executor.scala 290:56]
  wire [7:0] _GEN_2164 = 8'h2 < length_1 ? _GEN_2068 : _GEN_1972; // @[executor.scala 290:56]
  wire [7:0] _GEN_2165 = 8'h2 < length_1 ? _GEN_2069 : _GEN_1973; // @[executor.scala 290:56]
  wire [7:0] _GEN_2166 = 8'h2 < length_1 ? _GEN_2070 : _GEN_1974; // @[executor.scala 290:56]
  wire [7:0] _GEN_2167 = 8'h2 < length_1 ? _GEN_2071 : _GEN_1975; // @[executor.scala 290:56]
  wire [7:0] _GEN_2168 = 8'h2 < length_1 ? _GEN_2072 : _GEN_1976; // @[executor.scala 290:56]
  wire [7:0] _GEN_2169 = 8'h2 < length_1 ? _GEN_2073 : _GEN_1977; // @[executor.scala 290:56]
  wire [7:0] _GEN_2170 = 8'h2 < length_1 ? _GEN_2074 : _GEN_1978; // @[executor.scala 290:56]
  wire [7:0] _GEN_2171 = 8'h2 < length_1 ? _GEN_2075 : _GEN_1979; // @[executor.scala 290:56]
  wire [7:0] _GEN_2172 = 8'h2 < length_1 ? _GEN_2076 : _GEN_1980; // @[executor.scala 290:56]
  wire [7:0] _GEN_2173 = 8'h2 < length_1 ? _GEN_2077 : _GEN_1981; // @[executor.scala 290:56]
  wire [7:0] _GEN_2174 = 8'h2 < length_1 ? _GEN_2078 : _GEN_1982; // @[executor.scala 290:56]
  wire [7:0] _GEN_2175 = 8'h2 < length_1 ? _GEN_2079 : _GEN_1983; // @[executor.scala 290:56]
  wire [7:0] _GEN_2176 = 8'h2 < length_1 ? _GEN_2080 : _GEN_1984; // @[executor.scala 290:56]
  wire [7:0] _GEN_2177 = 8'h2 < length_1 ? _GEN_2081 : _GEN_1985; // @[executor.scala 290:56]
  wire [7:0] _GEN_2178 = 8'h2 < length_1 ? _GEN_2082 : _GEN_1986; // @[executor.scala 290:56]
  wire [7:0] _GEN_2179 = 8'h2 < length_1 ? _GEN_2083 : _GEN_1987; // @[executor.scala 290:56]
  wire [7:0] _GEN_2180 = 8'h2 < length_1 ? _GEN_2084 : _GEN_1988; // @[executor.scala 290:56]
  wire [7:0] _GEN_2181 = 8'h2 < length_1 ? _GEN_2085 : _GEN_1989; // @[executor.scala 290:56]
  wire [7:0] _GEN_2182 = 8'h2 < length_1 ? _GEN_2086 : _GEN_1990; // @[executor.scala 290:56]
  wire [7:0] _GEN_2183 = 8'h2 < length_1 ? _GEN_2087 : _GEN_1991; // @[executor.scala 290:56]
  wire [7:0] _GEN_2184 = 8'h2 < length_1 ? _GEN_2088 : _GEN_1992; // @[executor.scala 290:56]
  wire [7:0] _GEN_2185 = 8'h2 < length_1 ? _GEN_2089 : _GEN_1993; // @[executor.scala 290:56]
  wire [7:0] _GEN_2186 = 8'h2 < length_1 ? _GEN_2090 : _GEN_1994; // @[executor.scala 290:56]
  wire [7:0] _GEN_2187 = 8'h2 < length_1 ? _GEN_2091 : _GEN_1995; // @[executor.scala 290:56]
  wire [7:0] _GEN_2188 = 8'h2 < length_1 ? _GEN_2092 : _GEN_1996; // @[executor.scala 290:56]
  wire [7:0] _GEN_2189 = 8'h2 < length_1 ? _GEN_2093 : _GEN_1997; // @[executor.scala 290:56]
  wire [7:0] _GEN_2190 = 8'h2 < length_1 ? _GEN_2094 : _GEN_1998; // @[executor.scala 290:56]
  wire [7:0] _GEN_2191 = 8'h2 < length_1 ? _GEN_2095 : _GEN_1999; // @[executor.scala 290:56]
  wire [7:0] _GEN_2192 = 8'h2 < length_1 ? _GEN_2096 : _GEN_2000; // @[executor.scala 290:56]
  wire [7:0] _GEN_2193 = 8'h2 < length_1 ? _GEN_2097 : _GEN_2001; // @[executor.scala 290:56]
  wire [7:0] _GEN_2194 = 8'h2 < length_1 ? _GEN_2098 : _GEN_2002; // @[executor.scala 290:56]
  wire [7:0] _GEN_2195 = 8'h2 < length_1 ? _GEN_2099 : _GEN_2003; // @[executor.scala 290:56]
  wire [7:0] _GEN_2196 = 8'h2 < length_1 ? _GEN_2100 : _GEN_2004; // @[executor.scala 290:56]
  wire [7:0] _GEN_2197 = 8'h2 < length_1 ? _GEN_2101 : _GEN_2005; // @[executor.scala 290:56]
  wire [7:0] _GEN_2198 = 8'h2 < length_1 ? _GEN_2102 : _GEN_2006; // @[executor.scala 290:56]
  wire [7:0] _GEN_2199 = 8'h2 < length_1 ? _GEN_2103 : _GEN_2007; // @[executor.scala 290:56]
  wire [7:0] _GEN_2200 = 8'h2 < length_1 ? _GEN_2104 : _GEN_2008; // @[executor.scala 290:56]
  wire [7:0] _GEN_2201 = 8'h2 < length_1 ? _GEN_2105 : _GEN_2009; // @[executor.scala 290:56]
  wire [7:0] _GEN_2202 = 8'h2 < length_1 ? _GEN_2106 : _GEN_2010; // @[executor.scala 290:56]
  wire [7:0] _GEN_2203 = 8'h2 < length_1 ? _GEN_2107 : _GEN_2011; // @[executor.scala 290:56]
  wire [7:0] _GEN_2204 = 8'h2 < length_1 ? _GEN_2108 : _GEN_2012; // @[executor.scala 290:56]
  wire [7:0] _GEN_2205 = 8'h2 < length_1 ? _GEN_2109 : _GEN_2013; // @[executor.scala 290:56]
  wire [7:0] _GEN_2206 = 8'h2 < length_1 ? _GEN_2110 : _GEN_2014; // @[executor.scala 290:56]
  wire [7:0] _GEN_2207 = 8'h2 < length_1 ? _GEN_2111 : _GEN_2015; // @[executor.scala 290:56]
  wire [7:0] _GEN_2208 = 8'h2 < length_1 ? _GEN_2112 : _GEN_2016; // @[executor.scala 290:56]
  wire [7:0] field_byte_11 = field_1[39:32]; // @[executor.scala 287:53]
  wire [7:0] total_offset_11 = offset_1 + 8'h3; // @[executor.scala 289:53]
  wire [7:0] _GEN_2209 = 7'h0 == total_offset_11[6:0] ? field_byte_11 : _GEN_2113; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2210 = 7'h1 == total_offset_11[6:0] ? field_byte_11 : _GEN_2114; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2211 = 7'h2 == total_offset_11[6:0] ? field_byte_11 : _GEN_2115; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2212 = 7'h3 == total_offset_11[6:0] ? field_byte_11 : _GEN_2116; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2213 = 7'h4 == total_offset_11[6:0] ? field_byte_11 : _GEN_2117; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2214 = 7'h5 == total_offset_11[6:0] ? field_byte_11 : _GEN_2118; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2215 = 7'h6 == total_offset_11[6:0] ? field_byte_11 : _GEN_2119; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2216 = 7'h7 == total_offset_11[6:0] ? field_byte_11 : _GEN_2120; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2217 = 7'h8 == total_offset_11[6:0] ? field_byte_11 : _GEN_2121; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2218 = 7'h9 == total_offset_11[6:0] ? field_byte_11 : _GEN_2122; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2219 = 7'ha == total_offset_11[6:0] ? field_byte_11 : _GEN_2123; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2220 = 7'hb == total_offset_11[6:0] ? field_byte_11 : _GEN_2124; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2221 = 7'hc == total_offset_11[6:0] ? field_byte_11 : _GEN_2125; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2222 = 7'hd == total_offset_11[6:0] ? field_byte_11 : _GEN_2126; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2223 = 7'he == total_offset_11[6:0] ? field_byte_11 : _GEN_2127; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2224 = 7'hf == total_offset_11[6:0] ? field_byte_11 : _GEN_2128; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2225 = 7'h10 == total_offset_11[6:0] ? field_byte_11 : _GEN_2129; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2226 = 7'h11 == total_offset_11[6:0] ? field_byte_11 : _GEN_2130; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2227 = 7'h12 == total_offset_11[6:0] ? field_byte_11 : _GEN_2131; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2228 = 7'h13 == total_offset_11[6:0] ? field_byte_11 : _GEN_2132; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2229 = 7'h14 == total_offset_11[6:0] ? field_byte_11 : _GEN_2133; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2230 = 7'h15 == total_offset_11[6:0] ? field_byte_11 : _GEN_2134; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2231 = 7'h16 == total_offset_11[6:0] ? field_byte_11 : _GEN_2135; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2232 = 7'h17 == total_offset_11[6:0] ? field_byte_11 : _GEN_2136; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2233 = 7'h18 == total_offset_11[6:0] ? field_byte_11 : _GEN_2137; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2234 = 7'h19 == total_offset_11[6:0] ? field_byte_11 : _GEN_2138; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2235 = 7'h1a == total_offset_11[6:0] ? field_byte_11 : _GEN_2139; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2236 = 7'h1b == total_offset_11[6:0] ? field_byte_11 : _GEN_2140; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2237 = 7'h1c == total_offset_11[6:0] ? field_byte_11 : _GEN_2141; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2238 = 7'h1d == total_offset_11[6:0] ? field_byte_11 : _GEN_2142; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2239 = 7'h1e == total_offset_11[6:0] ? field_byte_11 : _GEN_2143; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2240 = 7'h1f == total_offset_11[6:0] ? field_byte_11 : _GEN_2144; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2241 = 7'h20 == total_offset_11[6:0] ? field_byte_11 : _GEN_2145; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2242 = 7'h21 == total_offset_11[6:0] ? field_byte_11 : _GEN_2146; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2243 = 7'h22 == total_offset_11[6:0] ? field_byte_11 : _GEN_2147; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2244 = 7'h23 == total_offset_11[6:0] ? field_byte_11 : _GEN_2148; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2245 = 7'h24 == total_offset_11[6:0] ? field_byte_11 : _GEN_2149; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2246 = 7'h25 == total_offset_11[6:0] ? field_byte_11 : _GEN_2150; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2247 = 7'h26 == total_offset_11[6:0] ? field_byte_11 : _GEN_2151; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2248 = 7'h27 == total_offset_11[6:0] ? field_byte_11 : _GEN_2152; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2249 = 7'h28 == total_offset_11[6:0] ? field_byte_11 : _GEN_2153; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2250 = 7'h29 == total_offset_11[6:0] ? field_byte_11 : _GEN_2154; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2251 = 7'h2a == total_offset_11[6:0] ? field_byte_11 : _GEN_2155; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2252 = 7'h2b == total_offset_11[6:0] ? field_byte_11 : _GEN_2156; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2253 = 7'h2c == total_offset_11[6:0] ? field_byte_11 : _GEN_2157; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2254 = 7'h2d == total_offset_11[6:0] ? field_byte_11 : _GEN_2158; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2255 = 7'h2e == total_offset_11[6:0] ? field_byte_11 : _GEN_2159; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2256 = 7'h2f == total_offset_11[6:0] ? field_byte_11 : _GEN_2160; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2257 = 7'h30 == total_offset_11[6:0] ? field_byte_11 : _GEN_2161; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2258 = 7'h31 == total_offset_11[6:0] ? field_byte_11 : _GEN_2162; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2259 = 7'h32 == total_offset_11[6:0] ? field_byte_11 : _GEN_2163; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2260 = 7'h33 == total_offset_11[6:0] ? field_byte_11 : _GEN_2164; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2261 = 7'h34 == total_offset_11[6:0] ? field_byte_11 : _GEN_2165; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2262 = 7'h35 == total_offset_11[6:0] ? field_byte_11 : _GEN_2166; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2263 = 7'h36 == total_offset_11[6:0] ? field_byte_11 : _GEN_2167; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2264 = 7'h37 == total_offset_11[6:0] ? field_byte_11 : _GEN_2168; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2265 = 7'h38 == total_offset_11[6:0] ? field_byte_11 : _GEN_2169; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2266 = 7'h39 == total_offset_11[6:0] ? field_byte_11 : _GEN_2170; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2267 = 7'h3a == total_offset_11[6:0] ? field_byte_11 : _GEN_2171; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2268 = 7'h3b == total_offset_11[6:0] ? field_byte_11 : _GEN_2172; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2269 = 7'h3c == total_offset_11[6:0] ? field_byte_11 : _GEN_2173; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2270 = 7'h3d == total_offset_11[6:0] ? field_byte_11 : _GEN_2174; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2271 = 7'h3e == total_offset_11[6:0] ? field_byte_11 : _GEN_2175; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2272 = 7'h3f == total_offset_11[6:0] ? field_byte_11 : _GEN_2176; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2273 = 7'h40 == total_offset_11[6:0] ? field_byte_11 : _GEN_2177; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2274 = 7'h41 == total_offset_11[6:0] ? field_byte_11 : _GEN_2178; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2275 = 7'h42 == total_offset_11[6:0] ? field_byte_11 : _GEN_2179; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2276 = 7'h43 == total_offset_11[6:0] ? field_byte_11 : _GEN_2180; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2277 = 7'h44 == total_offset_11[6:0] ? field_byte_11 : _GEN_2181; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2278 = 7'h45 == total_offset_11[6:0] ? field_byte_11 : _GEN_2182; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2279 = 7'h46 == total_offset_11[6:0] ? field_byte_11 : _GEN_2183; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2280 = 7'h47 == total_offset_11[6:0] ? field_byte_11 : _GEN_2184; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2281 = 7'h48 == total_offset_11[6:0] ? field_byte_11 : _GEN_2185; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2282 = 7'h49 == total_offset_11[6:0] ? field_byte_11 : _GEN_2186; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2283 = 7'h4a == total_offset_11[6:0] ? field_byte_11 : _GEN_2187; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2284 = 7'h4b == total_offset_11[6:0] ? field_byte_11 : _GEN_2188; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2285 = 7'h4c == total_offset_11[6:0] ? field_byte_11 : _GEN_2189; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2286 = 7'h4d == total_offset_11[6:0] ? field_byte_11 : _GEN_2190; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2287 = 7'h4e == total_offset_11[6:0] ? field_byte_11 : _GEN_2191; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2288 = 7'h4f == total_offset_11[6:0] ? field_byte_11 : _GEN_2192; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2289 = 7'h50 == total_offset_11[6:0] ? field_byte_11 : _GEN_2193; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2290 = 7'h51 == total_offset_11[6:0] ? field_byte_11 : _GEN_2194; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2291 = 7'h52 == total_offset_11[6:0] ? field_byte_11 : _GEN_2195; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2292 = 7'h53 == total_offset_11[6:0] ? field_byte_11 : _GEN_2196; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2293 = 7'h54 == total_offset_11[6:0] ? field_byte_11 : _GEN_2197; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2294 = 7'h55 == total_offset_11[6:0] ? field_byte_11 : _GEN_2198; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2295 = 7'h56 == total_offset_11[6:0] ? field_byte_11 : _GEN_2199; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2296 = 7'h57 == total_offset_11[6:0] ? field_byte_11 : _GEN_2200; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2297 = 7'h58 == total_offset_11[6:0] ? field_byte_11 : _GEN_2201; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2298 = 7'h59 == total_offset_11[6:0] ? field_byte_11 : _GEN_2202; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2299 = 7'h5a == total_offset_11[6:0] ? field_byte_11 : _GEN_2203; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2300 = 7'h5b == total_offset_11[6:0] ? field_byte_11 : _GEN_2204; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2301 = 7'h5c == total_offset_11[6:0] ? field_byte_11 : _GEN_2205; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2302 = 7'h5d == total_offset_11[6:0] ? field_byte_11 : _GEN_2206; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2303 = 7'h5e == total_offset_11[6:0] ? field_byte_11 : _GEN_2207; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2304 = 7'h5f == total_offset_11[6:0] ? field_byte_11 : _GEN_2208; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2305 = 8'h3 < length_1 ? _GEN_2209 : _GEN_2113; // @[executor.scala 290:56]
  wire [7:0] _GEN_2306 = 8'h3 < length_1 ? _GEN_2210 : _GEN_2114; // @[executor.scala 290:56]
  wire [7:0] _GEN_2307 = 8'h3 < length_1 ? _GEN_2211 : _GEN_2115; // @[executor.scala 290:56]
  wire [7:0] _GEN_2308 = 8'h3 < length_1 ? _GEN_2212 : _GEN_2116; // @[executor.scala 290:56]
  wire [7:0] _GEN_2309 = 8'h3 < length_1 ? _GEN_2213 : _GEN_2117; // @[executor.scala 290:56]
  wire [7:0] _GEN_2310 = 8'h3 < length_1 ? _GEN_2214 : _GEN_2118; // @[executor.scala 290:56]
  wire [7:0] _GEN_2311 = 8'h3 < length_1 ? _GEN_2215 : _GEN_2119; // @[executor.scala 290:56]
  wire [7:0] _GEN_2312 = 8'h3 < length_1 ? _GEN_2216 : _GEN_2120; // @[executor.scala 290:56]
  wire [7:0] _GEN_2313 = 8'h3 < length_1 ? _GEN_2217 : _GEN_2121; // @[executor.scala 290:56]
  wire [7:0] _GEN_2314 = 8'h3 < length_1 ? _GEN_2218 : _GEN_2122; // @[executor.scala 290:56]
  wire [7:0] _GEN_2315 = 8'h3 < length_1 ? _GEN_2219 : _GEN_2123; // @[executor.scala 290:56]
  wire [7:0] _GEN_2316 = 8'h3 < length_1 ? _GEN_2220 : _GEN_2124; // @[executor.scala 290:56]
  wire [7:0] _GEN_2317 = 8'h3 < length_1 ? _GEN_2221 : _GEN_2125; // @[executor.scala 290:56]
  wire [7:0] _GEN_2318 = 8'h3 < length_1 ? _GEN_2222 : _GEN_2126; // @[executor.scala 290:56]
  wire [7:0] _GEN_2319 = 8'h3 < length_1 ? _GEN_2223 : _GEN_2127; // @[executor.scala 290:56]
  wire [7:0] _GEN_2320 = 8'h3 < length_1 ? _GEN_2224 : _GEN_2128; // @[executor.scala 290:56]
  wire [7:0] _GEN_2321 = 8'h3 < length_1 ? _GEN_2225 : _GEN_2129; // @[executor.scala 290:56]
  wire [7:0] _GEN_2322 = 8'h3 < length_1 ? _GEN_2226 : _GEN_2130; // @[executor.scala 290:56]
  wire [7:0] _GEN_2323 = 8'h3 < length_1 ? _GEN_2227 : _GEN_2131; // @[executor.scala 290:56]
  wire [7:0] _GEN_2324 = 8'h3 < length_1 ? _GEN_2228 : _GEN_2132; // @[executor.scala 290:56]
  wire [7:0] _GEN_2325 = 8'h3 < length_1 ? _GEN_2229 : _GEN_2133; // @[executor.scala 290:56]
  wire [7:0] _GEN_2326 = 8'h3 < length_1 ? _GEN_2230 : _GEN_2134; // @[executor.scala 290:56]
  wire [7:0] _GEN_2327 = 8'h3 < length_1 ? _GEN_2231 : _GEN_2135; // @[executor.scala 290:56]
  wire [7:0] _GEN_2328 = 8'h3 < length_1 ? _GEN_2232 : _GEN_2136; // @[executor.scala 290:56]
  wire [7:0] _GEN_2329 = 8'h3 < length_1 ? _GEN_2233 : _GEN_2137; // @[executor.scala 290:56]
  wire [7:0] _GEN_2330 = 8'h3 < length_1 ? _GEN_2234 : _GEN_2138; // @[executor.scala 290:56]
  wire [7:0] _GEN_2331 = 8'h3 < length_1 ? _GEN_2235 : _GEN_2139; // @[executor.scala 290:56]
  wire [7:0] _GEN_2332 = 8'h3 < length_1 ? _GEN_2236 : _GEN_2140; // @[executor.scala 290:56]
  wire [7:0] _GEN_2333 = 8'h3 < length_1 ? _GEN_2237 : _GEN_2141; // @[executor.scala 290:56]
  wire [7:0] _GEN_2334 = 8'h3 < length_1 ? _GEN_2238 : _GEN_2142; // @[executor.scala 290:56]
  wire [7:0] _GEN_2335 = 8'h3 < length_1 ? _GEN_2239 : _GEN_2143; // @[executor.scala 290:56]
  wire [7:0] _GEN_2336 = 8'h3 < length_1 ? _GEN_2240 : _GEN_2144; // @[executor.scala 290:56]
  wire [7:0] _GEN_2337 = 8'h3 < length_1 ? _GEN_2241 : _GEN_2145; // @[executor.scala 290:56]
  wire [7:0] _GEN_2338 = 8'h3 < length_1 ? _GEN_2242 : _GEN_2146; // @[executor.scala 290:56]
  wire [7:0] _GEN_2339 = 8'h3 < length_1 ? _GEN_2243 : _GEN_2147; // @[executor.scala 290:56]
  wire [7:0] _GEN_2340 = 8'h3 < length_1 ? _GEN_2244 : _GEN_2148; // @[executor.scala 290:56]
  wire [7:0] _GEN_2341 = 8'h3 < length_1 ? _GEN_2245 : _GEN_2149; // @[executor.scala 290:56]
  wire [7:0] _GEN_2342 = 8'h3 < length_1 ? _GEN_2246 : _GEN_2150; // @[executor.scala 290:56]
  wire [7:0] _GEN_2343 = 8'h3 < length_1 ? _GEN_2247 : _GEN_2151; // @[executor.scala 290:56]
  wire [7:0] _GEN_2344 = 8'h3 < length_1 ? _GEN_2248 : _GEN_2152; // @[executor.scala 290:56]
  wire [7:0] _GEN_2345 = 8'h3 < length_1 ? _GEN_2249 : _GEN_2153; // @[executor.scala 290:56]
  wire [7:0] _GEN_2346 = 8'h3 < length_1 ? _GEN_2250 : _GEN_2154; // @[executor.scala 290:56]
  wire [7:0] _GEN_2347 = 8'h3 < length_1 ? _GEN_2251 : _GEN_2155; // @[executor.scala 290:56]
  wire [7:0] _GEN_2348 = 8'h3 < length_1 ? _GEN_2252 : _GEN_2156; // @[executor.scala 290:56]
  wire [7:0] _GEN_2349 = 8'h3 < length_1 ? _GEN_2253 : _GEN_2157; // @[executor.scala 290:56]
  wire [7:0] _GEN_2350 = 8'h3 < length_1 ? _GEN_2254 : _GEN_2158; // @[executor.scala 290:56]
  wire [7:0] _GEN_2351 = 8'h3 < length_1 ? _GEN_2255 : _GEN_2159; // @[executor.scala 290:56]
  wire [7:0] _GEN_2352 = 8'h3 < length_1 ? _GEN_2256 : _GEN_2160; // @[executor.scala 290:56]
  wire [7:0] _GEN_2353 = 8'h3 < length_1 ? _GEN_2257 : _GEN_2161; // @[executor.scala 290:56]
  wire [7:0] _GEN_2354 = 8'h3 < length_1 ? _GEN_2258 : _GEN_2162; // @[executor.scala 290:56]
  wire [7:0] _GEN_2355 = 8'h3 < length_1 ? _GEN_2259 : _GEN_2163; // @[executor.scala 290:56]
  wire [7:0] _GEN_2356 = 8'h3 < length_1 ? _GEN_2260 : _GEN_2164; // @[executor.scala 290:56]
  wire [7:0] _GEN_2357 = 8'h3 < length_1 ? _GEN_2261 : _GEN_2165; // @[executor.scala 290:56]
  wire [7:0] _GEN_2358 = 8'h3 < length_1 ? _GEN_2262 : _GEN_2166; // @[executor.scala 290:56]
  wire [7:0] _GEN_2359 = 8'h3 < length_1 ? _GEN_2263 : _GEN_2167; // @[executor.scala 290:56]
  wire [7:0] _GEN_2360 = 8'h3 < length_1 ? _GEN_2264 : _GEN_2168; // @[executor.scala 290:56]
  wire [7:0] _GEN_2361 = 8'h3 < length_1 ? _GEN_2265 : _GEN_2169; // @[executor.scala 290:56]
  wire [7:0] _GEN_2362 = 8'h3 < length_1 ? _GEN_2266 : _GEN_2170; // @[executor.scala 290:56]
  wire [7:0] _GEN_2363 = 8'h3 < length_1 ? _GEN_2267 : _GEN_2171; // @[executor.scala 290:56]
  wire [7:0] _GEN_2364 = 8'h3 < length_1 ? _GEN_2268 : _GEN_2172; // @[executor.scala 290:56]
  wire [7:0] _GEN_2365 = 8'h3 < length_1 ? _GEN_2269 : _GEN_2173; // @[executor.scala 290:56]
  wire [7:0] _GEN_2366 = 8'h3 < length_1 ? _GEN_2270 : _GEN_2174; // @[executor.scala 290:56]
  wire [7:0] _GEN_2367 = 8'h3 < length_1 ? _GEN_2271 : _GEN_2175; // @[executor.scala 290:56]
  wire [7:0] _GEN_2368 = 8'h3 < length_1 ? _GEN_2272 : _GEN_2176; // @[executor.scala 290:56]
  wire [7:0] _GEN_2369 = 8'h3 < length_1 ? _GEN_2273 : _GEN_2177; // @[executor.scala 290:56]
  wire [7:0] _GEN_2370 = 8'h3 < length_1 ? _GEN_2274 : _GEN_2178; // @[executor.scala 290:56]
  wire [7:0] _GEN_2371 = 8'h3 < length_1 ? _GEN_2275 : _GEN_2179; // @[executor.scala 290:56]
  wire [7:0] _GEN_2372 = 8'h3 < length_1 ? _GEN_2276 : _GEN_2180; // @[executor.scala 290:56]
  wire [7:0] _GEN_2373 = 8'h3 < length_1 ? _GEN_2277 : _GEN_2181; // @[executor.scala 290:56]
  wire [7:0] _GEN_2374 = 8'h3 < length_1 ? _GEN_2278 : _GEN_2182; // @[executor.scala 290:56]
  wire [7:0] _GEN_2375 = 8'h3 < length_1 ? _GEN_2279 : _GEN_2183; // @[executor.scala 290:56]
  wire [7:0] _GEN_2376 = 8'h3 < length_1 ? _GEN_2280 : _GEN_2184; // @[executor.scala 290:56]
  wire [7:0] _GEN_2377 = 8'h3 < length_1 ? _GEN_2281 : _GEN_2185; // @[executor.scala 290:56]
  wire [7:0] _GEN_2378 = 8'h3 < length_1 ? _GEN_2282 : _GEN_2186; // @[executor.scala 290:56]
  wire [7:0] _GEN_2379 = 8'h3 < length_1 ? _GEN_2283 : _GEN_2187; // @[executor.scala 290:56]
  wire [7:0] _GEN_2380 = 8'h3 < length_1 ? _GEN_2284 : _GEN_2188; // @[executor.scala 290:56]
  wire [7:0] _GEN_2381 = 8'h3 < length_1 ? _GEN_2285 : _GEN_2189; // @[executor.scala 290:56]
  wire [7:0] _GEN_2382 = 8'h3 < length_1 ? _GEN_2286 : _GEN_2190; // @[executor.scala 290:56]
  wire [7:0] _GEN_2383 = 8'h3 < length_1 ? _GEN_2287 : _GEN_2191; // @[executor.scala 290:56]
  wire [7:0] _GEN_2384 = 8'h3 < length_1 ? _GEN_2288 : _GEN_2192; // @[executor.scala 290:56]
  wire [7:0] _GEN_2385 = 8'h3 < length_1 ? _GEN_2289 : _GEN_2193; // @[executor.scala 290:56]
  wire [7:0] _GEN_2386 = 8'h3 < length_1 ? _GEN_2290 : _GEN_2194; // @[executor.scala 290:56]
  wire [7:0] _GEN_2387 = 8'h3 < length_1 ? _GEN_2291 : _GEN_2195; // @[executor.scala 290:56]
  wire [7:0] _GEN_2388 = 8'h3 < length_1 ? _GEN_2292 : _GEN_2196; // @[executor.scala 290:56]
  wire [7:0] _GEN_2389 = 8'h3 < length_1 ? _GEN_2293 : _GEN_2197; // @[executor.scala 290:56]
  wire [7:0] _GEN_2390 = 8'h3 < length_1 ? _GEN_2294 : _GEN_2198; // @[executor.scala 290:56]
  wire [7:0] _GEN_2391 = 8'h3 < length_1 ? _GEN_2295 : _GEN_2199; // @[executor.scala 290:56]
  wire [7:0] _GEN_2392 = 8'h3 < length_1 ? _GEN_2296 : _GEN_2200; // @[executor.scala 290:56]
  wire [7:0] _GEN_2393 = 8'h3 < length_1 ? _GEN_2297 : _GEN_2201; // @[executor.scala 290:56]
  wire [7:0] _GEN_2394 = 8'h3 < length_1 ? _GEN_2298 : _GEN_2202; // @[executor.scala 290:56]
  wire [7:0] _GEN_2395 = 8'h3 < length_1 ? _GEN_2299 : _GEN_2203; // @[executor.scala 290:56]
  wire [7:0] _GEN_2396 = 8'h3 < length_1 ? _GEN_2300 : _GEN_2204; // @[executor.scala 290:56]
  wire [7:0] _GEN_2397 = 8'h3 < length_1 ? _GEN_2301 : _GEN_2205; // @[executor.scala 290:56]
  wire [7:0] _GEN_2398 = 8'h3 < length_1 ? _GEN_2302 : _GEN_2206; // @[executor.scala 290:56]
  wire [7:0] _GEN_2399 = 8'h3 < length_1 ? _GEN_2303 : _GEN_2207; // @[executor.scala 290:56]
  wire [7:0] _GEN_2400 = 8'h3 < length_1 ? _GEN_2304 : _GEN_2208; // @[executor.scala 290:56]
  wire [7:0] field_byte_12 = field_1[31:24]; // @[executor.scala 287:53]
  wire [7:0] total_offset_12 = offset_1 + 8'h4; // @[executor.scala 289:53]
  wire [7:0] _GEN_2401 = 7'h0 == total_offset_12[6:0] ? field_byte_12 : _GEN_2305; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2402 = 7'h1 == total_offset_12[6:0] ? field_byte_12 : _GEN_2306; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2403 = 7'h2 == total_offset_12[6:0] ? field_byte_12 : _GEN_2307; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2404 = 7'h3 == total_offset_12[6:0] ? field_byte_12 : _GEN_2308; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2405 = 7'h4 == total_offset_12[6:0] ? field_byte_12 : _GEN_2309; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2406 = 7'h5 == total_offset_12[6:0] ? field_byte_12 : _GEN_2310; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2407 = 7'h6 == total_offset_12[6:0] ? field_byte_12 : _GEN_2311; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2408 = 7'h7 == total_offset_12[6:0] ? field_byte_12 : _GEN_2312; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2409 = 7'h8 == total_offset_12[6:0] ? field_byte_12 : _GEN_2313; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2410 = 7'h9 == total_offset_12[6:0] ? field_byte_12 : _GEN_2314; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2411 = 7'ha == total_offset_12[6:0] ? field_byte_12 : _GEN_2315; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2412 = 7'hb == total_offset_12[6:0] ? field_byte_12 : _GEN_2316; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2413 = 7'hc == total_offset_12[6:0] ? field_byte_12 : _GEN_2317; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2414 = 7'hd == total_offset_12[6:0] ? field_byte_12 : _GEN_2318; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2415 = 7'he == total_offset_12[6:0] ? field_byte_12 : _GEN_2319; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2416 = 7'hf == total_offset_12[6:0] ? field_byte_12 : _GEN_2320; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2417 = 7'h10 == total_offset_12[6:0] ? field_byte_12 : _GEN_2321; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2418 = 7'h11 == total_offset_12[6:0] ? field_byte_12 : _GEN_2322; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2419 = 7'h12 == total_offset_12[6:0] ? field_byte_12 : _GEN_2323; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2420 = 7'h13 == total_offset_12[6:0] ? field_byte_12 : _GEN_2324; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2421 = 7'h14 == total_offset_12[6:0] ? field_byte_12 : _GEN_2325; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2422 = 7'h15 == total_offset_12[6:0] ? field_byte_12 : _GEN_2326; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2423 = 7'h16 == total_offset_12[6:0] ? field_byte_12 : _GEN_2327; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2424 = 7'h17 == total_offset_12[6:0] ? field_byte_12 : _GEN_2328; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2425 = 7'h18 == total_offset_12[6:0] ? field_byte_12 : _GEN_2329; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2426 = 7'h19 == total_offset_12[6:0] ? field_byte_12 : _GEN_2330; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2427 = 7'h1a == total_offset_12[6:0] ? field_byte_12 : _GEN_2331; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2428 = 7'h1b == total_offset_12[6:0] ? field_byte_12 : _GEN_2332; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2429 = 7'h1c == total_offset_12[6:0] ? field_byte_12 : _GEN_2333; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2430 = 7'h1d == total_offset_12[6:0] ? field_byte_12 : _GEN_2334; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2431 = 7'h1e == total_offset_12[6:0] ? field_byte_12 : _GEN_2335; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2432 = 7'h1f == total_offset_12[6:0] ? field_byte_12 : _GEN_2336; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2433 = 7'h20 == total_offset_12[6:0] ? field_byte_12 : _GEN_2337; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2434 = 7'h21 == total_offset_12[6:0] ? field_byte_12 : _GEN_2338; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2435 = 7'h22 == total_offset_12[6:0] ? field_byte_12 : _GEN_2339; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2436 = 7'h23 == total_offset_12[6:0] ? field_byte_12 : _GEN_2340; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2437 = 7'h24 == total_offset_12[6:0] ? field_byte_12 : _GEN_2341; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2438 = 7'h25 == total_offset_12[6:0] ? field_byte_12 : _GEN_2342; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2439 = 7'h26 == total_offset_12[6:0] ? field_byte_12 : _GEN_2343; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2440 = 7'h27 == total_offset_12[6:0] ? field_byte_12 : _GEN_2344; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2441 = 7'h28 == total_offset_12[6:0] ? field_byte_12 : _GEN_2345; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2442 = 7'h29 == total_offset_12[6:0] ? field_byte_12 : _GEN_2346; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2443 = 7'h2a == total_offset_12[6:0] ? field_byte_12 : _GEN_2347; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2444 = 7'h2b == total_offset_12[6:0] ? field_byte_12 : _GEN_2348; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2445 = 7'h2c == total_offset_12[6:0] ? field_byte_12 : _GEN_2349; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2446 = 7'h2d == total_offset_12[6:0] ? field_byte_12 : _GEN_2350; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2447 = 7'h2e == total_offset_12[6:0] ? field_byte_12 : _GEN_2351; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2448 = 7'h2f == total_offset_12[6:0] ? field_byte_12 : _GEN_2352; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2449 = 7'h30 == total_offset_12[6:0] ? field_byte_12 : _GEN_2353; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2450 = 7'h31 == total_offset_12[6:0] ? field_byte_12 : _GEN_2354; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2451 = 7'h32 == total_offset_12[6:0] ? field_byte_12 : _GEN_2355; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2452 = 7'h33 == total_offset_12[6:0] ? field_byte_12 : _GEN_2356; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2453 = 7'h34 == total_offset_12[6:0] ? field_byte_12 : _GEN_2357; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2454 = 7'h35 == total_offset_12[6:0] ? field_byte_12 : _GEN_2358; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2455 = 7'h36 == total_offset_12[6:0] ? field_byte_12 : _GEN_2359; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2456 = 7'h37 == total_offset_12[6:0] ? field_byte_12 : _GEN_2360; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2457 = 7'h38 == total_offset_12[6:0] ? field_byte_12 : _GEN_2361; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2458 = 7'h39 == total_offset_12[6:0] ? field_byte_12 : _GEN_2362; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2459 = 7'h3a == total_offset_12[6:0] ? field_byte_12 : _GEN_2363; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2460 = 7'h3b == total_offset_12[6:0] ? field_byte_12 : _GEN_2364; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2461 = 7'h3c == total_offset_12[6:0] ? field_byte_12 : _GEN_2365; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2462 = 7'h3d == total_offset_12[6:0] ? field_byte_12 : _GEN_2366; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2463 = 7'h3e == total_offset_12[6:0] ? field_byte_12 : _GEN_2367; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2464 = 7'h3f == total_offset_12[6:0] ? field_byte_12 : _GEN_2368; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2465 = 7'h40 == total_offset_12[6:0] ? field_byte_12 : _GEN_2369; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2466 = 7'h41 == total_offset_12[6:0] ? field_byte_12 : _GEN_2370; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2467 = 7'h42 == total_offset_12[6:0] ? field_byte_12 : _GEN_2371; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2468 = 7'h43 == total_offset_12[6:0] ? field_byte_12 : _GEN_2372; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2469 = 7'h44 == total_offset_12[6:0] ? field_byte_12 : _GEN_2373; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2470 = 7'h45 == total_offset_12[6:0] ? field_byte_12 : _GEN_2374; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2471 = 7'h46 == total_offset_12[6:0] ? field_byte_12 : _GEN_2375; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2472 = 7'h47 == total_offset_12[6:0] ? field_byte_12 : _GEN_2376; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2473 = 7'h48 == total_offset_12[6:0] ? field_byte_12 : _GEN_2377; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2474 = 7'h49 == total_offset_12[6:0] ? field_byte_12 : _GEN_2378; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2475 = 7'h4a == total_offset_12[6:0] ? field_byte_12 : _GEN_2379; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2476 = 7'h4b == total_offset_12[6:0] ? field_byte_12 : _GEN_2380; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2477 = 7'h4c == total_offset_12[6:0] ? field_byte_12 : _GEN_2381; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2478 = 7'h4d == total_offset_12[6:0] ? field_byte_12 : _GEN_2382; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2479 = 7'h4e == total_offset_12[6:0] ? field_byte_12 : _GEN_2383; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2480 = 7'h4f == total_offset_12[6:0] ? field_byte_12 : _GEN_2384; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2481 = 7'h50 == total_offset_12[6:0] ? field_byte_12 : _GEN_2385; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2482 = 7'h51 == total_offset_12[6:0] ? field_byte_12 : _GEN_2386; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2483 = 7'h52 == total_offset_12[6:0] ? field_byte_12 : _GEN_2387; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2484 = 7'h53 == total_offset_12[6:0] ? field_byte_12 : _GEN_2388; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2485 = 7'h54 == total_offset_12[6:0] ? field_byte_12 : _GEN_2389; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2486 = 7'h55 == total_offset_12[6:0] ? field_byte_12 : _GEN_2390; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2487 = 7'h56 == total_offset_12[6:0] ? field_byte_12 : _GEN_2391; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2488 = 7'h57 == total_offset_12[6:0] ? field_byte_12 : _GEN_2392; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2489 = 7'h58 == total_offset_12[6:0] ? field_byte_12 : _GEN_2393; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2490 = 7'h59 == total_offset_12[6:0] ? field_byte_12 : _GEN_2394; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2491 = 7'h5a == total_offset_12[6:0] ? field_byte_12 : _GEN_2395; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2492 = 7'h5b == total_offset_12[6:0] ? field_byte_12 : _GEN_2396; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2493 = 7'h5c == total_offset_12[6:0] ? field_byte_12 : _GEN_2397; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2494 = 7'h5d == total_offset_12[6:0] ? field_byte_12 : _GEN_2398; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2495 = 7'h5e == total_offset_12[6:0] ? field_byte_12 : _GEN_2399; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2496 = 7'h5f == total_offset_12[6:0] ? field_byte_12 : _GEN_2400; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2497 = 8'h4 < length_1 ? _GEN_2401 : _GEN_2305; // @[executor.scala 290:56]
  wire [7:0] _GEN_2498 = 8'h4 < length_1 ? _GEN_2402 : _GEN_2306; // @[executor.scala 290:56]
  wire [7:0] _GEN_2499 = 8'h4 < length_1 ? _GEN_2403 : _GEN_2307; // @[executor.scala 290:56]
  wire [7:0] _GEN_2500 = 8'h4 < length_1 ? _GEN_2404 : _GEN_2308; // @[executor.scala 290:56]
  wire [7:0] _GEN_2501 = 8'h4 < length_1 ? _GEN_2405 : _GEN_2309; // @[executor.scala 290:56]
  wire [7:0] _GEN_2502 = 8'h4 < length_1 ? _GEN_2406 : _GEN_2310; // @[executor.scala 290:56]
  wire [7:0] _GEN_2503 = 8'h4 < length_1 ? _GEN_2407 : _GEN_2311; // @[executor.scala 290:56]
  wire [7:0] _GEN_2504 = 8'h4 < length_1 ? _GEN_2408 : _GEN_2312; // @[executor.scala 290:56]
  wire [7:0] _GEN_2505 = 8'h4 < length_1 ? _GEN_2409 : _GEN_2313; // @[executor.scala 290:56]
  wire [7:0] _GEN_2506 = 8'h4 < length_1 ? _GEN_2410 : _GEN_2314; // @[executor.scala 290:56]
  wire [7:0] _GEN_2507 = 8'h4 < length_1 ? _GEN_2411 : _GEN_2315; // @[executor.scala 290:56]
  wire [7:0] _GEN_2508 = 8'h4 < length_1 ? _GEN_2412 : _GEN_2316; // @[executor.scala 290:56]
  wire [7:0] _GEN_2509 = 8'h4 < length_1 ? _GEN_2413 : _GEN_2317; // @[executor.scala 290:56]
  wire [7:0] _GEN_2510 = 8'h4 < length_1 ? _GEN_2414 : _GEN_2318; // @[executor.scala 290:56]
  wire [7:0] _GEN_2511 = 8'h4 < length_1 ? _GEN_2415 : _GEN_2319; // @[executor.scala 290:56]
  wire [7:0] _GEN_2512 = 8'h4 < length_1 ? _GEN_2416 : _GEN_2320; // @[executor.scala 290:56]
  wire [7:0] _GEN_2513 = 8'h4 < length_1 ? _GEN_2417 : _GEN_2321; // @[executor.scala 290:56]
  wire [7:0] _GEN_2514 = 8'h4 < length_1 ? _GEN_2418 : _GEN_2322; // @[executor.scala 290:56]
  wire [7:0] _GEN_2515 = 8'h4 < length_1 ? _GEN_2419 : _GEN_2323; // @[executor.scala 290:56]
  wire [7:0] _GEN_2516 = 8'h4 < length_1 ? _GEN_2420 : _GEN_2324; // @[executor.scala 290:56]
  wire [7:0] _GEN_2517 = 8'h4 < length_1 ? _GEN_2421 : _GEN_2325; // @[executor.scala 290:56]
  wire [7:0] _GEN_2518 = 8'h4 < length_1 ? _GEN_2422 : _GEN_2326; // @[executor.scala 290:56]
  wire [7:0] _GEN_2519 = 8'h4 < length_1 ? _GEN_2423 : _GEN_2327; // @[executor.scala 290:56]
  wire [7:0] _GEN_2520 = 8'h4 < length_1 ? _GEN_2424 : _GEN_2328; // @[executor.scala 290:56]
  wire [7:0] _GEN_2521 = 8'h4 < length_1 ? _GEN_2425 : _GEN_2329; // @[executor.scala 290:56]
  wire [7:0] _GEN_2522 = 8'h4 < length_1 ? _GEN_2426 : _GEN_2330; // @[executor.scala 290:56]
  wire [7:0] _GEN_2523 = 8'h4 < length_1 ? _GEN_2427 : _GEN_2331; // @[executor.scala 290:56]
  wire [7:0] _GEN_2524 = 8'h4 < length_1 ? _GEN_2428 : _GEN_2332; // @[executor.scala 290:56]
  wire [7:0] _GEN_2525 = 8'h4 < length_1 ? _GEN_2429 : _GEN_2333; // @[executor.scala 290:56]
  wire [7:0] _GEN_2526 = 8'h4 < length_1 ? _GEN_2430 : _GEN_2334; // @[executor.scala 290:56]
  wire [7:0] _GEN_2527 = 8'h4 < length_1 ? _GEN_2431 : _GEN_2335; // @[executor.scala 290:56]
  wire [7:0] _GEN_2528 = 8'h4 < length_1 ? _GEN_2432 : _GEN_2336; // @[executor.scala 290:56]
  wire [7:0] _GEN_2529 = 8'h4 < length_1 ? _GEN_2433 : _GEN_2337; // @[executor.scala 290:56]
  wire [7:0] _GEN_2530 = 8'h4 < length_1 ? _GEN_2434 : _GEN_2338; // @[executor.scala 290:56]
  wire [7:0] _GEN_2531 = 8'h4 < length_1 ? _GEN_2435 : _GEN_2339; // @[executor.scala 290:56]
  wire [7:0] _GEN_2532 = 8'h4 < length_1 ? _GEN_2436 : _GEN_2340; // @[executor.scala 290:56]
  wire [7:0] _GEN_2533 = 8'h4 < length_1 ? _GEN_2437 : _GEN_2341; // @[executor.scala 290:56]
  wire [7:0] _GEN_2534 = 8'h4 < length_1 ? _GEN_2438 : _GEN_2342; // @[executor.scala 290:56]
  wire [7:0] _GEN_2535 = 8'h4 < length_1 ? _GEN_2439 : _GEN_2343; // @[executor.scala 290:56]
  wire [7:0] _GEN_2536 = 8'h4 < length_1 ? _GEN_2440 : _GEN_2344; // @[executor.scala 290:56]
  wire [7:0] _GEN_2537 = 8'h4 < length_1 ? _GEN_2441 : _GEN_2345; // @[executor.scala 290:56]
  wire [7:0] _GEN_2538 = 8'h4 < length_1 ? _GEN_2442 : _GEN_2346; // @[executor.scala 290:56]
  wire [7:0] _GEN_2539 = 8'h4 < length_1 ? _GEN_2443 : _GEN_2347; // @[executor.scala 290:56]
  wire [7:0] _GEN_2540 = 8'h4 < length_1 ? _GEN_2444 : _GEN_2348; // @[executor.scala 290:56]
  wire [7:0] _GEN_2541 = 8'h4 < length_1 ? _GEN_2445 : _GEN_2349; // @[executor.scala 290:56]
  wire [7:0] _GEN_2542 = 8'h4 < length_1 ? _GEN_2446 : _GEN_2350; // @[executor.scala 290:56]
  wire [7:0] _GEN_2543 = 8'h4 < length_1 ? _GEN_2447 : _GEN_2351; // @[executor.scala 290:56]
  wire [7:0] _GEN_2544 = 8'h4 < length_1 ? _GEN_2448 : _GEN_2352; // @[executor.scala 290:56]
  wire [7:0] _GEN_2545 = 8'h4 < length_1 ? _GEN_2449 : _GEN_2353; // @[executor.scala 290:56]
  wire [7:0] _GEN_2546 = 8'h4 < length_1 ? _GEN_2450 : _GEN_2354; // @[executor.scala 290:56]
  wire [7:0] _GEN_2547 = 8'h4 < length_1 ? _GEN_2451 : _GEN_2355; // @[executor.scala 290:56]
  wire [7:0] _GEN_2548 = 8'h4 < length_1 ? _GEN_2452 : _GEN_2356; // @[executor.scala 290:56]
  wire [7:0] _GEN_2549 = 8'h4 < length_1 ? _GEN_2453 : _GEN_2357; // @[executor.scala 290:56]
  wire [7:0] _GEN_2550 = 8'h4 < length_1 ? _GEN_2454 : _GEN_2358; // @[executor.scala 290:56]
  wire [7:0] _GEN_2551 = 8'h4 < length_1 ? _GEN_2455 : _GEN_2359; // @[executor.scala 290:56]
  wire [7:0] _GEN_2552 = 8'h4 < length_1 ? _GEN_2456 : _GEN_2360; // @[executor.scala 290:56]
  wire [7:0] _GEN_2553 = 8'h4 < length_1 ? _GEN_2457 : _GEN_2361; // @[executor.scala 290:56]
  wire [7:0] _GEN_2554 = 8'h4 < length_1 ? _GEN_2458 : _GEN_2362; // @[executor.scala 290:56]
  wire [7:0] _GEN_2555 = 8'h4 < length_1 ? _GEN_2459 : _GEN_2363; // @[executor.scala 290:56]
  wire [7:0] _GEN_2556 = 8'h4 < length_1 ? _GEN_2460 : _GEN_2364; // @[executor.scala 290:56]
  wire [7:0] _GEN_2557 = 8'h4 < length_1 ? _GEN_2461 : _GEN_2365; // @[executor.scala 290:56]
  wire [7:0] _GEN_2558 = 8'h4 < length_1 ? _GEN_2462 : _GEN_2366; // @[executor.scala 290:56]
  wire [7:0] _GEN_2559 = 8'h4 < length_1 ? _GEN_2463 : _GEN_2367; // @[executor.scala 290:56]
  wire [7:0] _GEN_2560 = 8'h4 < length_1 ? _GEN_2464 : _GEN_2368; // @[executor.scala 290:56]
  wire [7:0] _GEN_2561 = 8'h4 < length_1 ? _GEN_2465 : _GEN_2369; // @[executor.scala 290:56]
  wire [7:0] _GEN_2562 = 8'h4 < length_1 ? _GEN_2466 : _GEN_2370; // @[executor.scala 290:56]
  wire [7:0] _GEN_2563 = 8'h4 < length_1 ? _GEN_2467 : _GEN_2371; // @[executor.scala 290:56]
  wire [7:0] _GEN_2564 = 8'h4 < length_1 ? _GEN_2468 : _GEN_2372; // @[executor.scala 290:56]
  wire [7:0] _GEN_2565 = 8'h4 < length_1 ? _GEN_2469 : _GEN_2373; // @[executor.scala 290:56]
  wire [7:0] _GEN_2566 = 8'h4 < length_1 ? _GEN_2470 : _GEN_2374; // @[executor.scala 290:56]
  wire [7:0] _GEN_2567 = 8'h4 < length_1 ? _GEN_2471 : _GEN_2375; // @[executor.scala 290:56]
  wire [7:0] _GEN_2568 = 8'h4 < length_1 ? _GEN_2472 : _GEN_2376; // @[executor.scala 290:56]
  wire [7:0] _GEN_2569 = 8'h4 < length_1 ? _GEN_2473 : _GEN_2377; // @[executor.scala 290:56]
  wire [7:0] _GEN_2570 = 8'h4 < length_1 ? _GEN_2474 : _GEN_2378; // @[executor.scala 290:56]
  wire [7:0] _GEN_2571 = 8'h4 < length_1 ? _GEN_2475 : _GEN_2379; // @[executor.scala 290:56]
  wire [7:0] _GEN_2572 = 8'h4 < length_1 ? _GEN_2476 : _GEN_2380; // @[executor.scala 290:56]
  wire [7:0] _GEN_2573 = 8'h4 < length_1 ? _GEN_2477 : _GEN_2381; // @[executor.scala 290:56]
  wire [7:0] _GEN_2574 = 8'h4 < length_1 ? _GEN_2478 : _GEN_2382; // @[executor.scala 290:56]
  wire [7:0] _GEN_2575 = 8'h4 < length_1 ? _GEN_2479 : _GEN_2383; // @[executor.scala 290:56]
  wire [7:0] _GEN_2576 = 8'h4 < length_1 ? _GEN_2480 : _GEN_2384; // @[executor.scala 290:56]
  wire [7:0] _GEN_2577 = 8'h4 < length_1 ? _GEN_2481 : _GEN_2385; // @[executor.scala 290:56]
  wire [7:0] _GEN_2578 = 8'h4 < length_1 ? _GEN_2482 : _GEN_2386; // @[executor.scala 290:56]
  wire [7:0] _GEN_2579 = 8'h4 < length_1 ? _GEN_2483 : _GEN_2387; // @[executor.scala 290:56]
  wire [7:0] _GEN_2580 = 8'h4 < length_1 ? _GEN_2484 : _GEN_2388; // @[executor.scala 290:56]
  wire [7:0] _GEN_2581 = 8'h4 < length_1 ? _GEN_2485 : _GEN_2389; // @[executor.scala 290:56]
  wire [7:0] _GEN_2582 = 8'h4 < length_1 ? _GEN_2486 : _GEN_2390; // @[executor.scala 290:56]
  wire [7:0] _GEN_2583 = 8'h4 < length_1 ? _GEN_2487 : _GEN_2391; // @[executor.scala 290:56]
  wire [7:0] _GEN_2584 = 8'h4 < length_1 ? _GEN_2488 : _GEN_2392; // @[executor.scala 290:56]
  wire [7:0] _GEN_2585 = 8'h4 < length_1 ? _GEN_2489 : _GEN_2393; // @[executor.scala 290:56]
  wire [7:0] _GEN_2586 = 8'h4 < length_1 ? _GEN_2490 : _GEN_2394; // @[executor.scala 290:56]
  wire [7:0] _GEN_2587 = 8'h4 < length_1 ? _GEN_2491 : _GEN_2395; // @[executor.scala 290:56]
  wire [7:0] _GEN_2588 = 8'h4 < length_1 ? _GEN_2492 : _GEN_2396; // @[executor.scala 290:56]
  wire [7:0] _GEN_2589 = 8'h4 < length_1 ? _GEN_2493 : _GEN_2397; // @[executor.scala 290:56]
  wire [7:0] _GEN_2590 = 8'h4 < length_1 ? _GEN_2494 : _GEN_2398; // @[executor.scala 290:56]
  wire [7:0] _GEN_2591 = 8'h4 < length_1 ? _GEN_2495 : _GEN_2399; // @[executor.scala 290:56]
  wire [7:0] _GEN_2592 = 8'h4 < length_1 ? _GEN_2496 : _GEN_2400; // @[executor.scala 290:56]
  wire [7:0] field_byte_13 = field_1[23:16]; // @[executor.scala 287:53]
  wire [7:0] total_offset_13 = offset_1 + 8'h5; // @[executor.scala 289:53]
  wire [7:0] _GEN_2593 = 7'h0 == total_offset_13[6:0] ? field_byte_13 : _GEN_2497; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2594 = 7'h1 == total_offset_13[6:0] ? field_byte_13 : _GEN_2498; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2595 = 7'h2 == total_offset_13[6:0] ? field_byte_13 : _GEN_2499; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2596 = 7'h3 == total_offset_13[6:0] ? field_byte_13 : _GEN_2500; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2597 = 7'h4 == total_offset_13[6:0] ? field_byte_13 : _GEN_2501; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2598 = 7'h5 == total_offset_13[6:0] ? field_byte_13 : _GEN_2502; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2599 = 7'h6 == total_offset_13[6:0] ? field_byte_13 : _GEN_2503; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2600 = 7'h7 == total_offset_13[6:0] ? field_byte_13 : _GEN_2504; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2601 = 7'h8 == total_offset_13[6:0] ? field_byte_13 : _GEN_2505; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2602 = 7'h9 == total_offset_13[6:0] ? field_byte_13 : _GEN_2506; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2603 = 7'ha == total_offset_13[6:0] ? field_byte_13 : _GEN_2507; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2604 = 7'hb == total_offset_13[6:0] ? field_byte_13 : _GEN_2508; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2605 = 7'hc == total_offset_13[6:0] ? field_byte_13 : _GEN_2509; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2606 = 7'hd == total_offset_13[6:0] ? field_byte_13 : _GEN_2510; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2607 = 7'he == total_offset_13[6:0] ? field_byte_13 : _GEN_2511; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2608 = 7'hf == total_offset_13[6:0] ? field_byte_13 : _GEN_2512; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2609 = 7'h10 == total_offset_13[6:0] ? field_byte_13 : _GEN_2513; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2610 = 7'h11 == total_offset_13[6:0] ? field_byte_13 : _GEN_2514; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2611 = 7'h12 == total_offset_13[6:0] ? field_byte_13 : _GEN_2515; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2612 = 7'h13 == total_offset_13[6:0] ? field_byte_13 : _GEN_2516; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2613 = 7'h14 == total_offset_13[6:0] ? field_byte_13 : _GEN_2517; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2614 = 7'h15 == total_offset_13[6:0] ? field_byte_13 : _GEN_2518; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2615 = 7'h16 == total_offset_13[6:0] ? field_byte_13 : _GEN_2519; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2616 = 7'h17 == total_offset_13[6:0] ? field_byte_13 : _GEN_2520; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2617 = 7'h18 == total_offset_13[6:0] ? field_byte_13 : _GEN_2521; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2618 = 7'h19 == total_offset_13[6:0] ? field_byte_13 : _GEN_2522; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2619 = 7'h1a == total_offset_13[6:0] ? field_byte_13 : _GEN_2523; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2620 = 7'h1b == total_offset_13[6:0] ? field_byte_13 : _GEN_2524; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2621 = 7'h1c == total_offset_13[6:0] ? field_byte_13 : _GEN_2525; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2622 = 7'h1d == total_offset_13[6:0] ? field_byte_13 : _GEN_2526; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2623 = 7'h1e == total_offset_13[6:0] ? field_byte_13 : _GEN_2527; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2624 = 7'h1f == total_offset_13[6:0] ? field_byte_13 : _GEN_2528; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2625 = 7'h20 == total_offset_13[6:0] ? field_byte_13 : _GEN_2529; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2626 = 7'h21 == total_offset_13[6:0] ? field_byte_13 : _GEN_2530; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2627 = 7'h22 == total_offset_13[6:0] ? field_byte_13 : _GEN_2531; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2628 = 7'h23 == total_offset_13[6:0] ? field_byte_13 : _GEN_2532; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2629 = 7'h24 == total_offset_13[6:0] ? field_byte_13 : _GEN_2533; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2630 = 7'h25 == total_offset_13[6:0] ? field_byte_13 : _GEN_2534; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2631 = 7'h26 == total_offset_13[6:0] ? field_byte_13 : _GEN_2535; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2632 = 7'h27 == total_offset_13[6:0] ? field_byte_13 : _GEN_2536; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2633 = 7'h28 == total_offset_13[6:0] ? field_byte_13 : _GEN_2537; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2634 = 7'h29 == total_offset_13[6:0] ? field_byte_13 : _GEN_2538; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2635 = 7'h2a == total_offset_13[6:0] ? field_byte_13 : _GEN_2539; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2636 = 7'h2b == total_offset_13[6:0] ? field_byte_13 : _GEN_2540; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2637 = 7'h2c == total_offset_13[6:0] ? field_byte_13 : _GEN_2541; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2638 = 7'h2d == total_offset_13[6:0] ? field_byte_13 : _GEN_2542; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2639 = 7'h2e == total_offset_13[6:0] ? field_byte_13 : _GEN_2543; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2640 = 7'h2f == total_offset_13[6:0] ? field_byte_13 : _GEN_2544; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2641 = 7'h30 == total_offset_13[6:0] ? field_byte_13 : _GEN_2545; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2642 = 7'h31 == total_offset_13[6:0] ? field_byte_13 : _GEN_2546; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2643 = 7'h32 == total_offset_13[6:0] ? field_byte_13 : _GEN_2547; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2644 = 7'h33 == total_offset_13[6:0] ? field_byte_13 : _GEN_2548; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2645 = 7'h34 == total_offset_13[6:0] ? field_byte_13 : _GEN_2549; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2646 = 7'h35 == total_offset_13[6:0] ? field_byte_13 : _GEN_2550; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2647 = 7'h36 == total_offset_13[6:0] ? field_byte_13 : _GEN_2551; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2648 = 7'h37 == total_offset_13[6:0] ? field_byte_13 : _GEN_2552; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2649 = 7'h38 == total_offset_13[6:0] ? field_byte_13 : _GEN_2553; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2650 = 7'h39 == total_offset_13[6:0] ? field_byte_13 : _GEN_2554; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2651 = 7'h3a == total_offset_13[6:0] ? field_byte_13 : _GEN_2555; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2652 = 7'h3b == total_offset_13[6:0] ? field_byte_13 : _GEN_2556; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2653 = 7'h3c == total_offset_13[6:0] ? field_byte_13 : _GEN_2557; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2654 = 7'h3d == total_offset_13[6:0] ? field_byte_13 : _GEN_2558; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2655 = 7'h3e == total_offset_13[6:0] ? field_byte_13 : _GEN_2559; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2656 = 7'h3f == total_offset_13[6:0] ? field_byte_13 : _GEN_2560; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2657 = 7'h40 == total_offset_13[6:0] ? field_byte_13 : _GEN_2561; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2658 = 7'h41 == total_offset_13[6:0] ? field_byte_13 : _GEN_2562; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2659 = 7'h42 == total_offset_13[6:0] ? field_byte_13 : _GEN_2563; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2660 = 7'h43 == total_offset_13[6:0] ? field_byte_13 : _GEN_2564; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2661 = 7'h44 == total_offset_13[6:0] ? field_byte_13 : _GEN_2565; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2662 = 7'h45 == total_offset_13[6:0] ? field_byte_13 : _GEN_2566; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2663 = 7'h46 == total_offset_13[6:0] ? field_byte_13 : _GEN_2567; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2664 = 7'h47 == total_offset_13[6:0] ? field_byte_13 : _GEN_2568; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2665 = 7'h48 == total_offset_13[6:0] ? field_byte_13 : _GEN_2569; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2666 = 7'h49 == total_offset_13[6:0] ? field_byte_13 : _GEN_2570; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2667 = 7'h4a == total_offset_13[6:0] ? field_byte_13 : _GEN_2571; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2668 = 7'h4b == total_offset_13[6:0] ? field_byte_13 : _GEN_2572; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2669 = 7'h4c == total_offset_13[6:0] ? field_byte_13 : _GEN_2573; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2670 = 7'h4d == total_offset_13[6:0] ? field_byte_13 : _GEN_2574; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2671 = 7'h4e == total_offset_13[6:0] ? field_byte_13 : _GEN_2575; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2672 = 7'h4f == total_offset_13[6:0] ? field_byte_13 : _GEN_2576; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2673 = 7'h50 == total_offset_13[6:0] ? field_byte_13 : _GEN_2577; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2674 = 7'h51 == total_offset_13[6:0] ? field_byte_13 : _GEN_2578; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2675 = 7'h52 == total_offset_13[6:0] ? field_byte_13 : _GEN_2579; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2676 = 7'h53 == total_offset_13[6:0] ? field_byte_13 : _GEN_2580; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2677 = 7'h54 == total_offset_13[6:0] ? field_byte_13 : _GEN_2581; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2678 = 7'h55 == total_offset_13[6:0] ? field_byte_13 : _GEN_2582; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2679 = 7'h56 == total_offset_13[6:0] ? field_byte_13 : _GEN_2583; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2680 = 7'h57 == total_offset_13[6:0] ? field_byte_13 : _GEN_2584; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2681 = 7'h58 == total_offset_13[6:0] ? field_byte_13 : _GEN_2585; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2682 = 7'h59 == total_offset_13[6:0] ? field_byte_13 : _GEN_2586; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2683 = 7'h5a == total_offset_13[6:0] ? field_byte_13 : _GEN_2587; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2684 = 7'h5b == total_offset_13[6:0] ? field_byte_13 : _GEN_2588; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2685 = 7'h5c == total_offset_13[6:0] ? field_byte_13 : _GEN_2589; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2686 = 7'h5d == total_offset_13[6:0] ? field_byte_13 : _GEN_2590; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2687 = 7'h5e == total_offset_13[6:0] ? field_byte_13 : _GEN_2591; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2688 = 7'h5f == total_offset_13[6:0] ? field_byte_13 : _GEN_2592; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2689 = 8'h5 < length_1 ? _GEN_2593 : _GEN_2497; // @[executor.scala 290:56]
  wire [7:0] _GEN_2690 = 8'h5 < length_1 ? _GEN_2594 : _GEN_2498; // @[executor.scala 290:56]
  wire [7:0] _GEN_2691 = 8'h5 < length_1 ? _GEN_2595 : _GEN_2499; // @[executor.scala 290:56]
  wire [7:0] _GEN_2692 = 8'h5 < length_1 ? _GEN_2596 : _GEN_2500; // @[executor.scala 290:56]
  wire [7:0] _GEN_2693 = 8'h5 < length_1 ? _GEN_2597 : _GEN_2501; // @[executor.scala 290:56]
  wire [7:0] _GEN_2694 = 8'h5 < length_1 ? _GEN_2598 : _GEN_2502; // @[executor.scala 290:56]
  wire [7:0] _GEN_2695 = 8'h5 < length_1 ? _GEN_2599 : _GEN_2503; // @[executor.scala 290:56]
  wire [7:0] _GEN_2696 = 8'h5 < length_1 ? _GEN_2600 : _GEN_2504; // @[executor.scala 290:56]
  wire [7:0] _GEN_2697 = 8'h5 < length_1 ? _GEN_2601 : _GEN_2505; // @[executor.scala 290:56]
  wire [7:0] _GEN_2698 = 8'h5 < length_1 ? _GEN_2602 : _GEN_2506; // @[executor.scala 290:56]
  wire [7:0] _GEN_2699 = 8'h5 < length_1 ? _GEN_2603 : _GEN_2507; // @[executor.scala 290:56]
  wire [7:0] _GEN_2700 = 8'h5 < length_1 ? _GEN_2604 : _GEN_2508; // @[executor.scala 290:56]
  wire [7:0] _GEN_2701 = 8'h5 < length_1 ? _GEN_2605 : _GEN_2509; // @[executor.scala 290:56]
  wire [7:0] _GEN_2702 = 8'h5 < length_1 ? _GEN_2606 : _GEN_2510; // @[executor.scala 290:56]
  wire [7:0] _GEN_2703 = 8'h5 < length_1 ? _GEN_2607 : _GEN_2511; // @[executor.scala 290:56]
  wire [7:0] _GEN_2704 = 8'h5 < length_1 ? _GEN_2608 : _GEN_2512; // @[executor.scala 290:56]
  wire [7:0] _GEN_2705 = 8'h5 < length_1 ? _GEN_2609 : _GEN_2513; // @[executor.scala 290:56]
  wire [7:0] _GEN_2706 = 8'h5 < length_1 ? _GEN_2610 : _GEN_2514; // @[executor.scala 290:56]
  wire [7:0] _GEN_2707 = 8'h5 < length_1 ? _GEN_2611 : _GEN_2515; // @[executor.scala 290:56]
  wire [7:0] _GEN_2708 = 8'h5 < length_1 ? _GEN_2612 : _GEN_2516; // @[executor.scala 290:56]
  wire [7:0] _GEN_2709 = 8'h5 < length_1 ? _GEN_2613 : _GEN_2517; // @[executor.scala 290:56]
  wire [7:0] _GEN_2710 = 8'h5 < length_1 ? _GEN_2614 : _GEN_2518; // @[executor.scala 290:56]
  wire [7:0] _GEN_2711 = 8'h5 < length_1 ? _GEN_2615 : _GEN_2519; // @[executor.scala 290:56]
  wire [7:0] _GEN_2712 = 8'h5 < length_1 ? _GEN_2616 : _GEN_2520; // @[executor.scala 290:56]
  wire [7:0] _GEN_2713 = 8'h5 < length_1 ? _GEN_2617 : _GEN_2521; // @[executor.scala 290:56]
  wire [7:0] _GEN_2714 = 8'h5 < length_1 ? _GEN_2618 : _GEN_2522; // @[executor.scala 290:56]
  wire [7:0] _GEN_2715 = 8'h5 < length_1 ? _GEN_2619 : _GEN_2523; // @[executor.scala 290:56]
  wire [7:0] _GEN_2716 = 8'h5 < length_1 ? _GEN_2620 : _GEN_2524; // @[executor.scala 290:56]
  wire [7:0] _GEN_2717 = 8'h5 < length_1 ? _GEN_2621 : _GEN_2525; // @[executor.scala 290:56]
  wire [7:0] _GEN_2718 = 8'h5 < length_1 ? _GEN_2622 : _GEN_2526; // @[executor.scala 290:56]
  wire [7:0] _GEN_2719 = 8'h5 < length_1 ? _GEN_2623 : _GEN_2527; // @[executor.scala 290:56]
  wire [7:0] _GEN_2720 = 8'h5 < length_1 ? _GEN_2624 : _GEN_2528; // @[executor.scala 290:56]
  wire [7:0] _GEN_2721 = 8'h5 < length_1 ? _GEN_2625 : _GEN_2529; // @[executor.scala 290:56]
  wire [7:0] _GEN_2722 = 8'h5 < length_1 ? _GEN_2626 : _GEN_2530; // @[executor.scala 290:56]
  wire [7:0] _GEN_2723 = 8'h5 < length_1 ? _GEN_2627 : _GEN_2531; // @[executor.scala 290:56]
  wire [7:0] _GEN_2724 = 8'h5 < length_1 ? _GEN_2628 : _GEN_2532; // @[executor.scala 290:56]
  wire [7:0] _GEN_2725 = 8'h5 < length_1 ? _GEN_2629 : _GEN_2533; // @[executor.scala 290:56]
  wire [7:0] _GEN_2726 = 8'h5 < length_1 ? _GEN_2630 : _GEN_2534; // @[executor.scala 290:56]
  wire [7:0] _GEN_2727 = 8'h5 < length_1 ? _GEN_2631 : _GEN_2535; // @[executor.scala 290:56]
  wire [7:0] _GEN_2728 = 8'h5 < length_1 ? _GEN_2632 : _GEN_2536; // @[executor.scala 290:56]
  wire [7:0] _GEN_2729 = 8'h5 < length_1 ? _GEN_2633 : _GEN_2537; // @[executor.scala 290:56]
  wire [7:0] _GEN_2730 = 8'h5 < length_1 ? _GEN_2634 : _GEN_2538; // @[executor.scala 290:56]
  wire [7:0] _GEN_2731 = 8'h5 < length_1 ? _GEN_2635 : _GEN_2539; // @[executor.scala 290:56]
  wire [7:0] _GEN_2732 = 8'h5 < length_1 ? _GEN_2636 : _GEN_2540; // @[executor.scala 290:56]
  wire [7:0] _GEN_2733 = 8'h5 < length_1 ? _GEN_2637 : _GEN_2541; // @[executor.scala 290:56]
  wire [7:0] _GEN_2734 = 8'h5 < length_1 ? _GEN_2638 : _GEN_2542; // @[executor.scala 290:56]
  wire [7:0] _GEN_2735 = 8'h5 < length_1 ? _GEN_2639 : _GEN_2543; // @[executor.scala 290:56]
  wire [7:0] _GEN_2736 = 8'h5 < length_1 ? _GEN_2640 : _GEN_2544; // @[executor.scala 290:56]
  wire [7:0] _GEN_2737 = 8'h5 < length_1 ? _GEN_2641 : _GEN_2545; // @[executor.scala 290:56]
  wire [7:0] _GEN_2738 = 8'h5 < length_1 ? _GEN_2642 : _GEN_2546; // @[executor.scala 290:56]
  wire [7:0] _GEN_2739 = 8'h5 < length_1 ? _GEN_2643 : _GEN_2547; // @[executor.scala 290:56]
  wire [7:0] _GEN_2740 = 8'h5 < length_1 ? _GEN_2644 : _GEN_2548; // @[executor.scala 290:56]
  wire [7:0] _GEN_2741 = 8'h5 < length_1 ? _GEN_2645 : _GEN_2549; // @[executor.scala 290:56]
  wire [7:0] _GEN_2742 = 8'h5 < length_1 ? _GEN_2646 : _GEN_2550; // @[executor.scala 290:56]
  wire [7:0] _GEN_2743 = 8'h5 < length_1 ? _GEN_2647 : _GEN_2551; // @[executor.scala 290:56]
  wire [7:0] _GEN_2744 = 8'h5 < length_1 ? _GEN_2648 : _GEN_2552; // @[executor.scala 290:56]
  wire [7:0] _GEN_2745 = 8'h5 < length_1 ? _GEN_2649 : _GEN_2553; // @[executor.scala 290:56]
  wire [7:0] _GEN_2746 = 8'h5 < length_1 ? _GEN_2650 : _GEN_2554; // @[executor.scala 290:56]
  wire [7:0] _GEN_2747 = 8'h5 < length_1 ? _GEN_2651 : _GEN_2555; // @[executor.scala 290:56]
  wire [7:0] _GEN_2748 = 8'h5 < length_1 ? _GEN_2652 : _GEN_2556; // @[executor.scala 290:56]
  wire [7:0] _GEN_2749 = 8'h5 < length_1 ? _GEN_2653 : _GEN_2557; // @[executor.scala 290:56]
  wire [7:0] _GEN_2750 = 8'h5 < length_1 ? _GEN_2654 : _GEN_2558; // @[executor.scala 290:56]
  wire [7:0] _GEN_2751 = 8'h5 < length_1 ? _GEN_2655 : _GEN_2559; // @[executor.scala 290:56]
  wire [7:0] _GEN_2752 = 8'h5 < length_1 ? _GEN_2656 : _GEN_2560; // @[executor.scala 290:56]
  wire [7:0] _GEN_2753 = 8'h5 < length_1 ? _GEN_2657 : _GEN_2561; // @[executor.scala 290:56]
  wire [7:0] _GEN_2754 = 8'h5 < length_1 ? _GEN_2658 : _GEN_2562; // @[executor.scala 290:56]
  wire [7:0] _GEN_2755 = 8'h5 < length_1 ? _GEN_2659 : _GEN_2563; // @[executor.scala 290:56]
  wire [7:0] _GEN_2756 = 8'h5 < length_1 ? _GEN_2660 : _GEN_2564; // @[executor.scala 290:56]
  wire [7:0] _GEN_2757 = 8'h5 < length_1 ? _GEN_2661 : _GEN_2565; // @[executor.scala 290:56]
  wire [7:0] _GEN_2758 = 8'h5 < length_1 ? _GEN_2662 : _GEN_2566; // @[executor.scala 290:56]
  wire [7:0] _GEN_2759 = 8'h5 < length_1 ? _GEN_2663 : _GEN_2567; // @[executor.scala 290:56]
  wire [7:0] _GEN_2760 = 8'h5 < length_1 ? _GEN_2664 : _GEN_2568; // @[executor.scala 290:56]
  wire [7:0] _GEN_2761 = 8'h5 < length_1 ? _GEN_2665 : _GEN_2569; // @[executor.scala 290:56]
  wire [7:0] _GEN_2762 = 8'h5 < length_1 ? _GEN_2666 : _GEN_2570; // @[executor.scala 290:56]
  wire [7:0] _GEN_2763 = 8'h5 < length_1 ? _GEN_2667 : _GEN_2571; // @[executor.scala 290:56]
  wire [7:0] _GEN_2764 = 8'h5 < length_1 ? _GEN_2668 : _GEN_2572; // @[executor.scala 290:56]
  wire [7:0] _GEN_2765 = 8'h5 < length_1 ? _GEN_2669 : _GEN_2573; // @[executor.scala 290:56]
  wire [7:0] _GEN_2766 = 8'h5 < length_1 ? _GEN_2670 : _GEN_2574; // @[executor.scala 290:56]
  wire [7:0] _GEN_2767 = 8'h5 < length_1 ? _GEN_2671 : _GEN_2575; // @[executor.scala 290:56]
  wire [7:0] _GEN_2768 = 8'h5 < length_1 ? _GEN_2672 : _GEN_2576; // @[executor.scala 290:56]
  wire [7:0] _GEN_2769 = 8'h5 < length_1 ? _GEN_2673 : _GEN_2577; // @[executor.scala 290:56]
  wire [7:0] _GEN_2770 = 8'h5 < length_1 ? _GEN_2674 : _GEN_2578; // @[executor.scala 290:56]
  wire [7:0] _GEN_2771 = 8'h5 < length_1 ? _GEN_2675 : _GEN_2579; // @[executor.scala 290:56]
  wire [7:0] _GEN_2772 = 8'h5 < length_1 ? _GEN_2676 : _GEN_2580; // @[executor.scala 290:56]
  wire [7:0] _GEN_2773 = 8'h5 < length_1 ? _GEN_2677 : _GEN_2581; // @[executor.scala 290:56]
  wire [7:0] _GEN_2774 = 8'h5 < length_1 ? _GEN_2678 : _GEN_2582; // @[executor.scala 290:56]
  wire [7:0] _GEN_2775 = 8'h5 < length_1 ? _GEN_2679 : _GEN_2583; // @[executor.scala 290:56]
  wire [7:0] _GEN_2776 = 8'h5 < length_1 ? _GEN_2680 : _GEN_2584; // @[executor.scala 290:56]
  wire [7:0] _GEN_2777 = 8'h5 < length_1 ? _GEN_2681 : _GEN_2585; // @[executor.scala 290:56]
  wire [7:0] _GEN_2778 = 8'h5 < length_1 ? _GEN_2682 : _GEN_2586; // @[executor.scala 290:56]
  wire [7:0] _GEN_2779 = 8'h5 < length_1 ? _GEN_2683 : _GEN_2587; // @[executor.scala 290:56]
  wire [7:0] _GEN_2780 = 8'h5 < length_1 ? _GEN_2684 : _GEN_2588; // @[executor.scala 290:56]
  wire [7:0] _GEN_2781 = 8'h5 < length_1 ? _GEN_2685 : _GEN_2589; // @[executor.scala 290:56]
  wire [7:0] _GEN_2782 = 8'h5 < length_1 ? _GEN_2686 : _GEN_2590; // @[executor.scala 290:56]
  wire [7:0] _GEN_2783 = 8'h5 < length_1 ? _GEN_2687 : _GEN_2591; // @[executor.scala 290:56]
  wire [7:0] _GEN_2784 = 8'h5 < length_1 ? _GEN_2688 : _GEN_2592; // @[executor.scala 290:56]
  wire [7:0] field_byte_14 = field_1[15:8]; // @[executor.scala 287:53]
  wire [7:0] total_offset_14 = offset_1 + 8'h6; // @[executor.scala 289:53]
  wire [7:0] _GEN_2785 = 7'h0 == total_offset_14[6:0] ? field_byte_14 : _GEN_2689; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2786 = 7'h1 == total_offset_14[6:0] ? field_byte_14 : _GEN_2690; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2787 = 7'h2 == total_offset_14[6:0] ? field_byte_14 : _GEN_2691; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2788 = 7'h3 == total_offset_14[6:0] ? field_byte_14 : _GEN_2692; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2789 = 7'h4 == total_offset_14[6:0] ? field_byte_14 : _GEN_2693; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2790 = 7'h5 == total_offset_14[6:0] ? field_byte_14 : _GEN_2694; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2791 = 7'h6 == total_offset_14[6:0] ? field_byte_14 : _GEN_2695; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2792 = 7'h7 == total_offset_14[6:0] ? field_byte_14 : _GEN_2696; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2793 = 7'h8 == total_offset_14[6:0] ? field_byte_14 : _GEN_2697; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2794 = 7'h9 == total_offset_14[6:0] ? field_byte_14 : _GEN_2698; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2795 = 7'ha == total_offset_14[6:0] ? field_byte_14 : _GEN_2699; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2796 = 7'hb == total_offset_14[6:0] ? field_byte_14 : _GEN_2700; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2797 = 7'hc == total_offset_14[6:0] ? field_byte_14 : _GEN_2701; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2798 = 7'hd == total_offset_14[6:0] ? field_byte_14 : _GEN_2702; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2799 = 7'he == total_offset_14[6:0] ? field_byte_14 : _GEN_2703; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2800 = 7'hf == total_offset_14[6:0] ? field_byte_14 : _GEN_2704; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2801 = 7'h10 == total_offset_14[6:0] ? field_byte_14 : _GEN_2705; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2802 = 7'h11 == total_offset_14[6:0] ? field_byte_14 : _GEN_2706; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2803 = 7'h12 == total_offset_14[6:0] ? field_byte_14 : _GEN_2707; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2804 = 7'h13 == total_offset_14[6:0] ? field_byte_14 : _GEN_2708; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2805 = 7'h14 == total_offset_14[6:0] ? field_byte_14 : _GEN_2709; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2806 = 7'h15 == total_offset_14[6:0] ? field_byte_14 : _GEN_2710; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2807 = 7'h16 == total_offset_14[6:0] ? field_byte_14 : _GEN_2711; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2808 = 7'h17 == total_offset_14[6:0] ? field_byte_14 : _GEN_2712; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2809 = 7'h18 == total_offset_14[6:0] ? field_byte_14 : _GEN_2713; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2810 = 7'h19 == total_offset_14[6:0] ? field_byte_14 : _GEN_2714; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2811 = 7'h1a == total_offset_14[6:0] ? field_byte_14 : _GEN_2715; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2812 = 7'h1b == total_offset_14[6:0] ? field_byte_14 : _GEN_2716; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2813 = 7'h1c == total_offset_14[6:0] ? field_byte_14 : _GEN_2717; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2814 = 7'h1d == total_offset_14[6:0] ? field_byte_14 : _GEN_2718; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2815 = 7'h1e == total_offset_14[6:0] ? field_byte_14 : _GEN_2719; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2816 = 7'h1f == total_offset_14[6:0] ? field_byte_14 : _GEN_2720; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2817 = 7'h20 == total_offset_14[6:0] ? field_byte_14 : _GEN_2721; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2818 = 7'h21 == total_offset_14[6:0] ? field_byte_14 : _GEN_2722; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2819 = 7'h22 == total_offset_14[6:0] ? field_byte_14 : _GEN_2723; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2820 = 7'h23 == total_offset_14[6:0] ? field_byte_14 : _GEN_2724; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2821 = 7'h24 == total_offset_14[6:0] ? field_byte_14 : _GEN_2725; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2822 = 7'h25 == total_offset_14[6:0] ? field_byte_14 : _GEN_2726; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2823 = 7'h26 == total_offset_14[6:0] ? field_byte_14 : _GEN_2727; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2824 = 7'h27 == total_offset_14[6:0] ? field_byte_14 : _GEN_2728; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2825 = 7'h28 == total_offset_14[6:0] ? field_byte_14 : _GEN_2729; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2826 = 7'h29 == total_offset_14[6:0] ? field_byte_14 : _GEN_2730; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2827 = 7'h2a == total_offset_14[6:0] ? field_byte_14 : _GEN_2731; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2828 = 7'h2b == total_offset_14[6:0] ? field_byte_14 : _GEN_2732; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2829 = 7'h2c == total_offset_14[6:0] ? field_byte_14 : _GEN_2733; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2830 = 7'h2d == total_offset_14[6:0] ? field_byte_14 : _GEN_2734; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2831 = 7'h2e == total_offset_14[6:0] ? field_byte_14 : _GEN_2735; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2832 = 7'h2f == total_offset_14[6:0] ? field_byte_14 : _GEN_2736; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2833 = 7'h30 == total_offset_14[6:0] ? field_byte_14 : _GEN_2737; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2834 = 7'h31 == total_offset_14[6:0] ? field_byte_14 : _GEN_2738; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2835 = 7'h32 == total_offset_14[6:0] ? field_byte_14 : _GEN_2739; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2836 = 7'h33 == total_offset_14[6:0] ? field_byte_14 : _GEN_2740; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2837 = 7'h34 == total_offset_14[6:0] ? field_byte_14 : _GEN_2741; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2838 = 7'h35 == total_offset_14[6:0] ? field_byte_14 : _GEN_2742; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2839 = 7'h36 == total_offset_14[6:0] ? field_byte_14 : _GEN_2743; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2840 = 7'h37 == total_offset_14[6:0] ? field_byte_14 : _GEN_2744; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2841 = 7'h38 == total_offset_14[6:0] ? field_byte_14 : _GEN_2745; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2842 = 7'h39 == total_offset_14[6:0] ? field_byte_14 : _GEN_2746; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2843 = 7'h3a == total_offset_14[6:0] ? field_byte_14 : _GEN_2747; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2844 = 7'h3b == total_offset_14[6:0] ? field_byte_14 : _GEN_2748; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2845 = 7'h3c == total_offset_14[6:0] ? field_byte_14 : _GEN_2749; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2846 = 7'h3d == total_offset_14[6:0] ? field_byte_14 : _GEN_2750; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2847 = 7'h3e == total_offset_14[6:0] ? field_byte_14 : _GEN_2751; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2848 = 7'h3f == total_offset_14[6:0] ? field_byte_14 : _GEN_2752; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2849 = 7'h40 == total_offset_14[6:0] ? field_byte_14 : _GEN_2753; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2850 = 7'h41 == total_offset_14[6:0] ? field_byte_14 : _GEN_2754; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2851 = 7'h42 == total_offset_14[6:0] ? field_byte_14 : _GEN_2755; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2852 = 7'h43 == total_offset_14[6:0] ? field_byte_14 : _GEN_2756; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2853 = 7'h44 == total_offset_14[6:0] ? field_byte_14 : _GEN_2757; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2854 = 7'h45 == total_offset_14[6:0] ? field_byte_14 : _GEN_2758; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2855 = 7'h46 == total_offset_14[6:0] ? field_byte_14 : _GEN_2759; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2856 = 7'h47 == total_offset_14[6:0] ? field_byte_14 : _GEN_2760; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2857 = 7'h48 == total_offset_14[6:0] ? field_byte_14 : _GEN_2761; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2858 = 7'h49 == total_offset_14[6:0] ? field_byte_14 : _GEN_2762; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2859 = 7'h4a == total_offset_14[6:0] ? field_byte_14 : _GEN_2763; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2860 = 7'h4b == total_offset_14[6:0] ? field_byte_14 : _GEN_2764; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2861 = 7'h4c == total_offset_14[6:0] ? field_byte_14 : _GEN_2765; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2862 = 7'h4d == total_offset_14[6:0] ? field_byte_14 : _GEN_2766; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2863 = 7'h4e == total_offset_14[6:0] ? field_byte_14 : _GEN_2767; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2864 = 7'h4f == total_offset_14[6:0] ? field_byte_14 : _GEN_2768; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2865 = 7'h50 == total_offset_14[6:0] ? field_byte_14 : _GEN_2769; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2866 = 7'h51 == total_offset_14[6:0] ? field_byte_14 : _GEN_2770; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2867 = 7'h52 == total_offset_14[6:0] ? field_byte_14 : _GEN_2771; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2868 = 7'h53 == total_offset_14[6:0] ? field_byte_14 : _GEN_2772; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2869 = 7'h54 == total_offset_14[6:0] ? field_byte_14 : _GEN_2773; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2870 = 7'h55 == total_offset_14[6:0] ? field_byte_14 : _GEN_2774; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2871 = 7'h56 == total_offset_14[6:0] ? field_byte_14 : _GEN_2775; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2872 = 7'h57 == total_offset_14[6:0] ? field_byte_14 : _GEN_2776; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2873 = 7'h58 == total_offset_14[6:0] ? field_byte_14 : _GEN_2777; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2874 = 7'h59 == total_offset_14[6:0] ? field_byte_14 : _GEN_2778; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2875 = 7'h5a == total_offset_14[6:0] ? field_byte_14 : _GEN_2779; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2876 = 7'h5b == total_offset_14[6:0] ? field_byte_14 : _GEN_2780; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2877 = 7'h5c == total_offset_14[6:0] ? field_byte_14 : _GEN_2781; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2878 = 7'h5d == total_offset_14[6:0] ? field_byte_14 : _GEN_2782; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2879 = 7'h5e == total_offset_14[6:0] ? field_byte_14 : _GEN_2783; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2880 = 7'h5f == total_offset_14[6:0] ? field_byte_14 : _GEN_2784; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2881 = 8'h6 < length_1 ? _GEN_2785 : _GEN_2689; // @[executor.scala 290:56]
  wire [7:0] _GEN_2882 = 8'h6 < length_1 ? _GEN_2786 : _GEN_2690; // @[executor.scala 290:56]
  wire [7:0] _GEN_2883 = 8'h6 < length_1 ? _GEN_2787 : _GEN_2691; // @[executor.scala 290:56]
  wire [7:0] _GEN_2884 = 8'h6 < length_1 ? _GEN_2788 : _GEN_2692; // @[executor.scala 290:56]
  wire [7:0] _GEN_2885 = 8'h6 < length_1 ? _GEN_2789 : _GEN_2693; // @[executor.scala 290:56]
  wire [7:0] _GEN_2886 = 8'h6 < length_1 ? _GEN_2790 : _GEN_2694; // @[executor.scala 290:56]
  wire [7:0] _GEN_2887 = 8'h6 < length_1 ? _GEN_2791 : _GEN_2695; // @[executor.scala 290:56]
  wire [7:0] _GEN_2888 = 8'h6 < length_1 ? _GEN_2792 : _GEN_2696; // @[executor.scala 290:56]
  wire [7:0] _GEN_2889 = 8'h6 < length_1 ? _GEN_2793 : _GEN_2697; // @[executor.scala 290:56]
  wire [7:0] _GEN_2890 = 8'h6 < length_1 ? _GEN_2794 : _GEN_2698; // @[executor.scala 290:56]
  wire [7:0] _GEN_2891 = 8'h6 < length_1 ? _GEN_2795 : _GEN_2699; // @[executor.scala 290:56]
  wire [7:0] _GEN_2892 = 8'h6 < length_1 ? _GEN_2796 : _GEN_2700; // @[executor.scala 290:56]
  wire [7:0] _GEN_2893 = 8'h6 < length_1 ? _GEN_2797 : _GEN_2701; // @[executor.scala 290:56]
  wire [7:0] _GEN_2894 = 8'h6 < length_1 ? _GEN_2798 : _GEN_2702; // @[executor.scala 290:56]
  wire [7:0] _GEN_2895 = 8'h6 < length_1 ? _GEN_2799 : _GEN_2703; // @[executor.scala 290:56]
  wire [7:0] _GEN_2896 = 8'h6 < length_1 ? _GEN_2800 : _GEN_2704; // @[executor.scala 290:56]
  wire [7:0] _GEN_2897 = 8'h6 < length_1 ? _GEN_2801 : _GEN_2705; // @[executor.scala 290:56]
  wire [7:0] _GEN_2898 = 8'h6 < length_1 ? _GEN_2802 : _GEN_2706; // @[executor.scala 290:56]
  wire [7:0] _GEN_2899 = 8'h6 < length_1 ? _GEN_2803 : _GEN_2707; // @[executor.scala 290:56]
  wire [7:0] _GEN_2900 = 8'h6 < length_1 ? _GEN_2804 : _GEN_2708; // @[executor.scala 290:56]
  wire [7:0] _GEN_2901 = 8'h6 < length_1 ? _GEN_2805 : _GEN_2709; // @[executor.scala 290:56]
  wire [7:0] _GEN_2902 = 8'h6 < length_1 ? _GEN_2806 : _GEN_2710; // @[executor.scala 290:56]
  wire [7:0] _GEN_2903 = 8'h6 < length_1 ? _GEN_2807 : _GEN_2711; // @[executor.scala 290:56]
  wire [7:0] _GEN_2904 = 8'h6 < length_1 ? _GEN_2808 : _GEN_2712; // @[executor.scala 290:56]
  wire [7:0] _GEN_2905 = 8'h6 < length_1 ? _GEN_2809 : _GEN_2713; // @[executor.scala 290:56]
  wire [7:0] _GEN_2906 = 8'h6 < length_1 ? _GEN_2810 : _GEN_2714; // @[executor.scala 290:56]
  wire [7:0] _GEN_2907 = 8'h6 < length_1 ? _GEN_2811 : _GEN_2715; // @[executor.scala 290:56]
  wire [7:0] _GEN_2908 = 8'h6 < length_1 ? _GEN_2812 : _GEN_2716; // @[executor.scala 290:56]
  wire [7:0] _GEN_2909 = 8'h6 < length_1 ? _GEN_2813 : _GEN_2717; // @[executor.scala 290:56]
  wire [7:0] _GEN_2910 = 8'h6 < length_1 ? _GEN_2814 : _GEN_2718; // @[executor.scala 290:56]
  wire [7:0] _GEN_2911 = 8'h6 < length_1 ? _GEN_2815 : _GEN_2719; // @[executor.scala 290:56]
  wire [7:0] _GEN_2912 = 8'h6 < length_1 ? _GEN_2816 : _GEN_2720; // @[executor.scala 290:56]
  wire [7:0] _GEN_2913 = 8'h6 < length_1 ? _GEN_2817 : _GEN_2721; // @[executor.scala 290:56]
  wire [7:0] _GEN_2914 = 8'h6 < length_1 ? _GEN_2818 : _GEN_2722; // @[executor.scala 290:56]
  wire [7:0] _GEN_2915 = 8'h6 < length_1 ? _GEN_2819 : _GEN_2723; // @[executor.scala 290:56]
  wire [7:0] _GEN_2916 = 8'h6 < length_1 ? _GEN_2820 : _GEN_2724; // @[executor.scala 290:56]
  wire [7:0] _GEN_2917 = 8'h6 < length_1 ? _GEN_2821 : _GEN_2725; // @[executor.scala 290:56]
  wire [7:0] _GEN_2918 = 8'h6 < length_1 ? _GEN_2822 : _GEN_2726; // @[executor.scala 290:56]
  wire [7:0] _GEN_2919 = 8'h6 < length_1 ? _GEN_2823 : _GEN_2727; // @[executor.scala 290:56]
  wire [7:0] _GEN_2920 = 8'h6 < length_1 ? _GEN_2824 : _GEN_2728; // @[executor.scala 290:56]
  wire [7:0] _GEN_2921 = 8'h6 < length_1 ? _GEN_2825 : _GEN_2729; // @[executor.scala 290:56]
  wire [7:0] _GEN_2922 = 8'h6 < length_1 ? _GEN_2826 : _GEN_2730; // @[executor.scala 290:56]
  wire [7:0] _GEN_2923 = 8'h6 < length_1 ? _GEN_2827 : _GEN_2731; // @[executor.scala 290:56]
  wire [7:0] _GEN_2924 = 8'h6 < length_1 ? _GEN_2828 : _GEN_2732; // @[executor.scala 290:56]
  wire [7:0] _GEN_2925 = 8'h6 < length_1 ? _GEN_2829 : _GEN_2733; // @[executor.scala 290:56]
  wire [7:0] _GEN_2926 = 8'h6 < length_1 ? _GEN_2830 : _GEN_2734; // @[executor.scala 290:56]
  wire [7:0] _GEN_2927 = 8'h6 < length_1 ? _GEN_2831 : _GEN_2735; // @[executor.scala 290:56]
  wire [7:0] _GEN_2928 = 8'h6 < length_1 ? _GEN_2832 : _GEN_2736; // @[executor.scala 290:56]
  wire [7:0] _GEN_2929 = 8'h6 < length_1 ? _GEN_2833 : _GEN_2737; // @[executor.scala 290:56]
  wire [7:0] _GEN_2930 = 8'h6 < length_1 ? _GEN_2834 : _GEN_2738; // @[executor.scala 290:56]
  wire [7:0] _GEN_2931 = 8'h6 < length_1 ? _GEN_2835 : _GEN_2739; // @[executor.scala 290:56]
  wire [7:0] _GEN_2932 = 8'h6 < length_1 ? _GEN_2836 : _GEN_2740; // @[executor.scala 290:56]
  wire [7:0] _GEN_2933 = 8'h6 < length_1 ? _GEN_2837 : _GEN_2741; // @[executor.scala 290:56]
  wire [7:0] _GEN_2934 = 8'h6 < length_1 ? _GEN_2838 : _GEN_2742; // @[executor.scala 290:56]
  wire [7:0] _GEN_2935 = 8'h6 < length_1 ? _GEN_2839 : _GEN_2743; // @[executor.scala 290:56]
  wire [7:0] _GEN_2936 = 8'h6 < length_1 ? _GEN_2840 : _GEN_2744; // @[executor.scala 290:56]
  wire [7:0] _GEN_2937 = 8'h6 < length_1 ? _GEN_2841 : _GEN_2745; // @[executor.scala 290:56]
  wire [7:0] _GEN_2938 = 8'h6 < length_1 ? _GEN_2842 : _GEN_2746; // @[executor.scala 290:56]
  wire [7:0] _GEN_2939 = 8'h6 < length_1 ? _GEN_2843 : _GEN_2747; // @[executor.scala 290:56]
  wire [7:0] _GEN_2940 = 8'h6 < length_1 ? _GEN_2844 : _GEN_2748; // @[executor.scala 290:56]
  wire [7:0] _GEN_2941 = 8'h6 < length_1 ? _GEN_2845 : _GEN_2749; // @[executor.scala 290:56]
  wire [7:0] _GEN_2942 = 8'h6 < length_1 ? _GEN_2846 : _GEN_2750; // @[executor.scala 290:56]
  wire [7:0] _GEN_2943 = 8'h6 < length_1 ? _GEN_2847 : _GEN_2751; // @[executor.scala 290:56]
  wire [7:0] _GEN_2944 = 8'h6 < length_1 ? _GEN_2848 : _GEN_2752; // @[executor.scala 290:56]
  wire [7:0] _GEN_2945 = 8'h6 < length_1 ? _GEN_2849 : _GEN_2753; // @[executor.scala 290:56]
  wire [7:0] _GEN_2946 = 8'h6 < length_1 ? _GEN_2850 : _GEN_2754; // @[executor.scala 290:56]
  wire [7:0] _GEN_2947 = 8'h6 < length_1 ? _GEN_2851 : _GEN_2755; // @[executor.scala 290:56]
  wire [7:0] _GEN_2948 = 8'h6 < length_1 ? _GEN_2852 : _GEN_2756; // @[executor.scala 290:56]
  wire [7:0] _GEN_2949 = 8'h6 < length_1 ? _GEN_2853 : _GEN_2757; // @[executor.scala 290:56]
  wire [7:0] _GEN_2950 = 8'h6 < length_1 ? _GEN_2854 : _GEN_2758; // @[executor.scala 290:56]
  wire [7:0] _GEN_2951 = 8'h6 < length_1 ? _GEN_2855 : _GEN_2759; // @[executor.scala 290:56]
  wire [7:0] _GEN_2952 = 8'h6 < length_1 ? _GEN_2856 : _GEN_2760; // @[executor.scala 290:56]
  wire [7:0] _GEN_2953 = 8'h6 < length_1 ? _GEN_2857 : _GEN_2761; // @[executor.scala 290:56]
  wire [7:0] _GEN_2954 = 8'h6 < length_1 ? _GEN_2858 : _GEN_2762; // @[executor.scala 290:56]
  wire [7:0] _GEN_2955 = 8'h6 < length_1 ? _GEN_2859 : _GEN_2763; // @[executor.scala 290:56]
  wire [7:0] _GEN_2956 = 8'h6 < length_1 ? _GEN_2860 : _GEN_2764; // @[executor.scala 290:56]
  wire [7:0] _GEN_2957 = 8'h6 < length_1 ? _GEN_2861 : _GEN_2765; // @[executor.scala 290:56]
  wire [7:0] _GEN_2958 = 8'h6 < length_1 ? _GEN_2862 : _GEN_2766; // @[executor.scala 290:56]
  wire [7:0] _GEN_2959 = 8'h6 < length_1 ? _GEN_2863 : _GEN_2767; // @[executor.scala 290:56]
  wire [7:0] _GEN_2960 = 8'h6 < length_1 ? _GEN_2864 : _GEN_2768; // @[executor.scala 290:56]
  wire [7:0] _GEN_2961 = 8'h6 < length_1 ? _GEN_2865 : _GEN_2769; // @[executor.scala 290:56]
  wire [7:0] _GEN_2962 = 8'h6 < length_1 ? _GEN_2866 : _GEN_2770; // @[executor.scala 290:56]
  wire [7:0] _GEN_2963 = 8'h6 < length_1 ? _GEN_2867 : _GEN_2771; // @[executor.scala 290:56]
  wire [7:0] _GEN_2964 = 8'h6 < length_1 ? _GEN_2868 : _GEN_2772; // @[executor.scala 290:56]
  wire [7:0] _GEN_2965 = 8'h6 < length_1 ? _GEN_2869 : _GEN_2773; // @[executor.scala 290:56]
  wire [7:0] _GEN_2966 = 8'h6 < length_1 ? _GEN_2870 : _GEN_2774; // @[executor.scala 290:56]
  wire [7:0] _GEN_2967 = 8'h6 < length_1 ? _GEN_2871 : _GEN_2775; // @[executor.scala 290:56]
  wire [7:0] _GEN_2968 = 8'h6 < length_1 ? _GEN_2872 : _GEN_2776; // @[executor.scala 290:56]
  wire [7:0] _GEN_2969 = 8'h6 < length_1 ? _GEN_2873 : _GEN_2777; // @[executor.scala 290:56]
  wire [7:0] _GEN_2970 = 8'h6 < length_1 ? _GEN_2874 : _GEN_2778; // @[executor.scala 290:56]
  wire [7:0] _GEN_2971 = 8'h6 < length_1 ? _GEN_2875 : _GEN_2779; // @[executor.scala 290:56]
  wire [7:0] _GEN_2972 = 8'h6 < length_1 ? _GEN_2876 : _GEN_2780; // @[executor.scala 290:56]
  wire [7:0] _GEN_2973 = 8'h6 < length_1 ? _GEN_2877 : _GEN_2781; // @[executor.scala 290:56]
  wire [7:0] _GEN_2974 = 8'h6 < length_1 ? _GEN_2878 : _GEN_2782; // @[executor.scala 290:56]
  wire [7:0] _GEN_2975 = 8'h6 < length_1 ? _GEN_2879 : _GEN_2783; // @[executor.scala 290:56]
  wire [7:0] _GEN_2976 = 8'h6 < length_1 ? _GEN_2880 : _GEN_2784; // @[executor.scala 290:56]
  wire [7:0] field_byte_15 = field_1[7:0]; // @[executor.scala 287:53]
  wire [7:0] total_offset_15 = offset_1 + 8'h7; // @[executor.scala 289:53]
  wire [7:0] _GEN_2977 = 7'h0 == total_offset_15[6:0] ? field_byte_15 : _GEN_2881; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2978 = 7'h1 == total_offset_15[6:0] ? field_byte_15 : _GEN_2882; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2979 = 7'h2 == total_offset_15[6:0] ? field_byte_15 : _GEN_2883; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2980 = 7'h3 == total_offset_15[6:0] ? field_byte_15 : _GEN_2884; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2981 = 7'h4 == total_offset_15[6:0] ? field_byte_15 : _GEN_2885; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2982 = 7'h5 == total_offset_15[6:0] ? field_byte_15 : _GEN_2886; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2983 = 7'h6 == total_offset_15[6:0] ? field_byte_15 : _GEN_2887; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2984 = 7'h7 == total_offset_15[6:0] ? field_byte_15 : _GEN_2888; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2985 = 7'h8 == total_offset_15[6:0] ? field_byte_15 : _GEN_2889; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2986 = 7'h9 == total_offset_15[6:0] ? field_byte_15 : _GEN_2890; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2987 = 7'ha == total_offset_15[6:0] ? field_byte_15 : _GEN_2891; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2988 = 7'hb == total_offset_15[6:0] ? field_byte_15 : _GEN_2892; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2989 = 7'hc == total_offset_15[6:0] ? field_byte_15 : _GEN_2893; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2990 = 7'hd == total_offset_15[6:0] ? field_byte_15 : _GEN_2894; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2991 = 7'he == total_offset_15[6:0] ? field_byte_15 : _GEN_2895; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2992 = 7'hf == total_offset_15[6:0] ? field_byte_15 : _GEN_2896; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2993 = 7'h10 == total_offset_15[6:0] ? field_byte_15 : _GEN_2897; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2994 = 7'h11 == total_offset_15[6:0] ? field_byte_15 : _GEN_2898; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2995 = 7'h12 == total_offset_15[6:0] ? field_byte_15 : _GEN_2899; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2996 = 7'h13 == total_offset_15[6:0] ? field_byte_15 : _GEN_2900; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2997 = 7'h14 == total_offset_15[6:0] ? field_byte_15 : _GEN_2901; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2998 = 7'h15 == total_offset_15[6:0] ? field_byte_15 : _GEN_2902; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_2999 = 7'h16 == total_offset_15[6:0] ? field_byte_15 : _GEN_2903; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3000 = 7'h17 == total_offset_15[6:0] ? field_byte_15 : _GEN_2904; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3001 = 7'h18 == total_offset_15[6:0] ? field_byte_15 : _GEN_2905; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3002 = 7'h19 == total_offset_15[6:0] ? field_byte_15 : _GEN_2906; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3003 = 7'h1a == total_offset_15[6:0] ? field_byte_15 : _GEN_2907; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3004 = 7'h1b == total_offset_15[6:0] ? field_byte_15 : _GEN_2908; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3005 = 7'h1c == total_offset_15[6:0] ? field_byte_15 : _GEN_2909; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3006 = 7'h1d == total_offset_15[6:0] ? field_byte_15 : _GEN_2910; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3007 = 7'h1e == total_offset_15[6:0] ? field_byte_15 : _GEN_2911; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3008 = 7'h1f == total_offset_15[6:0] ? field_byte_15 : _GEN_2912; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3009 = 7'h20 == total_offset_15[6:0] ? field_byte_15 : _GEN_2913; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3010 = 7'h21 == total_offset_15[6:0] ? field_byte_15 : _GEN_2914; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3011 = 7'h22 == total_offset_15[6:0] ? field_byte_15 : _GEN_2915; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3012 = 7'h23 == total_offset_15[6:0] ? field_byte_15 : _GEN_2916; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3013 = 7'h24 == total_offset_15[6:0] ? field_byte_15 : _GEN_2917; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3014 = 7'h25 == total_offset_15[6:0] ? field_byte_15 : _GEN_2918; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3015 = 7'h26 == total_offset_15[6:0] ? field_byte_15 : _GEN_2919; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3016 = 7'h27 == total_offset_15[6:0] ? field_byte_15 : _GEN_2920; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3017 = 7'h28 == total_offset_15[6:0] ? field_byte_15 : _GEN_2921; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3018 = 7'h29 == total_offset_15[6:0] ? field_byte_15 : _GEN_2922; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3019 = 7'h2a == total_offset_15[6:0] ? field_byte_15 : _GEN_2923; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3020 = 7'h2b == total_offset_15[6:0] ? field_byte_15 : _GEN_2924; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3021 = 7'h2c == total_offset_15[6:0] ? field_byte_15 : _GEN_2925; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3022 = 7'h2d == total_offset_15[6:0] ? field_byte_15 : _GEN_2926; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3023 = 7'h2e == total_offset_15[6:0] ? field_byte_15 : _GEN_2927; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3024 = 7'h2f == total_offset_15[6:0] ? field_byte_15 : _GEN_2928; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3025 = 7'h30 == total_offset_15[6:0] ? field_byte_15 : _GEN_2929; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3026 = 7'h31 == total_offset_15[6:0] ? field_byte_15 : _GEN_2930; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3027 = 7'h32 == total_offset_15[6:0] ? field_byte_15 : _GEN_2931; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3028 = 7'h33 == total_offset_15[6:0] ? field_byte_15 : _GEN_2932; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3029 = 7'h34 == total_offset_15[6:0] ? field_byte_15 : _GEN_2933; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3030 = 7'h35 == total_offset_15[6:0] ? field_byte_15 : _GEN_2934; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3031 = 7'h36 == total_offset_15[6:0] ? field_byte_15 : _GEN_2935; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3032 = 7'h37 == total_offset_15[6:0] ? field_byte_15 : _GEN_2936; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3033 = 7'h38 == total_offset_15[6:0] ? field_byte_15 : _GEN_2937; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3034 = 7'h39 == total_offset_15[6:0] ? field_byte_15 : _GEN_2938; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3035 = 7'h3a == total_offset_15[6:0] ? field_byte_15 : _GEN_2939; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3036 = 7'h3b == total_offset_15[6:0] ? field_byte_15 : _GEN_2940; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3037 = 7'h3c == total_offset_15[6:0] ? field_byte_15 : _GEN_2941; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3038 = 7'h3d == total_offset_15[6:0] ? field_byte_15 : _GEN_2942; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3039 = 7'h3e == total_offset_15[6:0] ? field_byte_15 : _GEN_2943; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3040 = 7'h3f == total_offset_15[6:0] ? field_byte_15 : _GEN_2944; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3041 = 7'h40 == total_offset_15[6:0] ? field_byte_15 : _GEN_2945; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3042 = 7'h41 == total_offset_15[6:0] ? field_byte_15 : _GEN_2946; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3043 = 7'h42 == total_offset_15[6:0] ? field_byte_15 : _GEN_2947; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3044 = 7'h43 == total_offset_15[6:0] ? field_byte_15 : _GEN_2948; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3045 = 7'h44 == total_offset_15[6:0] ? field_byte_15 : _GEN_2949; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3046 = 7'h45 == total_offset_15[6:0] ? field_byte_15 : _GEN_2950; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3047 = 7'h46 == total_offset_15[6:0] ? field_byte_15 : _GEN_2951; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3048 = 7'h47 == total_offset_15[6:0] ? field_byte_15 : _GEN_2952; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3049 = 7'h48 == total_offset_15[6:0] ? field_byte_15 : _GEN_2953; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3050 = 7'h49 == total_offset_15[6:0] ? field_byte_15 : _GEN_2954; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3051 = 7'h4a == total_offset_15[6:0] ? field_byte_15 : _GEN_2955; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3052 = 7'h4b == total_offset_15[6:0] ? field_byte_15 : _GEN_2956; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3053 = 7'h4c == total_offset_15[6:0] ? field_byte_15 : _GEN_2957; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3054 = 7'h4d == total_offset_15[6:0] ? field_byte_15 : _GEN_2958; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3055 = 7'h4e == total_offset_15[6:0] ? field_byte_15 : _GEN_2959; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3056 = 7'h4f == total_offset_15[6:0] ? field_byte_15 : _GEN_2960; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3057 = 7'h50 == total_offset_15[6:0] ? field_byte_15 : _GEN_2961; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3058 = 7'h51 == total_offset_15[6:0] ? field_byte_15 : _GEN_2962; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3059 = 7'h52 == total_offset_15[6:0] ? field_byte_15 : _GEN_2963; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3060 = 7'h53 == total_offset_15[6:0] ? field_byte_15 : _GEN_2964; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3061 = 7'h54 == total_offset_15[6:0] ? field_byte_15 : _GEN_2965; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3062 = 7'h55 == total_offset_15[6:0] ? field_byte_15 : _GEN_2966; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3063 = 7'h56 == total_offset_15[6:0] ? field_byte_15 : _GEN_2967; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3064 = 7'h57 == total_offset_15[6:0] ? field_byte_15 : _GEN_2968; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3065 = 7'h58 == total_offset_15[6:0] ? field_byte_15 : _GEN_2969; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3066 = 7'h59 == total_offset_15[6:0] ? field_byte_15 : _GEN_2970; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3067 = 7'h5a == total_offset_15[6:0] ? field_byte_15 : _GEN_2971; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3068 = 7'h5b == total_offset_15[6:0] ? field_byte_15 : _GEN_2972; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3069 = 7'h5c == total_offset_15[6:0] ? field_byte_15 : _GEN_2973; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3070 = 7'h5d == total_offset_15[6:0] ? field_byte_15 : _GEN_2974; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3071 = 7'h5e == total_offset_15[6:0] ? field_byte_15 : _GEN_2975; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3072 = 7'h5f == total_offset_15[6:0] ? field_byte_15 : _GEN_2976; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3073 = 8'h7 < length_1 ? _GEN_2977 : _GEN_2881; // @[executor.scala 290:56]
  wire [7:0] _GEN_3074 = 8'h7 < length_1 ? _GEN_2978 : _GEN_2882; // @[executor.scala 290:56]
  wire [7:0] _GEN_3075 = 8'h7 < length_1 ? _GEN_2979 : _GEN_2883; // @[executor.scala 290:56]
  wire [7:0] _GEN_3076 = 8'h7 < length_1 ? _GEN_2980 : _GEN_2884; // @[executor.scala 290:56]
  wire [7:0] _GEN_3077 = 8'h7 < length_1 ? _GEN_2981 : _GEN_2885; // @[executor.scala 290:56]
  wire [7:0] _GEN_3078 = 8'h7 < length_1 ? _GEN_2982 : _GEN_2886; // @[executor.scala 290:56]
  wire [7:0] _GEN_3079 = 8'h7 < length_1 ? _GEN_2983 : _GEN_2887; // @[executor.scala 290:56]
  wire [7:0] _GEN_3080 = 8'h7 < length_1 ? _GEN_2984 : _GEN_2888; // @[executor.scala 290:56]
  wire [7:0] _GEN_3081 = 8'h7 < length_1 ? _GEN_2985 : _GEN_2889; // @[executor.scala 290:56]
  wire [7:0] _GEN_3082 = 8'h7 < length_1 ? _GEN_2986 : _GEN_2890; // @[executor.scala 290:56]
  wire [7:0] _GEN_3083 = 8'h7 < length_1 ? _GEN_2987 : _GEN_2891; // @[executor.scala 290:56]
  wire [7:0] _GEN_3084 = 8'h7 < length_1 ? _GEN_2988 : _GEN_2892; // @[executor.scala 290:56]
  wire [7:0] _GEN_3085 = 8'h7 < length_1 ? _GEN_2989 : _GEN_2893; // @[executor.scala 290:56]
  wire [7:0] _GEN_3086 = 8'h7 < length_1 ? _GEN_2990 : _GEN_2894; // @[executor.scala 290:56]
  wire [7:0] _GEN_3087 = 8'h7 < length_1 ? _GEN_2991 : _GEN_2895; // @[executor.scala 290:56]
  wire [7:0] _GEN_3088 = 8'h7 < length_1 ? _GEN_2992 : _GEN_2896; // @[executor.scala 290:56]
  wire [7:0] _GEN_3089 = 8'h7 < length_1 ? _GEN_2993 : _GEN_2897; // @[executor.scala 290:56]
  wire [7:0] _GEN_3090 = 8'h7 < length_1 ? _GEN_2994 : _GEN_2898; // @[executor.scala 290:56]
  wire [7:0] _GEN_3091 = 8'h7 < length_1 ? _GEN_2995 : _GEN_2899; // @[executor.scala 290:56]
  wire [7:0] _GEN_3092 = 8'h7 < length_1 ? _GEN_2996 : _GEN_2900; // @[executor.scala 290:56]
  wire [7:0] _GEN_3093 = 8'h7 < length_1 ? _GEN_2997 : _GEN_2901; // @[executor.scala 290:56]
  wire [7:0] _GEN_3094 = 8'h7 < length_1 ? _GEN_2998 : _GEN_2902; // @[executor.scala 290:56]
  wire [7:0] _GEN_3095 = 8'h7 < length_1 ? _GEN_2999 : _GEN_2903; // @[executor.scala 290:56]
  wire [7:0] _GEN_3096 = 8'h7 < length_1 ? _GEN_3000 : _GEN_2904; // @[executor.scala 290:56]
  wire [7:0] _GEN_3097 = 8'h7 < length_1 ? _GEN_3001 : _GEN_2905; // @[executor.scala 290:56]
  wire [7:0] _GEN_3098 = 8'h7 < length_1 ? _GEN_3002 : _GEN_2906; // @[executor.scala 290:56]
  wire [7:0] _GEN_3099 = 8'h7 < length_1 ? _GEN_3003 : _GEN_2907; // @[executor.scala 290:56]
  wire [7:0] _GEN_3100 = 8'h7 < length_1 ? _GEN_3004 : _GEN_2908; // @[executor.scala 290:56]
  wire [7:0] _GEN_3101 = 8'h7 < length_1 ? _GEN_3005 : _GEN_2909; // @[executor.scala 290:56]
  wire [7:0] _GEN_3102 = 8'h7 < length_1 ? _GEN_3006 : _GEN_2910; // @[executor.scala 290:56]
  wire [7:0] _GEN_3103 = 8'h7 < length_1 ? _GEN_3007 : _GEN_2911; // @[executor.scala 290:56]
  wire [7:0] _GEN_3104 = 8'h7 < length_1 ? _GEN_3008 : _GEN_2912; // @[executor.scala 290:56]
  wire [7:0] _GEN_3105 = 8'h7 < length_1 ? _GEN_3009 : _GEN_2913; // @[executor.scala 290:56]
  wire [7:0] _GEN_3106 = 8'h7 < length_1 ? _GEN_3010 : _GEN_2914; // @[executor.scala 290:56]
  wire [7:0] _GEN_3107 = 8'h7 < length_1 ? _GEN_3011 : _GEN_2915; // @[executor.scala 290:56]
  wire [7:0] _GEN_3108 = 8'h7 < length_1 ? _GEN_3012 : _GEN_2916; // @[executor.scala 290:56]
  wire [7:0] _GEN_3109 = 8'h7 < length_1 ? _GEN_3013 : _GEN_2917; // @[executor.scala 290:56]
  wire [7:0] _GEN_3110 = 8'h7 < length_1 ? _GEN_3014 : _GEN_2918; // @[executor.scala 290:56]
  wire [7:0] _GEN_3111 = 8'h7 < length_1 ? _GEN_3015 : _GEN_2919; // @[executor.scala 290:56]
  wire [7:0] _GEN_3112 = 8'h7 < length_1 ? _GEN_3016 : _GEN_2920; // @[executor.scala 290:56]
  wire [7:0] _GEN_3113 = 8'h7 < length_1 ? _GEN_3017 : _GEN_2921; // @[executor.scala 290:56]
  wire [7:0] _GEN_3114 = 8'h7 < length_1 ? _GEN_3018 : _GEN_2922; // @[executor.scala 290:56]
  wire [7:0] _GEN_3115 = 8'h7 < length_1 ? _GEN_3019 : _GEN_2923; // @[executor.scala 290:56]
  wire [7:0] _GEN_3116 = 8'h7 < length_1 ? _GEN_3020 : _GEN_2924; // @[executor.scala 290:56]
  wire [7:0] _GEN_3117 = 8'h7 < length_1 ? _GEN_3021 : _GEN_2925; // @[executor.scala 290:56]
  wire [7:0] _GEN_3118 = 8'h7 < length_1 ? _GEN_3022 : _GEN_2926; // @[executor.scala 290:56]
  wire [7:0] _GEN_3119 = 8'h7 < length_1 ? _GEN_3023 : _GEN_2927; // @[executor.scala 290:56]
  wire [7:0] _GEN_3120 = 8'h7 < length_1 ? _GEN_3024 : _GEN_2928; // @[executor.scala 290:56]
  wire [7:0] _GEN_3121 = 8'h7 < length_1 ? _GEN_3025 : _GEN_2929; // @[executor.scala 290:56]
  wire [7:0] _GEN_3122 = 8'h7 < length_1 ? _GEN_3026 : _GEN_2930; // @[executor.scala 290:56]
  wire [7:0] _GEN_3123 = 8'h7 < length_1 ? _GEN_3027 : _GEN_2931; // @[executor.scala 290:56]
  wire [7:0] _GEN_3124 = 8'h7 < length_1 ? _GEN_3028 : _GEN_2932; // @[executor.scala 290:56]
  wire [7:0] _GEN_3125 = 8'h7 < length_1 ? _GEN_3029 : _GEN_2933; // @[executor.scala 290:56]
  wire [7:0] _GEN_3126 = 8'h7 < length_1 ? _GEN_3030 : _GEN_2934; // @[executor.scala 290:56]
  wire [7:0] _GEN_3127 = 8'h7 < length_1 ? _GEN_3031 : _GEN_2935; // @[executor.scala 290:56]
  wire [7:0] _GEN_3128 = 8'h7 < length_1 ? _GEN_3032 : _GEN_2936; // @[executor.scala 290:56]
  wire [7:0] _GEN_3129 = 8'h7 < length_1 ? _GEN_3033 : _GEN_2937; // @[executor.scala 290:56]
  wire [7:0] _GEN_3130 = 8'h7 < length_1 ? _GEN_3034 : _GEN_2938; // @[executor.scala 290:56]
  wire [7:0] _GEN_3131 = 8'h7 < length_1 ? _GEN_3035 : _GEN_2939; // @[executor.scala 290:56]
  wire [7:0] _GEN_3132 = 8'h7 < length_1 ? _GEN_3036 : _GEN_2940; // @[executor.scala 290:56]
  wire [7:0] _GEN_3133 = 8'h7 < length_1 ? _GEN_3037 : _GEN_2941; // @[executor.scala 290:56]
  wire [7:0] _GEN_3134 = 8'h7 < length_1 ? _GEN_3038 : _GEN_2942; // @[executor.scala 290:56]
  wire [7:0] _GEN_3135 = 8'h7 < length_1 ? _GEN_3039 : _GEN_2943; // @[executor.scala 290:56]
  wire [7:0] _GEN_3136 = 8'h7 < length_1 ? _GEN_3040 : _GEN_2944; // @[executor.scala 290:56]
  wire [7:0] _GEN_3137 = 8'h7 < length_1 ? _GEN_3041 : _GEN_2945; // @[executor.scala 290:56]
  wire [7:0] _GEN_3138 = 8'h7 < length_1 ? _GEN_3042 : _GEN_2946; // @[executor.scala 290:56]
  wire [7:0] _GEN_3139 = 8'h7 < length_1 ? _GEN_3043 : _GEN_2947; // @[executor.scala 290:56]
  wire [7:0] _GEN_3140 = 8'h7 < length_1 ? _GEN_3044 : _GEN_2948; // @[executor.scala 290:56]
  wire [7:0] _GEN_3141 = 8'h7 < length_1 ? _GEN_3045 : _GEN_2949; // @[executor.scala 290:56]
  wire [7:0] _GEN_3142 = 8'h7 < length_1 ? _GEN_3046 : _GEN_2950; // @[executor.scala 290:56]
  wire [7:0] _GEN_3143 = 8'h7 < length_1 ? _GEN_3047 : _GEN_2951; // @[executor.scala 290:56]
  wire [7:0] _GEN_3144 = 8'h7 < length_1 ? _GEN_3048 : _GEN_2952; // @[executor.scala 290:56]
  wire [7:0] _GEN_3145 = 8'h7 < length_1 ? _GEN_3049 : _GEN_2953; // @[executor.scala 290:56]
  wire [7:0] _GEN_3146 = 8'h7 < length_1 ? _GEN_3050 : _GEN_2954; // @[executor.scala 290:56]
  wire [7:0] _GEN_3147 = 8'h7 < length_1 ? _GEN_3051 : _GEN_2955; // @[executor.scala 290:56]
  wire [7:0] _GEN_3148 = 8'h7 < length_1 ? _GEN_3052 : _GEN_2956; // @[executor.scala 290:56]
  wire [7:0] _GEN_3149 = 8'h7 < length_1 ? _GEN_3053 : _GEN_2957; // @[executor.scala 290:56]
  wire [7:0] _GEN_3150 = 8'h7 < length_1 ? _GEN_3054 : _GEN_2958; // @[executor.scala 290:56]
  wire [7:0] _GEN_3151 = 8'h7 < length_1 ? _GEN_3055 : _GEN_2959; // @[executor.scala 290:56]
  wire [7:0] _GEN_3152 = 8'h7 < length_1 ? _GEN_3056 : _GEN_2960; // @[executor.scala 290:56]
  wire [7:0] _GEN_3153 = 8'h7 < length_1 ? _GEN_3057 : _GEN_2961; // @[executor.scala 290:56]
  wire [7:0] _GEN_3154 = 8'h7 < length_1 ? _GEN_3058 : _GEN_2962; // @[executor.scala 290:56]
  wire [7:0] _GEN_3155 = 8'h7 < length_1 ? _GEN_3059 : _GEN_2963; // @[executor.scala 290:56]
  wire [7:0] _GEN_3156 = 8'h7 < length_1 ? _GEN_3060 : _GEN_2964; // @[executor.scala 290:56]
  wire [7:0] _GEN_3157 = 8'h7 < length_1 ? _GEN_3061 : _GEN_2965; // @[executor.scala 290:56]
  wire [7:0] _GEN_3158 = 8'h7 < length_1 ? _GEN_3062 : _GEN_2966; // @[executor.scala 290:56]
  wire [7:0] _GEN_3159 = 8'h7 < length_1 ? _GEN_3063 : _GEN_2967; // @[executor.scala 290:56]
  wire [7:0] _GEN_3160 = 8'h7 < length_1 ? _GEN_3064 : _GEN_2968; // @[executor.scala 290:56]
  wire [7:0] _GEN_3161 = 8'h7 < length_1 ? _GEN_3065 : _GEN_2969; // @[executor.scala 290:56]
  wire [7:0] _GEN_3162 = 8'h7 < length_1 ? _GEN_3066 : _GEN_2970; // @[executor.scala 290:56]
  wire [7:0] _GEN_3163 = 8'h7 < length_1 ? _GEN_3067 : _GEN_2971; // @[executor.scala 290:56]
  wire [7:0] _GEN_3164 = 8'h7 < length_1 ? _GEN_3068 : _GEN_2972; // @[executor.scala 290:56]
  wire [7:0] _GEN_3165 = 8'h7 < length_1 ? _GEN_3069 : _GEN_2973; // @[executor.scala 290:56]
  wire [7:0] _GEN_3166 = 8'h7 < length_1 ? _GEN_3070 : _GEN_2974; // @[executor.scala 290:56]
  wire [7:0] _GEN_3167 = 8'h7 < length_1 ? _GEN_3071 : _GEN_2975; // @[executor.scala 290:56]
  wire [7:0] _GEN_3168 = 8'h7 < length_1 ? _GEN_3072 : _GEN_2976; // @[executor.scala 290:56]
  wire [63:0] _GEN_3169 = length_1 == 8'h0 ? field_1 : _GEN_1536; // @[executor.scala 283:67 executor.scala 284:51]
  wire [7:0] _GEN_3170 = length_1 == 8'h0 ? _GEN_1537 : _GEN_3073; // @[executor.scala 283:67]
  wire [7:0] _GEN_3171 = length_1 == 8'h0 ? _GEN_1538 : _GEN_3074; // @[executor.scala 283:67]
  wire [7:0] _GEN_3172 = length_1 == 8'h0 ? _GEN_1539 : _GEN_3075; // @[executor.scala 283:67]
  wire [7:0] _GEN_3173 = length_1 == 8'h0 ? _GEN_1540 : _GEN_3076; // @[executor.scala 283:67]
  wire [7:0] _GEN_3174 = length_1 == 8'h0 ? _GEN_1541 : _GEN_3077; // @[executor.scala 283:67]
  wire [7:0] _GEN_3175 = length_1 == 8'h0 ? _GEN_1542 : _GEN_3078; // @[executor.scala 283:67]
  wire [7:0] _GEN_3176 = length_1 == 8'h0 ? _GEN_1543 : _GEN_3079; // @[executor.scala 283:67]
  wire [7:0] _GEN_3177 = length_1 == 8'h0 ? _GEN_1544 : _GEN_3080; // @[executor.scala 283:67]
  wire [7:0] _GEN_3178 = length_1 == 8'h0 ? _GEN_1545 : _GEN_3081; // @[executor.scala 283:67]
  wire [7:0] _GEN_3179 = length_1 == 8'h0 ? _GEN_1546 : _GEN_3082; // @[executor.scala 283:67]
  wire [7:0] _GEN_3180 = length_1 == 8'h0 ? _GEN_1547 : _GEN_3083; // @[executor.scala 283:67]
  wire [7:0] _GEN_3181 = length_1 == 8'h0 ? _GEN_1548 : _GEN_3084; // @[executor.scala 283:67]
  wire [7:0] _GEN_3182 = length_1 == 8'h0 ? _GEN_1549 : _GEN_3085; // @[executor.scala 283:67]
  wire [7:0] _GEN_3183 = length_1 == 8'h0 ? _GEN_1550 : _GEN_3086; // @[executor.scala 283:67]
  wire [7:0] _GEN_3184 = length_1 == 8'h0 ? _GEN_1551 : _GEN_3087; // @[executor.scala 283:67]
  wire [7:0] _GEN_3185 = length_1 == 8'h0 ? _GEN_1552 : _GEN_3088; // @[executor.scala 283:67]
  wire [7:0] _GEN_3186 = length_1 == 8'h0 ? _GEN_1553 : _GEN_3089; // @[executor.scala 283:67]
  wire [7:0] _GEN_3187 = length_1 == 8'h0 ? _GEN_1554 : _GEN_3090; // @[executor.scala 283:67]
  wire [7:0] _GEN_3188 = length_1 == 8'h0 ? _GEN_1555 : _GEN_3091; // @[executor.scala 283:67]
  wire [7:0] _GEN_3189 = length_1 == 8'h0 ? _GEN_1556 : _GEN_3092; // @[executor.scala 283:67]
  wire [7:0] _GEN_3190 = length_1 == 8'h0 ? _GEN_1557 : _GEN_3093; // @[executor.scala 283:67]
  wire [7:0] _GEN_3191 = length_1 == 8'h0 ? _GEN_1558 : _GEN_3094; // @[executor.scala 283:67]
  wire [7:0] _GEN_3192 = length_1 == 8'h0 ? _GEN_1559 : _GEN_3095; // @[executor.scala 283:67]
  wire [7:0] _GEN_3193 = length_1 == 8'h0 ? _GEN_1560 : _GEN_3096; // @[executor.scala 283:67]
  wire [7:0] _GEN_3194 = length_1 == 8'h0 ? _GEN_1561 : _GEN_3097; // @[executor.scala 283:67]
  wire [7:0] _GEN_3195 = length_1 == 8'h0 ? _GEN_1562 : _GEN_3098; // @[executor.scala 283:67]
  wire [7:0] _GEN_3196 = length_1 == 8'h0 ? _GEN_1563 : _GEN_3099; // @[executor.scala 283:67]
  wire [7:0] _GEN_3197 = length_1 == 8'h0 ? _GEN_1564 : _GEN_3100; // @[executor.scala 283:67]
  wire [7:0] _GEN_3198 = length_1 == 8'h0 ? _GEN_1565 : _GEN_3101; // @[executor.scala 283:67]
  wire [7:0] _GEN_3199 = length_1 == 8'h0 ? _GEN_1566 : _GEN_3102; // @[executor.scala 283:67]
  wire [7:0] _GEN_3200 = length_1 == 8'h0 ? _GEN_1567 : _GEN_3103; // @[executor.scala 283:67]
  wire [7:0] _GEN_3201 = length_1 == 8'h0 ? _GEN_1568 : _GEN_3104; // @[executor.scala 283:67]
  wire [7:0] _GEN_3202 = length_1 == 8'h0 ? _GEN_1569 : _GEN_3105; // @[executor.scala 283:67]
  wire [7:0] _GEN_3203 = length_1 == 8'h0 ? _GEN_1570 : _GEN_3106; // @[executor.scala 283:67]
  wire [7:0] _GEN_3204 = length_1 == 8'h0 ? _GEN_1571 : _GEN_3107; // @[executor.scala 283:67]
  wire [7:0] _GEN_3205 = length_1 == 8'h0 ? _GEN_1572 : _GEN_3108; // @[executor.scala 283:67]
  wire [7:0] _GEN_3206 = length_1 == 8'h0 ? _GEN_1573 : _GEN_3109; // @[executor.scala 283:67]
  wire [7:0] _GEN_3207 = length_1 == 8'h0 ? _GEN_1574 : _GEN_3110; // @[executor.scala 283:67]
  wire [7:0] _GEN_3208 = length_1 == 8'h0 ? _GEN_1575 : _GEN_3111; // @[executor.scala 283:67]
  wire [7:0] _GEN_3209 = length_1 == 8'h0 ? _GEN_1576 : _GEN_3112; // @[executor.scala 283:67]
  wire [7:0] _GEN_3210 = length_1 == 8'h0 ? _GEN_1577 : _GEN_3113; // @[executor.scala 283:67]
  wire [7:0] _GEN_3211 = length_1 == 8'h0 ? _GEN_1578 : _GEN_3114; // @[executor.scala 283:67]
  wire [7:0] _GEN_3212 = length_1 == 8'h0 ? _GEN_1579 : _GEN_3115; // @[executor.scala 283:67]
  wire [7:0] _GEN_3213 = length_1 == 8'h0 ? _GEN_1580 : _GEN_3116; // @[executor.scala 283:67]
  wire [7:0] _GEN_3214 = length_1 == 8'h0 ? _GEN_1581 : _GEN_3117; // @[executor.scala 283:67]
  wire [7:0] _GEN_3215 = length_1 == 8'h0 ? _GEN_1582 : _GEN_3118; // @[executor.scala 283:67]
  wire [7:0] _GEN_3216 = length_1 == 8'h0 ? _GEN_1583 : _GEN_3119; // @[executor.scala 283:67]
  wire [7:0] _GEN_3217 = length_1 == 8'h0 ? _GEN_1584 : _GEN_3120; // @[executor.scala 283:67]
  wire [7:0] _GEN_3218 = length_1 == 8'h0 ? _GEN_1585 : _GEN_3121; // @[executor.scala 283:67]
  wire [7:0] _GEN_3219 = length_1 == 8'h0 ? _GEN_1586 : _GEN_3122; // @[executor.scala 283:67]
  wire [7:0] _GEN_3220 = length_1 == 8'h0 ? _GEN_1587 : _GEN_3123; // @[executor.scala 283:67]
  wire [7:0] _GEN_3221 = length_1 == 8'h0 ? _GEN_1588 : _GEN_3124; // @[executor.scala 283:67]
  wire [7:0] _GEN_3222 = length_1 == 8'h0 ? _GEN_1589 : _GEN_3125; // @[executor.scala 283:67]
  wire [7:0] _GEN_3223 = length_1 == 8'h0 ? _GEN_1590 : _GEN_3126; // @[executor.scala 283:67]
  wire [7:0] _GEN_3224 = length_1 == 8'h0 ? _GEN_1591 : _GEN_3127; // @[executor.scala 283:67]
  wire [7:0] _GEN_3225 = length_1 == 8'h0 ? _GEN_1592 : _GEN_3128; // @[executor.scala 283:67]
  wire [7:0] _GEN_3226 = length_1 == 8'h0 ? _GEN_1593 : _GEN_3129; // @[executor.scala 283:67]
  wire [7:0] _GEN_3227 = length_1 == 8'h0 ? _GEN_1594 : _GEN_3130; // @[executor.scala 283:67]
  wire [7:0] _GEN_3228 = length_1 == 8'h0 ? _GEN_1595 : _GEN_3131; // @[executor.scala 283:67]
  wire [7:0] _GEN_3229 = length_1 == 8'h0 ? _GEN_1596 : _GEN_3132; // @[executor.scala 283:67]
  wire [7:0] _GEN_3230 = length_1 == 8'h0 ? _GEN_1597 : _GEN_3133; // @[executor.scala 283:67]
  wire [7:0] _GEN_3231 = length_1 == 8'h0 ? _GEN_1598 : _GEN_3134; // @[executor.scala 283:67]
  wire [7:0] _GEN_3232 = length_1 == 8'h0 ? _GEN_1599 : _GEN_3135; // @[executor.scala 283:67]
  wire [7:0] _GEN_3233 = length_1 == 8'h0 ? _GEN_1600 : _GEN_3136; // @[executor.scala 283:67]
  wire [7:0] _GEN_3234 = length_1 == 8'h0 ? _GEN_1601 : _GEN_3137; // @[executor.scala 283:67]
  wire [7:0] _GEN_3235 = length_1 == 8'h0 ? _GEN_1602 : _GEN_3138; // @[executor.scala 283:67]
  wire [7:0] _GEN_3236 = length_1 == 8'h0 ? _GEN_1603 : _GEN_3139; // @[executor.scala 283:67]
  wire [7:0] _GEN_3237 = length_1 == 8'h0 ? _GEN_1604 : _GEN_3140; // @[executor.scala 283:67]
  wire [7:0] _GEN_3238 = length_1 == 8'h0 ? _GEN_1605 : _GEN_3141; // @[executor.scala 283:67]
  wire [7:0] _GEN_3239 = length_1 == 8'h0 ? _GEN_1606 : _GEN_3142; // @[executor.scala 283:67]
  wire [7:0] _GEN_3240 = length_1 == 8'h0 ? _GEN_1607 : _GEN_3143; // @[executor.scala 283:67]
  wire [7:0] _GEN_3241 = length_1 == 8'h0 ? _GEN_1608 : _GEN_3144; // @[executor.scala 283:67]
  wire [7:0] _GEN_3242 = length_1 == 8'h0 ? _GEN_1609 : _GEN_3145; // @[executor.scala 283:67]
  wire [7:0] _GEN_3243 = length_1 == 8'h0 ? _GEN_1610 : _GEN_3146; // @[executor.scala 283:67]
  wire [7:0] _GEN_3244 = length_1 == 8'h0 ? _GEN_1611 : _GEN_3147; // @[executor.scala 283:67]
  wire [7:0] _GEN_3245 = length_1 == 8'h0 ? _GEN_1612 : _GEN_3148; // @[executor.scala 283:67]
  wire [7:0] _GEN_3246 = length_1 == 8'h0 ? _GEN_1613 : _GEN_3149; // @[executor.scala 283:67]
  wire [7:0] _GEN_3247 = length_1 == 8'h0 ? _GEN_1614 : _GEN_3150; // @[executor.scala 283:67]
  wire [7:0] _GEN_3248 = length_1 == 8'h0 ? _GEN_1615 : _GEN_3151; // @[executor.scala 283:67]
  wire [7:0] _GEN_3249 = length_1 == 8'h0 ? _GEN_1616 : _GEN_3152; // @[executor.scala 283:67]
  wire [7:0] _GEN_3250 = length_1 == 8'h0 ? _GEN_1617 : _GEN_3153; // @[executor.scala 283:67]
  wire [7:0] _GEN_3251 = length_1 == 8'h0 ? _GEN_1618 : _GEN_3154; // @[executor.scala 283:67]
  wire [7:0] _GEN_3252 = length_1 == 8'h0 ? _GEN_1619 : _GEN_3155; // @[executor.scala 283:67]
  wire [7:0] _GEN_3253 = length_1 == 8'h0 ? _GEN_1620 : _GEN_3156; // @[executor.scala 283:67]
  wire [7:0] _GEN_3254 = length_1 == 8'h0 ? _GEN_1621 : _GEN_3157; // @[executor.scala 283:67]
  wire [7:0] _GEN_3255 = length_1 == 8'h0 ? _GEN_1622 : _GEN_3158; // @[executor.scala 283:67]
  wire [7:0] _GEN_3256 = length_1 == 8'h0 ? _GEN_1623 : _GEN_3159; // @[executor.scala 283:67]
  wire [7:0] _GEN_3257 = length_1 == 8'h0 ? _GEN_1624 : _GEN_3160; // @[executor.scala 283:67]
  wire [7:0] _GEN_3258 = length_1 == 8'h0 ? _GEN_1625 : _GEN_3161; // @[executor.scala 283:67]
  wire [7:0] _GEN_3259 = length_1 == 8'h0 ? _GEN_1626 : _GEN_3162; // @[executor.scala 283:67]
  wire [7:0] _GEN_3260 = length_1 == 8'h0 ? _GEN_1627 : _GEN_3163; // @[executor.scala 283:67]
  wire [7:0] _GEN_3261 = length_1 == 8'h0 ? _GEN_1628 : _GEN_3164; // @[executor.scala 283:67]
  wire [7:0] _GEN_3262 = length_1 == 8'h0 ? _GEN_1629 : _GEN_3165; // @[executor.scala 283:67]
  wire [7:0] _GEN_3263 = length_1 == 8'h0 ? _GEN_1630 : _GEN_3166; // @[executor.scala 283:67]
  wire [7:0] _GEN_3264 = length_1 == 8'h0 ? _GEN_1631 : _GEN_3167; // @[executor.scala 283:67]
  wire [7:0] _GEN_3265 = length_1 == 8'h0 ? _GEN_1632 : _GEN_3168; // @[executor.scala 283:67]
  wire [7:0] field_byte_16 = field_2[63:56]; // @[executor.scala 287:53]
  wire [8:0] _total_offset_T_16 = {{1'd0}, offset_2}; // @[executor.scala 289:53]
  wire [7:0] total_offset_16 = _total_offset_T_16[7:0]; // @[executor.scala 289:53]
  wire [7:0] _GEN_3266 = 7'h0 == total_offset_16[6:0] ? field_byte_16 : _GEN_3170; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3267 = 7'h1 == total_offset_16[6:0] ? field_byte_16 : _GEN_3171; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3268 = 7'h2 == total_offset_16[6:0] ? field_byte_16 : _GEN_3172; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3269 = 7'h3 == total_offset_16[6:0] ? field_byte_16 : _GEN_3173; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3270 = 7'h4 == total_offset_16[6:0] ? field_byte_16 : _GEN_3174; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3271 = 7'h5 == total_offset_16[6:0] ? field_byte_16 : _GEN_3175; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3272 = 7'h6 == total_offset_16[6:0] ? field_byte_16 : _GEN_3176; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3273 = 7'h7 == total_offset_16[6:0] ? field_byte_16 : _GEN_3177; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3274 = 7'h8 == total_offset_16[6:0] ? field_byte_16 : _GEN_3178; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3275 = 7'h9 == total_offset_16[6:0] ? field_byte_16 : _GEN_3179; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3276 = 7'ha == total_offset_16[6:0] ? field_byte_16 : _GEN_3180; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3277 = 7'hb == total_offset_16[6:0] ? field_byte_16 : _GEN_3181; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3278 = 7'hc == total_offset_16[6:0] ? field_byte_16 : _GEN_3182; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3279 = 7'hd == total_offset_16[6:0] ? field_byte_16 : _GEN_3183; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3280 = 7'he == total_offset_16[6:0] ? field_byte_16 : _GEN_3184; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3281 = 7'hf == total_offset_16[6:0] ? field_byte_16 : _GEN_3185; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3282 = 7'h10 == total_offset_16[6:0] ? field_byte_16 : _GEN_3186; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3283 = 7'h11 == total_offset_16[6:0] ? field_byte_16 : _GEN_3187; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3284 = 7'h12 == total_offset_16[6:0] ? field_byte_16 : _GEN_3188; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3285 = 7'h13 == total_offset_16[6:0] ? field_byte_16 : _GEN_3189; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3286 = 7'h14 == total_offset_16[6:0] ? field_byte_16 : _GEN_3190; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3287 = 7'h15 == total_offset_16[6:0] ? field_byte_16 : _GEN_3191; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3288 = 7'h16 == total_offset_16[6:0] ? field_byte_16 : _GEN_3192; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3289 = 7'h17 == total_offset_16[6:0] ? field_byte_16 : _GEN_3193; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3290 = 7'h18 == total_offset_16[6:0] ? field_byte_16 : _GEN_3194; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3291 = 7'h19 == total_offset_16[6:0] ? field_byte_16 : _GEN_3195; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3292 = 7'h1a == total_offset_16[6:0] ? field_byte_16 : _GEN_3196; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3293 = 7'h1b == total_offset_16[6:0] ? field_byte_16 : _GEN_3197; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3294 = 7'h1c == total_offset_16[6:0] ? field_byte_16 : _GEN_3198; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3295 = 7'h1d == total_offset_16[6:0] ? field_byte_16 : _GEN_3199; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3296 = 7'h1e == total_offset_16[6:0] ? field_byte_16 : _GEN_3200; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3297 = 7'h1f == total_offset_16[6:0] ? field_byte_16 : _GEN_3201; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3298 = 7'h20 == total_offset_16[6:0] ? field_byte_16 : _GEN_3202; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3299 = 7'h21 == total_offset_16[6:0] ? field_byte_16 : _GEN_3203; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3300 = 7'h22 == total_offset_16[6:0] ? field_byte_16 : _GEN_3204; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3301 = 7'h23 == total_offset_16[6:0] ? field_byte_16 : _GEN_3205; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3302 = 7'h24 == total_offset_16[6:0] ? field_byte_16 : _GEN_3206; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3303 = 7'h25 == total_offset_16[6:0] ? field_byte_16 : _GEN_3207; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3304 = 7'h26 == total_offset_16[6:0] ? field_byte_16 : _GEN_3208; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3305 = 7'h27 == total_offset_16[6:0] ? field_byte_16 : _GEN_3209; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3306 = 7'h28 == total_offset_16[6:0] ? field_byte_16 : _GEN_3210; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3307 = 7'h29 == total_offset_16[6:0] ? field_byte_16 : _GEN_3211; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3308 = 7'h2a == total_offset_16[6:0] ? field_byte_16 : _GEN_3212; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3309 = 7'h2b == total_offset_16[6:0] ? field_byte_16 : _GEN_3213; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3310 = 7'h2c == total_offset_16[6:0] ? field_byte_16 : _GEN_3214; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3311 = 7'h2d == total_offset_16[6:0] ? field_byte_16 : _GEN_3215; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3312 = 7'h2e == total_offset_16[6:0] ? field_byte_16 : _GEN_3216; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3313 = 7'h2f == total_offset_16[6:0] ? field_byte_16 : _GEN_3217; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3314 = 7'h30 == total_offset_16[6:0] ? field_byte_16 : _GEN_3218; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3315 = 7'h31 == total_offset_16[6:0] ? field_byte_16 : _GEN_3219; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3316 = 7'h32 == total_offset_16[6:0] ? field_byte_16 : _GEN_3220; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3317 = 7'h33 == total_offset_16[6:0] ? field_byte_16 : _GEN_3221; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3318 = 7'h34 == total_offset_16[6:0] ? field_byte_16 : _GEN_3222; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3319 = 7'h35 == total_offset_16[6:0] ? field_byte_16 : _GEN_3223; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3320 = 7'h36 == total_offset_16[6:0] ? field_byte_16 : _GEN_3224; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3321 = 7'h37 == total_offset_16[6:0] ? field_byte_16 : _GEN_3225; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3322 = 7'h38 == total_offset_16[6:0] ? field_byte_16 : _GEN_3226; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3323 = 7'h39 == total_offset_16[6:0] ? field_byte_16 : _GEN_3227; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3324 = 7'h3a == total_offset_16[6:0] ? field_byte_16 : _GEN_3228; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3325 = 7'h3b == total_offset_16[6:0] ? field_byte_16 : _GEN_3229; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3326 = 7'h3c == total_offset_16[6:0] ? field_byte_16 : _GEN_3230; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3327 = 7'h3d == total_offset_16[6:0] ? field_byte_16 : _GEN_3231; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3328 = 7'h3e == total_offset_16[6:0] ? field_byte_16 : _GEN_3232; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3329 = 7'h3f == total_offset_16[6:0] ? field_byte_16 : _GEN_3233; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3330 = 7'h40 == total_offset_16[6:0] ? field_byte_16 : _GEN_3234; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3331 = 7'h41 == total_offset_16[6:0] ? field_byte_16 : _GEN_3235; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3332 = 7'h42 == total_offset_16[6:0] ? field_byte_16 : _GEN_3236; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3333 = 7'h43 == total_offset_16[6:0] ? field_byte_16 : _GEN_3237; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3334 = 7'h44 == total_offset_16[6:0] ? field_byte_16 : _GEN_3238; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3335 = 7'h45 == total_offset_16[6:0] ? field_byte_16 : _GEN_3239; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3336 = 7'h46 == total_offset_16[6:0] ? field_byte_16 : _GEN_3240; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3337 = 7'h47 == total_offset_16[6:0] ? field_byte_16 : _GEN_3241; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3338 = 7'h48 == total_offset_16[6:0] ? field_byte_16 : _GEN_3242; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3339 = 7'h49 == total_offset_16[6:0] ? field_byte_16 : _GEN_3243; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3340 = 7'h4a == total_offset_16[6:0] ? field_byte_16 : _GEN_3244; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3341 = 7'h4b == total_offset_16[6:0] ? field_byte_16 : _GEN_3245; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3342 = 7'h4c == total_offset_16[6:0] ? field_byte_16 : _GEN_3246; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3343 = 7'h4d == total_offset_16[6:0] ? field_byte_16 : _GEN_3247; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3344 = 7'h4e == total_offset_16[6:0] ? field_byte_16 : _GEN_3248; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3345 = 7'h4f == total_offset_16[6:0] ? field_byte_16 : _GEN_3249; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3346 = 7'h50 == total_offset_16[6:0] ? field_byte_16 : _GEN_3250; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3347 = 7'h51 == total_offset_16[6:0] ? field_byte_16 : _GEN_3251; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3348 = 7'h52 == total_offset_16[6:0] ? field_byte_16 : _GEN_3252; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3349 = 7'h53 == total_offset_16[6:0] ? field_byte_16 : _GEN_3253; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3350 = 7'h54 == total_offset_16[6:0] ? field_byte_16 : _GEN_3254; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3351 = 7'h55 == total_offset_16[6:0] ? field_byte_16 : _GEN_3255; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3352 = 7'h56 == total_offset_16[6:0] ? field_byte_16 : _GEN_3256; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3353 = 7'h57 == total_offset_16[6:0] ? field_byte_16 : _GEN_3257; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3354 = 7'h58 == total_offset_16[6:0] ? field_byte_16 : _GEN_3258; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3355 = 7'h59 == total_offset_16[6:0] ? field_byte_16 : _GEN_3259; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3356 = 7'h5a == total_offset_16[6:0] ? field_byte_16 : _GEN_3260; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3357 = 7'h5b == total_offset_16[6:0] ? field_byte_16 : _GEN_3261; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3358 = 7'h5c == total_offset_16[6:0] ? field_byte_16 : _GEN_3262; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3359 = 7'h5d == total_offset_16[6:0] ? field_byte_16 : _GEN_3263; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3360 = 7'h5e == total_offset_16[6:0] ? field_byte_16 : _GEN_3264; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3361 = 7'h5f == total_offset_16[6:0] ? field_byte_16 : _GEN_3265; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3362 = 8'h0 < length_2 ? _GEN_3266 : _GEN_3170; // @[executor.scala 290:56]
  wire [7:0] _GEN_3363 = 8'h0 < length_2 ? _GEN_3267 : _GEN_3171; // @[executor.scala 290:56]
  wire [7:0] _GEN_3364 = 8'h0 < length_2 ? _GEN_3268 : _GEN_3172; // @[executor.scala 290:56]
  wire [7:0] _GEN_3365 = 8'h0 < length_2 ? _GEN_3269 : _GEN_3173; // @[executor.scala 290:56]
  wire [7:0] _GEN_3366 = 8'h0 < length_2 ? _GEN_3270 : _GEN_3174; // @[executor.scala 290:56]
  wire [7:0] _GEN_3367 = 8'h0 < length_2 ? _GEN_3271 : _GEN_3175; // @[executor.scala 290:56]
  wire [7:0] _GEN_3368 = 8'h0 < length_2 ? _GEN_3272 : _GEN_3176; // @[executor.scala 290:56]
  wire [7:0] _GEN_3369 = 8'h0 < length_2 ? _GEN_3273 : _GEN_3177; // @[executor.scala 290:56]
  wire [7:0] _GEN_3370 = 8'h0 < length_2 ? _GEN_3274 : _GEN_3178; // @[executor.scala 290:56]
  wire [7:0] _GEN_3371 = 8'h0 < length_2 ? _GEN_3275 : _GEN_3179; // @[executor.scala 290:56]
  wire [7:0] _GEN_3372 = 8'h0 < length_2 ? _GEN_3276 : _GEN_3180; // @[executor.scala 290:56]
  wire [7:0] _GEN_3373 = 8'h0 < length_2 ? _GEN_3277 : _GEN_3181; // @[executor.scala 290:56]
  wire [7:0] _GEN_3374 = 8'h0 < length_2 ? _GEN_3278 : _GEN_3182; // @[executor.scala 290:56]
  wire [7:0] _GEN_3375 = 8'h0 < length_2 ? _GEN_3279 : _GEN_3183; // @[executor.scala 290:56]
  wire [7:0] _GEN_3376 = 8'h0 < length_2 ? _GEN_3280 : _GEN_3184; // @[executor.scala 290:56]
  wire [7:0] _GEN_3377 = 8'h0 < length_2 ? _GEN_3281 : _GEN_3185; // @[executor.scala 290:56]
  wire [7:0] _GEN_3378 = 8'h0 < length_2 ? _GEN_3282 : _GEN_3186; // @[executor.scala 290:56]
  wire [7:0] _GEN_3379 = 8'h0 < length_2 ? _GEN_3283 : _GEN_3187; // @[executor.scala 290:56]
  wire [7:0] _GEN_3380 = 8'h0 < length_2 ? _GEN_3284 : _GEN_3188; // @[executor.scala 290:56]
  wire [7:0] _GEN_3381 = 8'h0 < length_2 ? _GEN_3285 : _GEN_3189; // @[executor.scala 290:56]
  wire [7:0] _GEN_3382 = 8'h0 < length_2 ? _GEN_3286 : _GEN_3190; // @[executor.scala 290:56]
  wire [7:0] _GEN_3383 = 8'h0 < length_2 ? _GEN_3287 : _GEN_3191; // @[executor.scala 290:56]
  wire [7:0] _GEN_3384 = 8'h0 < length_2 ? _GEN_3288 : _GEN_3192; // @[executor.scala 290:56]
  wire [7:0] _GEN_3385 = 8'h0 < length_2 ? _GEN_3289 : _GEN_3193; // @[executor.scala 290:56]
  wire [7:0] _GEN_3386 = 8'h0 < length_2 ? _GEN_3290 : _GEN_3194; // @[executor.scala 290:56]
  wire [7:0] _GEN_3387 = 8'h0 < length_2 ? _GEN_3291 : _GEN_3195; // @[executor.scala 290:56]
  wire [7:0] _GEN_3388 = 8'h0 < length_2 ? _GEN_3292 : _GEN_3196; // @[executor.scala 290:56]
  wire [7:0] _GEN_3389 = 8'h0 < length_2 ? _GEN_3293 : _GEN_3197; // @[executor.scala 290:56]
  wire [7:0] _GEN_3390 = 8'h0 < length_2 ? _GEN_3294 : _GEN_3198; // @[executor.scala 290:56]
  wire [7:0] _GEN_3391 = 8'h0 < length_2 ? _GEN_3295 : _GEN_3199; // @[executor.scala 290:56]
  wire [7:0] _GEN_3392 = 8'h0 < length_2 ? _GEN_3296 : _GEN_3200; // @[executor.scala 290:56]
  wire [7:0] _GEN_3393 = 8'h0 < length_2 ? _GEN_3297 : _GEN_3201; // @[executor.scala 290:56]
  wire [7:0] _GEN_3394 = 8'h0 < length_2 ? _GEN_3298 : _GEN_3202; // @[executor.scala 290:56]
  wire [7:0] _GEN_3395 = 8'h0 < length_2 ? _GEN_3299 : _GEN_3203; // @[executor.scala 290:56]
  wire [7:0] _GEN_3396 = 8'h0 < length_2 ? _GEN_3300 : _GEN_3204; // @[executor.scala 290:56]
  wire [7:0] _GEN_3397 = 8'h0 < length_2 ? _GEN_3301 : _GEN_3205; // @[executor.scala 290:56]
  wire [7:0] _GEN_3398 = 8'h0 < length_2 ? _GEN_3302 : _GEN_3206; // @[executor.scala 290:56]
  wire [7:0] _GEN_3399 = 8'h0 < length_2 ? _GEN_3303 : _GEN_3207; // @[executor.scala 290:56]
  wire [7:0] _GEN_3400 = 8'h0 < length_2 ? _GEN_3304 : _GEN_3208; // @[executor.scala 290:56]
  wire [7:0] _GEN_3401 = 8'h0 < length_2 ? _GEN_3305 : _GEN_3209; // @[executor.scala 290:56]
  wire [7:0] _GEN_3402 = 8'h0 < length_2 ? _GEN_3306 : _GEN_3210; // @[executor.scala 290:56]
  wire [7:0] _GEN_3403 = 8'h0 < length_2 ? _GEN_3307 : _GEN_3211; // @[executor.scala 290:56]
  wire [7:0] _GEN_3404 = 8'h0 < length_2 ? _GEN_3308 : _GEN_3212; // @[executor.scala 290:56]
  wire [7:0] _GEN_3405 = 8'h0 < length_2 ? _GEN_3309 : _GEN_3213; // @[executor.scala 290:56]
  wire [7:0] _GEN_3406 = 8'h0 < length_2 ? _GEN_3310 : _GEN_3214; // @[executor.scala 290:56]
  wire [7:0] _GEN_3407 = 8'h0 < length_2 ? _GEN_3311 : _GEN_3215; // @[executor.scala 290:56]
  wire [7:0] _GEN_3408 = 8'h0 < length_2 ? _GEN_3312 : _GEN_3216; // @[executor.scala 290:56]
  wire [7:0] _GEN_3409 = 8'h0 < length_2 ? _GEN_3313 : _GEN_3217; // @[executor.scala 290:56]
  wire [7:0] _GEN_3410 = 8'h0 < length_2 ? _GEN_3314 : _GEN_3218; // @[executor.scala 290:56]
  wire [7:0] _GEN_3411 = 8'h0 < length_2 ? _GEN_3315 : _GEN_3219; // @[executor.scala 290:56]
  wire [7:0] _GEN_3412 = 8'h0 < length_2 ? _GEN_3316 : _GEN_3220; // @[executor.scala 290:56]
  wire [7:0] _GEN_3413 = 8'h0 < length_2 ? _GEN_3317 : _GEN_3221; // @[executor.scala 290:56]
  wire [7:0] _GEN_3414 = 8'h0 < length_2 ? _GEN_3318 : _GEN_3222; // @[executor.scala 290:56]
  wire [7:0] _GEN_3415 = 8'h0 < length_2 ? _GEN_3319 : _GEN_3223; // @[executor.scala 290:56]
  wire [7:0] _GEN_3416 = 8'h0 < length_2 ? _GEN_3320 : _GEN_3224; // @[executor.scala 290:56]
  wire [7:0] _GEN_3417 = 8'h0 < length_2 ? _GEN_3321 : _GEN_3225; // @[executor.scala 290:56]
  wire [7:0] _GEN_3418 = 8'h0 < length_2 ? _GEN_3322 : _GEN_3226; // @[executor.scala 290:56]
  wire [7:0] _GEN_3419 = 8'h0 < length_2 ? _GEN_3323 : _GEN_3227; // @[executor.scala 290:56]
  wire [7:0] _GEN_3420 = 8'h0 < length_2 ? _GEN_3324 : _GEN_3228; // @[executor.scala 290:56]
  wire [7:0] _GEN_3421 = 8'h0 < length_2 ? _GEN_3325 : _GEN_3229; // @[executor.scala 290:56]
  wire [7:0] _GEN_3422 = 8'h0 < length_2 ? _GEN_3326 : _GEN_3230; // @[executor.scala 290:56]
  wire [7:0] _GEN_3423 = 8'h0 < length_2 ? _GEN_3327 : _GEN_3231; // @[executor.scala 290:56]
  wire [7:0] _GEN_3424 = 8'h0 < length_2 ? _GEN_3328 : _GEN_3232; // @[executor.scala 290:56]
  wire [7:0] _GEN_3425 = 8'h0 < length_2 ? _GEN_3329 : _GEN_3233; // @[executor.scala 290:56]
  wire [7:0] _GEN_3426 = 8'h0 < length_2 ? _GEN_3330 : _GEN_3234; // @[executor.scala 290:56]
  wire [7:0] _GEN_3427 = 8'h0 < length_2 ? _GEN_3331 : _GEN_3235; // @[executor.scala 290:56]
  wire [7:0] _GEN_3428 = 8'h0 < length_2 ? _GEN_3332 : _GEN_3236; // @[executor.scala 290:56]
  wire [7:0] _GEN_3429 = 8'h0 < length_2 ? _GEN_3333 : _GEN_3237; // @[executor.scala 290:56]
  wire [7:0] _GEN_3430 = 8'h0 < length_2 ? _GEN_3334 : _GEN_3238; // @[executor.scala 290:56]
  wire [7:0] _GEN_3431 = 8'h0 < length_2 ? _GEN_3335 : _GEN_3239; // @[executor.scala 290:56]
  wire [7:0] _GEN_3432 = 8'h0 < length_2 ? _GEN_3336 : _GEN_3240; // @[executor.scala 290:56]
  wire [7:0] _GEN_3433 = 8'h0 < length_2 ? _GEN_3337 : _GEN_3241; // @[executor.scala 290:56]
  wire [7:0] _GEN_3434 = 8'h0 < length_2 ? _GEN_3338 : _GEN_3242; // @[executor.scala 290:56]
  wire [7:0] _GEN_3435 = 8'h0 < length_2 ? _GEN_3339 : _GEN_3243; // @[executor.scala 290:56]
  wire [7:0] _GEN_3436 = 8'h0 < length_2 ? _GEN_3340 : _GEN_3244; // @[executor.scala 290:56]
  wire [7:0] _GEN_3437 = 8'h0 < length_2 ? _GEN_3341 : _GEN_3245; // @[executor.scala 290:56]
  wire [7:0] _GEN_3438 = 8'h0 < length_2 ? _GEN_3342 : _GEN_3246; // @[executor.scala 290:56]
  wire [7:0] _GEN_3439 = 8'h0 < length_2 ? _GEN_3343 : _GEN_3247; // @[executor.scala 290:56]
  wire [7:0] _GEN_3440 = 8'h0 < length_2 ? _GEN_3344 : _GEN_3248; // @[executor.scala 290:56]
  wire [7:0] _GEN_3441 = 8'h0 < length_2 ? _GEN_3345 : _GEN_3249; // @[executor.scala 290:56]
  wire [7:0] _GEN_3442 = 8'h0 < length_2 ? _GEN_3346 : _GEN_3250; // @[executor.scala 290:56]
  wire [7:0] _GEN_3443 = 8'h0 < length_2 ? _GEN_3347 : _GEN_3251; // @[executor.scala 290:56]
  wire [7:0] _GEN_3444 = 8'h0 < length_2 ? _GEN_3348 : _GEN_3252; // @[executor.scala 290:56]
  wire [7:0] _GEN_3445 = 8'h0 < length_2 ? _GEN_3349 : _GEN_3253; // @[executor.scala 290:56]
  wire [7:0] _GEN_3446 = 8'h0 < length_2 ? _GEN_3350 : _GEN_3254; // @[executor.scala 290:56]
  wire [7:0] _GEN_3447 = 8'h0 < length_2 ? _GEN_3351 : _GEN_3255; // @[executor.scala 290:56]
  wire [7:0] _GEN_3448 = 8'h0 < length_2 ? _GEN_3352 : _GEN_3256; // @[executor.scala 290:56]
  wire [7:0] _GEN_3449 = 8'h0 < length_2 ? _GEN_3353 : _GEN_3257; // @[executor.scala 290:56]
  wire [7:0] _GEN_3450 = 8'h0 < length_2 ? _GEN_3354 : _GEN_3258; // @[executor.scala 290:56]
  wire [7:0] _GEN_3451 = 8'h0 < length_2 ? _GEN_3355 : _GEN_3259; // @[executor.scala 290:56]
  wire [7:0] _GEN_3452 = 8'h0 < length_2 ? _GEN_3356 : _GEN_3260; // @[executor.scala 290:56]
  wire [7:0] _GEN_3453 = 8'h0 < length_2 ? _GEN_3357 : _GEN_3261; // @[executor.scala 290:56]
  wire [7:0] _GEN_3454 = 8'h0 < length_2 ? _GEN_3358 : _GEN_3262; // @[executor.scala 290:56]
  wire [7:0] _GEN_3455 = 8'h0 < length_2 ? _GEN_3359 : _GEN_3263; // @[executor.scala 290:56]
  wire [7:0] _GEN_3456 = 8'h0 < length_2 ? _GEN_3360 : _GEN_3264; // @[executor.scala 290:56]
  wire [7:0] _GEN_3457 = 8'h0 < length_2 ? _GEN_3361 : _GEN_3265; // @[executor.scala 290:56]
  wire [7:0] field_byte_17 = field_2[55:48]; // @[executor.scala 287:53]
  wire [7:0] total_offset_17 = offset_2 + 8'h1; // @[executor.scala 289:53]
  wire [7:0] _GEN_3458 = 7'h0 == total_offset_17[6:0] ? field_byte_17 : _GEN_3362; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3459 = 7'h1 == total_offset_17[6:0] ? field_byte_17 : _GEN_3363; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3460 = 7'h2 == total_offset_17[6:0] ? field_byte_17 : _GEN_3364; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3461 = 7'h3 == total_offset_17[6:0] ? field_byte_17 : _GEN_3365; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3462 = 7'h4 == total_offset_17[6:0] ? field_byte_17 : _GEN_3366; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3463 = 7'h5 == total_offset_17[6:0] ? field_byte_17 : _GEN_3367; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3464 = 7'h6 == total_offset_17[6:0] ? field_byte_17 : _GEN_3368; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3465 = 7'h7 == total_offset_17[6:0] ? field_byte_17 : _GEN_3369; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3466 = 7'h8 == total_offset_17[6:0] ? field_byte_17 : _GEN_3370; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3467 = 7'h9 == total_offset_17[6:0] ? field_byte_17 : _GEN_3371; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3468 = 7'ha == total_offset_17[6:0] ? field_byte_17 : _GEN_3372; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3469 = 7'hb == total_offset_17[6:0] ? field_byte_17 : _GEN_3373; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3470 = 7'hc == total_offset_17[6:0] ? field_byte_17 : _GEN_3374; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3471 = 7'hd == total_offset_17[6:0] ? field_byte_17 : _GEN_3375; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3472 = 7'he == total_offset_17[6:0] ? field_byte_17 : _GEN_3376; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3473 = 7'hf == total_offset_17[6:0] ? field_byte_17 : _GEN_3377; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3474 = 7'h10 == total_offset_17[6:0] ? field_byte_17 : _GEN_3378; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3475 = 7'h11 == total_offset_17[6:0] ? field_byte_17 : _GEN_3379; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3476 = 7'h12 == total_offset_17[6:0] ? field_byte_17 : _GEN_3380; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3477 = 7'h13 == total_offset_17[6:0] ? field_byte_17 : _GEN_3381; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3478 = 7'h14 == total_offset_17[6:0] ? field_byte_17 : _GEN_3382; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3479 = 7'h15 == total_offset_17[6:0] ? field_byte_17 : _GEN_3383; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3480 = 7'h16 == total_offset_17[6:0] ? field_byte_17 : _GEN_3384; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3481 = 7'h17 == total_offset_17[6:0] ? field_byte_17 : _GEN_3385; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3482 = 7'h18 == total_offset_17[6:0] ? field_byte_17 : _GEN_3386; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3483 = 7'h19 == total_offset_17[6:0] ? field_byte_17 : _GEN_3387; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3484 = 7'h1a == total_offset_17[6:0] ? field_byte_17 : _GEN_3388; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3485 = 7'h1b == total_offset_17[6:0] ? field_byte_17 : _GEN_3389; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3486 = 7'h1c == total_offset_17[6:0] ? field_byte_17 : _GEN_3390; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3487 = 7'h1d == total_offset_17[6:0] ? field_byte_17 : _GEN_3391; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3488 = 7'h1e == total_offset_17[6:0] ? field_byte_17 : _GEN_3392; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3489 = 7'h1f == total_offset_17[6:0] ? field_byte_17 : _GEN_3393; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3490 = 7'h20 == total_offset_17[6:0] ? field_byte_17 : _GEN_3394; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3491 = 7'h21 == total_offset_17[6:0] ? field_byte_17 : _GEN_3395; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3492 = 7'h22 == total_offset_17[6:0] ? field_byte_17 : _GEN_3396; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3493 = 7'h23 == total_offset_17[6:0] ? field_byte_17 : _GEN_3397; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3494 = 7'h24 == total_offset_17[6:0] ? field_byte_17 : _GEN_3398; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3495 = 7'h25 == total_offset_17[6:0] ? field_byte_17 : _GEN_3399; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3496 = 7'h26 == total_offset_17[6:0] ? field_byte_17 : _GEN_3400; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3497 = 7'h27 == total_offset_17[6:0] ? field_byte_17 : _GEN_3401; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3498 = 7'h28 == total_offset_17[6:0] ? field_byte_17 : _GEN_3402; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3499 = 7'h29 == total_offset_17[6:0] ? field_byte_17 : _GEN_3403; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3500 = 7'h2a == total_offset_17[6:0] ? field_byte_17 : _GEN_3404; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3501 = 7'h2b == total_offset_17[6:0] ? field_byte_17 : _GEN_3405; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3502 = 7'h2c == total_offset_17[6:0] ? field_byte_17 : _GEN_3406; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3503 = 7'h2d == total_offset_17[6:0] ? field_byte_17 : _GEN_3407; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3504 = 7'h2e == total_offset_17[6:0] ? field_byte_17 : _GEN_3408; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3505 = 7'h2f == total_offset_17[6:0] ? field_byte_17 : _GEN_3409; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3506 = 7'h30 == total_offset_17[6:0] ? field_byte_17 : _GEN_3410; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3507 = 7'h31 == total_offset_17[6:0] ? field_byte_17 : _GEN_3411; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3508 = 7'h32 == total_offset_17[6:0] ? field_byte_17 : _GEN_3412; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3509 = 7'h33 == total_offset_17[6:0] ? field_byte_17 : _GEN_3413; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3510 = 7'h34 == total_offset_17[6:0] ? field_byte_17 : _GEN_3414; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3511 = 7'h35 == total_offset_17[6:0] ? field_byte_17 : _GEN_3415; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3512 = 7'h36 == total_offset_17[6:0] ? field_byte_17 : _GEN_3416; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3513 = 7'h37 == total_offset_17[6:0] ? field_byte_17 : _GEN_3417; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3514 = 7'h38 == total_offset_17[6:0] ? field_byte_17 : _GEN_3418; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3515 = 7'h39 == total_offset_17[6:0] ? field_byte_17 : _GEN_3419; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3516 = 7'h3a == total_offset_17[6:0] ? field_byte_17 : _GEN_3420; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3517 = 7'h3b == total_offset_17[6:0] ? field_byte_17 : _GEN_3421; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3518 = 7'h3c == total_offset_17[6:0] ? field_byte_17 : _GEN_3422; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3519 = 7'h3d == total_offset_17[6:0] ? field_byte_17 : _GEN_3423; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3520 = 7'h3e == total_offset_17[6:0] ? field_byte_17 : _GEN_3424; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3521 = 7'h3f == total_offset_17[6:0] ? field_byte_17 : _GEN_3425; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3522 = 7'h40 == total_offset_17[6:0] ? field_byte_17 : _GEN_3426; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3523 = 7'h41 == total_offset_17[6:0] ? field_byte_17 : _GEN_3427; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3524 = 7'h42 == total_offset_17[6:0] ? field_byte_17 : _GEN_3428; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3525 = 7'h43 == total_offset_17[6:0] ? field_byte_17 : _GEN_3429; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3526 = 7'h44 == total_offset_17[6:0] ? field_byte_17 : _GEN_3430; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3527 = 7'h45 == total_offset_17[6:0] ? field_byte_17 : _GEN_3431; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3528 = 7'h46 == total_offset_17[6:0] ? field_byte_17 : _GEN_3432; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3529 = 7'h47 == total_offset_17[6:0] ? field_byte_17 : _GEN_3433; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3530 = 7'h48 == total_offset_17[6:0] ? field_byte_17 : _GEN_3434; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3531 = 7'h49 == total_offset_17[6:0] ? field_byte_17 : _GEN_3435; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3532 = 7'h4a == total_offset_17[6:0] ? field_byte_17 : _GEN_3436; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3533 = 7'h4b == total_offset_17[6:0] ? field_byte_17 : _GEN_3437; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3534 = 7'h4c == total_offset_17[6:0] ? field_byte_17 : _GEN_3438; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3535 = 7'h4d == total_offset_17[6:0] ? field_byte_17 : _GEN_3439; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3536 = 7'h4e == total_offset_17[6:0] ? field_byte_17 : _GEN_3440; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3537 = 7'h4f == total_offset_17[6:0] ? field_byte_17 : _GEN_3441; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3538 = 7'h50 == total_offset_17[6:0] ? field_byte_17 : _GEN_3442; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3539 = 7'h51 == total_offset_17[6:0] ? field_byte_17 : _GEN_3443; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3540 = 7'h52 == total_offset_17[6:0] ? field_byte_17 : _GEN_3444; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3541 = 7'h53 == total_offset_17[6:0] ? field_byte_17 : _GEN_3445; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3542 = 7'h54 == total_offset_17[6:0] ? field_byte_17 : _GEN_3446; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3543 = 7'h55 == total_offset_17[6:0] ? field_byte_17 : _GEN_3447; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3544 = 7'h56 == total_offset_17[6:0] ? field_byte_17 : _GEN_3448; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3545 = 7'h57 == total_offset_17[6:0] ? field_byte_17 : _GEN_3449; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3546 = 7'h58 == total_offset_17[6:0] ? field_byte_17 : _GEN_3450; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3547 = 7'h59 == total_offset_17[6:0] ? field_byte_17 : _GEN_3451; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3548 = 7'h5a == total_offset_17[6:0] ? field_byte_17 : _GEN_3452; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3549 = 7'h5b == total_offset_17[6:0] ? field_byte_17 : _GEN_3453; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3550 = 7'h5c == total_offset_17[6:0] ? field_byte_17 : _GEN_3454; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3551 = 7'h5d == total_offset_17[6:0] ? field_byte_17 : _GEN_3455; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3552 = 7'h5e == total_offset_17[6:0] ? field_byte_17 : _GEN_3456; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3553 = 7'h5f == total_offset_17[6:0] ? field_byte_17 : _GEN_3457; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3554 = 8'h1 < length_2 ? _GEN_3458 : _GEN_3362; // @[executor.scala 290:56]
  wire [7:0] _GEN_3555 = 8'h1 < length_2 ? _GEN_3459 : _GEN_3363; // @[executor.scala 290:56]
  wire [7:0] _GEN_3556 = 8'h1 < length_2 ? _GEN_3460 : _GEN_3364; // @[executor.scala 290:56]
  wire [7:0] _GEN_3557 = 8'h1 < length_2 ? _GEN_3461 : _GEN_3365; // @[executor.scala 290:56]
  wire [7:0] _GEN_3558 = 8'h1 < length_2 ? _GEN_3462 : _GEN_3366; // @[executor.scala 290:56]
  wire [7:0] _GEN_3559 = 8'h1 < length_2 ? _GEN_3463 : _GEN_3367; // @[executor.scala 290:56]
  wire [7:0] _GEN_3560 = 8'h1 < length_2 ? _GEN_3464 : _GEN_3368; // @[executor.scala 290:56]
  wire [7:0] _GEN_3561 = 8'h1 < length_2 ? _GEN_3465 : _GEN_3369; // @[executor.scala 290:56]
  wire [7:0] _GEN_3562 = 8'h1 < length_2 ? _GEN_3466 : _GEN_3370; // @[executor.scala 290:56]
  wire [7:0] _GEN_3563 = 8'h1 < length_2 ? _GEN_3467 : _GEN_3371; // @[executor.scala 290:56]
  wire [7:0] _GEN_3564 = 8'h1 < length_2 ? _GEN_3468 : _GEN_3372; // @[executor.scala 290:56]
  wire [7:0] _GEN_3565 = 8'h1 < length_2 ? _GEN_3469 : _GEN_3373; // @[executor.scala 290:56]
  wire [7:0] _GEN_3566 = 8'h1 < length_2 ? _GEN_3470 : _GEN_3374; // @[executor.scala 290:56]
  wire [7:0] _GEN_3567 = 8'h1 < length_2 ? _GEN_3471 : _GEN_3375; // @[executor.scala 290:56]
  wire [7:0] _GEN_3568 = 8'h1 < length_2 ? _GEN_3472 : _GEN_3376; // @[executor.scala 290:56]
  wire [7:0] _GEN_3569 = 8'h1 < length_2 ? _GEN_3473 : _GEN_3377; // @[executor.scala 290:56]
  wire [7:0] _GEN_3570 = 8'h1 < length_2 ? _GEN_3474 : _GEN_3378; // @[executor.scala 290:56]
  wire [7:0] _GEN_3571 = 8'h1 < length_2 ? _GEN_3475 : _GEN_3379; // @[executor.scala 290:56]
  wire [7:0] _GEN_3572 = 8'h1 < length_2 ? _GEN_3476 : _GEN_3380; // @[executor.scala 290:56]
  wire [7:0] _GEN_3573 = 8'h1 < length_2 ? _GEN_3477 : _GEN_3381; // @[executor.scala 290:56]
  wire [7:0] _GEN_3574 = 8'h1 < length_2 ? _GEN_3478 : _GEN_3382; // @[executor.scala 290:56]
  wire [7:0] _GEN_3575 = 8'h1 < length_2 ? _GEN_3479 : _GEN_3383; // @[executor.scala 290:56]
  wire [7:0] _GEN_3576 = 8'h1 < length_2 ? _GEN_3480 : _GEN_3384; // @[executor.scala 290:56]
  wire [7:0] _GEN_3577 = 8'h1 < length_2 ? _GEN_3481 : _GEN_3385; // @[executor.scala 290:56]
  wire [7:0] _GEN_3578 = 8'h1 < length_2 ? _GEN_3482 : _GEN_3386; // @[executor.scala 290:56]
  wire [7:0] _GEN_3579 = 8'h1 < length_2 ? _GEN_3483 : _GEN_3387; // @[executor.scala 290:56]
  wire [7:0] _GEN_3580 = 8'h1 < length_2 ? _GEN_3484 : _GEN_3388; // @[executor.scala 290:56]
  wire [7:0] _GEN_3581 = 8'h1 < length_2 ? _GEN_3485 : _GEN_3389; // @[executor.scala 290:56]
  wire [7:0] _GEN_3582 = 8'h1 < length_2 ? _GEN_3486 : _GEN_3390; // @[executor.scala 290:56]
  wire [7:0] _GEN_3583 = 8'h1 < length_2 ? _GEN_3487 : _GEN_3391; // @[executor.scala 290:56]
  wire [7:0] _GEN_3584 = 8'h1 < length_2 ? _GEN_3488 : _GEN_3392; // @[executor.scala 290:56]
  wire [7:0] _GEN_3585 = 8'h1 < length_2 ? _GEN_3489 : _GEN_3393; // @[executor.scala 290:56]
  wire [7:0] _GEN_3586 = 8'h1 < length_2 ? _GEN_3490 : _GEN_3394; // @[executor.scala 290:56]
  wire [7:0] _GEN_3587 = 8'h1 < length_2 ? _GEN_3491 : _GEN_3395; // @[executor.scala 290:56]
  wire [7:0] _GEN_3588 = 8'h1 < length_2 ? _GEN_3492 : _GEN_3396; // @[executor.scala 290:56]
  wire [7:0] _GEN_3589 = 8'h1 < length_2 ? _GEN_3493 : _GEN_3397; // @[executor.scala 290:56]
  wire [7:0] _GEN_3590 = 8'h1 < length_2 ? _GEN_3494 : _GEN_3398; // @[executor.scala 290:56]
  wire [7:0] _GEN_3591 = 8'h1 < length_2 ? _GEN_3495 : _GEN_3399; // @[executor.scala 290:56]
  wire [7:0] _GEN_3592 = 8'h1 < length_2 ? _GEN_3496 : _GEN_3400; // @[executor.scala 290:56]
  wire [7:0] _GEN_3593 = 8'h1 < length_2 ? _GEN_3497 : _GEN_3401; // @[executor.scala 290:56]
  wire [7:0] _GEN_3594 = 8'h1 < length_2 ? _GEN_3498 : _GEN_3402; // @[executor.scala 290:56]
  wire [7:0] _GEN_3595 = 8'h1 < length_2 ? _GEN_3499 : _GEN_3403; // @[executor.scala 290:56]
  wire [7:0] _GEN_3596 = 8'h1 < length_2 ? _GEN_3500 : _GEN_3404; // @[executor.scala 290:56]
  wire [7:0] _GEN_3597 = 8'h1 < length_2 ? _GEN_3501 : _GEN_3405; // @[executor.scala 290:56]
  wire [7:0] _GEN_3598 = 8'h1 < length_2 ? _GEN_3502 : _GEN_3406; // @[executor.scala 290:56]
  wire [7:0] _GEN_3599 = 8'h1 < length_2 ? _GEN_3503 : _GEN_3407; // @[executor.scala 290:56]
  wire [7:0] _GEN_3600 = 8'h1 < length_2 ? _GEN_3504 : _GEN_3408; // @[executor.scala 290:56]
  wire [7:0] _GEN_3601 = 8'h1 < length_2 ? _GEN_3505 : _GEN_3409; // @[executor.scala 290:56]
  wire [7:0] _GEN_3602 = 8'h1 < length_2 ? _GEN_3506 : _GEN_3410; // @[executor.scala 290:56]
  wire [7:0] _GEN_3603 = 8'h1 < length_2 ? _GEN_3507 : _GEN_3411; // @[executor.scala 290:56]
  wire [7:0] _GEN_3604 = 8'h1 < length_2 ? _GEN_3508 : _GEN_3412; // @[executor.scala 290:56]
  wire [7:0] _GEN_3605 = 8'h1 < length_2 ? _GEN_3509 : _GEN_3413; // @[executor.scala 290:56]
  wire [7:0] _GEN_3606 = 8'h1 < length_2 ? _GEN_3510 : _GEN_3414; // @[executor.scala 290:56]
  wire [7:0] _GEN_3607 = 8'h1 < length_2 ? _GEN_3511 : _GEN_3415; // @[executor.scala 290:56]
  wire [7:0] _GEN_3608 = 8'h1 < length_2 ? _GEN_3512 : _GEN_3416; // @[executor.scala 290:56]
  wire [7:0] _GEN_3609 = 8'h1 < length_2 ? _GEN_3513 : _GEN_3417; // @[executor.scala 290:56]
  wire [7:0] _GEN_3610 = 8'h1 < length_2 ? _GEN_3514 : _GEN_3418; // @[executor.scala 290:56]
  wire [7:0] _GEN_3611 = 8'h1 < length_2 ? _GEN_3515 : _GEN_3419; // @[executor.scala 290:56]
  wire [7:0] _GEN_3612 = 8'h1 < length_2 ? _GEN_3516 : _GEN_3420; // @[executor.scala 290:56]
  wire [7:0] _GEN_3613 = 8'h1 < length_2 ? _GEN_3517 : _GEN_3421; // @[executor.scala 290:56]
  wire [7:0] _GEN_3614 = 8'h1 < length_2 ? _GEN_3518 : _GEN_3422; // @[executor.scala 290:56]
  wire [7:0] _GEN_3615 = 8'h1 < length_2 ? _GEN_3519 : _GEN_3423; // @[executor.scala 290:56]
  wire [7:0] _GEN_3616 = 8'h1 < length_2 ? _GEN_3520 : _GEN_3424; // @[executor.scala 290:56]
  wire [7:0] _GEN_3617 = 8'h1 < length_2 ? _GEN_3521 : _GEN_3425; // @[executor.scala 290:56]
  wire [7:0] _GEN_3618 = 8'h1 < length_2 ? _GEN_3522 : _GEN_3426; // @[executor.scala 290:56]
  wire [7:0] _GEN_3619 = 8'h1 < length_2 ? _GEN_3523 : _GEN_3427; // @[executor.scala 290:56]
  wire [7:0] _GEN_3620 = 8'h1 < length_2 ? _GEN_3524 : _GEN_3428; // @[executor.scala 290:56]
  wire [7:0] _GEN_3621 = 8'h1 < length_2 ? _GEN_3525 : _GEN_3429; // @[executor.scala 290:56]
  wire [7:0] _GEN_3622 = 8'h1 < length_2 ? _GEN_3526 : _GEN_3430; // @[executor.scala 290:56]
  wire [7:0] _GEN_3623 = 8'h1 < length_2 ? _GEN_3527 : _GEN_3431; // @[executor.scala 290:56]
  wire [7:0] _GEN_3624 = 8'h1 < length_2 ? _GEN_3528 : _GEN_3432; // @[executor.scala 290:56]
  wire [7:0] _GEN_3625 = 8'h1 < length_2 ? _GEN_3529 : _GEN_3433; // @[executor.scala 290:56]
  wire [7:0] _GEN_3626 = 8'h1 < length_2 ? _GEN_3530 : _GEN_3434; // @[executor.scala 290:56]
  wire [7:0] _GEN_3627 = 8'h1 < length_2 ? _GEN_3531 : _GEN_3435; // @[executor.scala 290:56]
  wire [7:0] _GEN_3628 = 8'h1 < length_2 ? _GEN_3532 : _GEN_3436; // @[executor.scala 290:56]
  wire [7:0] _GEN_3629 = 8'h1 < length_2 ? _GEN_3533 : _GEN_3437; // @[executor.scala 290:56]
  wire [7:0] _GEN_3630 = 8'h1 < length_2 ? _GEN_3534 : _GEN_3438; // @[executor.scala 290:56]
  wire [7:0] _GEN_3631 = 8'h1 < length_2 ? _GEN_3535 : _GEN_3439; // @[executor.scala 290:56]
  wire [7:0] _GEN_3632 = 8'h1 < length_2 ? _GEN_3536 : _GEN_3440; // @[executor.scala 290:56]
  wire [7:0] _GEN_3633 = 8'h1 < length_2 ? _GEN_3537 : _GEN_3441; // @[executor.scala 290:56]
  wire [7:0] _GEN_3634 = 8'h1 < length_2 ? _GEN_3538 : _GEN_3442; // @[executor.scala 290:56]
  wire [7:0] _GEN_3635 = 8'h1 < length_2 ? _GEN_3539 : _GEN_3443; // @[executor.scala 290:56]
  wire [7:0] _GEN_3636 = 8'h1 < length_2 ? _GEN_3540 : _GEN_3444; // @[executor.scala 290:56]
  wire [7:0] _GEN_3637 = 8'h1 < length_2 ? _GEN_3541 : _GEN_3445; // @[executor.scala 290:56]
  wire [7:0] _GEN_3638 = 8'h1 < length_2 ? _GEN_3542 : _GEN_3446; // @[executor.scala 290:56]
  wire [7:0] _GEN_3639 = 8'h1 < length_2 ? _GEN_3543 : _GEN_3447; // @[executor.scala 290:56]
  wire [7:0] _GEN_3640 = 8'h1 < length_2 ? _GEN_3544 : _GEN_3448; // @[executor.scala 290:56]
  wire [7:0] _GEN_3641 = 8'h1 < length_2 ? _GEN_3545 : _GEN_3449; // @[executor.scala 290:56]
  wire [7:0] _GEN_3642 = 8'h1 < length_2 ? _GEN_3546 : _GEN_3450; // @[executor.scala 290:56]
  wire [7:0] _GEN_3643 = 8'h1 < length_2 ? _GEN_3547 : _GEN_3451; // @[executor.scala 290:56]
  wire [7:0] _GEN_3644 = 8'h1 < length_2 ? _GEN_3548 : _GEN_3452; // @[executor.scala 290:56]
  wire [7:0] _GEN_3645 = 8'h1 < length_2 ? _GEN_3549 : _GEN_3453; // @[executor.scala 290:56]
  wire [7:0] _GEN_3646 = 8'h1 < length_2 ? _GEN_3550 : _GEN_3454; // @[executor.scala 290:56]
  wire [7:0] _GEN_3647 = 8'h1 < length_2 ? _GEN_3551 : _GEN_3455; // @[executor.scala 290:56]
  wire [7:0] _GEN_3648 = 8'h1 < length_2 ? _GEN_3552 : _GEN_3456; // @[executor.scala 290:56]
  wire [7:0] _GEN_3649 = 8'h1 < length_2 ? _GEN_3553 : _GEN_3457; // @[executor.scala 290:56]
  wire [7:0] field_byte_18 = field_2[47:40]; // @[executor.scala 287:53]
  wire [7:0] total_offset_18 = offset_2 + 8'h2; // @[executor.scala 289:53]
  wire [7:0] _GEN_3650 = 7'h0 == total_offset_18[6:0] ? field_byte_18 : _GEN_3554; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3651 = 7'h1 == total_offset_18[6:0] ? field_byte_18 : _GEN_3555; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3652 = 7'h2 == total_offset_18[6:0] ? field_byte_18 : _GEN_3556; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3653 = 7'h3 == total_offset_18[6:0] ? field_byte_18 : _GEN_3557; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3654 = 7'h4 == total_offset_18[6:0] ? field_byte_18 : _GEN_3558; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3655 = 7'h5 == total_offset_18[6:0] ? field_byte_18 : _GEN_3559; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3656 = 7'h6 == total_offset_18[6:0] ? field_byte_18 : _GEN_3560; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3657 = 7'h7 == total_offset_18[6:0] ? field_byte_18 : _GEN_3561; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3658 = 7'h8 == total_offset_18[6:0] ? field_byte_18 : _GEN_3562; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3659 = 7'h9 == total_offset_18[6:0] ? field_byte_18 : _GEN_3563; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3660 = 7'ha == total_offset_18[6:0] ? field_byte_18 : _GEN_3564; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3661 = 7'hb == total_offset_18[6:0] ? field_byte_18 : _GEN_3565; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3662 = 7'hc == total_offset_18[6:0] ? field_byte_18 : _GEN_3566; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3663 = 7'hd == total_offset_18[6:0] ? field_byte_18 : _GEN_3567; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3664 = 7'he == total_offset_18[6:0] ? field_byte_18 : _GEN_3568; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3665 = 7'hf == total_offset_18[6:0] ? field_byte_18 : _GEN_3569; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3666 = 7'h10 == total_offset_18[6:0] ? field_byte_18 : _GEN_3570; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3667 = 7'h11 == total_offset_18[6:0] ? field_byte_18 : _GEN_3571; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3668 = 7'h12 == total_offset_18[6:0] ? field_byte_18 : _GEN_3572; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3669 = 7'h13 == total_offset_18[6:0] ? field_byte_18 : _GEN_3573; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3670 = 7'h14 == total_offset_18[6:0] ? field_byte_18 : _GEN_3574; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3671 = 7'h15 == total_offset_18[6:0] ? field_byte_18 : _GEN_3575; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3672 = 7'h16 == total_offset_18[6:0] ? field_byte_18 : _GEN_3576; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3673 = 7'h17 == total_offset_18[6:0] ? field_byte_18 : _GEN_3577; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3674 = 7'h18 == total_offset_18[6:0] ? field_byte_18 : _GEN_3578; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3675 = 7'h19 == total_offset_18[6:0] ? field_byte_18 : _GEN_3579; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3676 = 7'h1a == total_offset_18[6:0] ? field_byte_18 : _GEN_3580; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3677 = 7'h1b == total_offset_18[6:0] ? field_byte_18 : _GEN_3581; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3678 = 7'h1c == total_offset_18[6:0] ? field_byte_18 : _GEN_3582; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3679 = 7'h1d == total_offset_18[6:0] ? field_byte_18 : _GEN_3583; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3680 = 7'h1e == total_offset_18[6:0] ? field_byte_18 : _GEN_3584; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3681 = 7'h1f == total_offset_18[6:0] ? field_byte_18 : _GEN_3585; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3682 = 7'h20 == total_offset_18[6:0] ? field_byte_18 : _GEN_3586; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3683 = 7'h21 == total_offset_18[6:0] ? field_byte_18 : _GEN_3587; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3684 = 7'h22 == total_offset_18[6:0] ? field_byte_18 : _GEN_3588; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3685 = 7'h23 == total_offset_18[6:0] ? field_byte_18 : _GEN_3589; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3686 = 7'h24 == total_offset_18[6:0] ? field_byte_18 : _GEN_3590; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3687 = 7'h25 == total_offset_18[6:0] ? field_byte_18 : _GEN_3591; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3688 = 7'h26 == total_offset_18[6:0] ? field_byte_18 : _GEN_3592; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3689 = 7'h27 == total_offset_18[6:0] ? field_byte_18 : _GEN_3593; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3690 = 7'h28 == total_offset_18[6:0] ? field_byte_18 : _GEN_3594; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3691 = 7'h29 == total_offset_18[6:0] ? field_byte_18 : _GEN_3595; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3692 = 7'h2a == total_offset_18[6:0] ? field_byte_18 : _GEN_3596; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3693 = 7'h2b == total_offset_18[6:0] ? field_byte_18 : _GEN_3597; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3694 = 7'h2c == total_offset_18[6:0] ? field_byte_18 : _GEN_3598; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3695 = 7'h2d == total_offset_18[6:0] ? field_byte_18 : _GEN_3599; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3696 = 7'h2e == total_offset_18[6:0] ? field_byte_18 : _GEN_3600; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3697 = 7'h2f == total_offset_18[6:0] ? field_byte_18 : _GEN_3601; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3698 = 7'h30 == total_offset_18[6:0] ? field_byte_18 : _GEN_3602; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3699 = 7'h31 == total_offset_18[6:0] ? field_byte_18 : _GEN_3603; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3700 = 7'h32 == total_offset_18[6:0] ? field_byte_18 : _GEN_3604; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3701 = 7'h33 == total_offset_18[6:0] ? field_byte_18 : _GEN_3605; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3702 = 7'h34 == total_offset_18[6:0] ? field_byte_18 : _GEN_3606; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3703 = 7'h35 == total_offset_18[6:0] ? field_byte_18 : _GEN_3607; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3704 = 7'h36 == total_offset_18[6:0] ? field_byte_18 : _GEN_3608; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3705 = 7'h37 == total_offset_18[6:0] ? field_byte_18 : _GEN_3609; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3706 = 7'h38 == total_offset_18[6:0] ? field_byte_18 : _GEN_3610; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3707 = 7'h39 == total_offset_18[6:0] ? field_byte_18 : _GEN_3611; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3708 = 7'h3a == total_offset_18[6:0] ? field_byte_18 : _GEN_3612; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3709 = 7'h3b == total_offset_18[6:0] ? field_byte_18 : _GEN_3613; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3710 = 7'h3c == total_offset_18[6:0] ? field_byte_18 : _GEN_3614; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3711 = 7'h3d == total_offset_18[6:0] ? field_byte_18 : _GEN_3615; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3712 = 7'h3e == total_offset_18[6:0] ? field_byte_18 : _GEN_3616; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3713 = 7'h3f == total_offset_18[6:0] ? field_byte_18 : _GEN_3617; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3714 = 7'h40 == total_offset_18[6:0] ? field_byte_18 : _GEN_3618; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3715 = 7'h41 == total_offset_18[6:0] ? field_byte_18 : _GEN_3619; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3716 = 7'h42 == total_offset_18[6:0] ? field_byte_18 : _GEN_3620; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3717 = 7'h43 == total_offset_18[6:0] ? field_byte_18 : _GEN_3621; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3718 = 7'h44 == total_offset_18[6:0] ? field_byte_18 : _GEN_3622; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3719 = 7'h45 == total_offset_18[6:0] ? field_byte_18 : _GEN_3623; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3720 = 7'h46 == total_offset_18[6:0] ? field_byte_18 : _GEN_3624; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3721 = 7'h47 == total_offset_18[6:0] ? field_byte_18 : _GEN_3625; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3722 = 7'h48 == total_offset_18[6:0] ? field_byte_18 : _GEN_3626; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3723 = 7'h49 == total_offset_18[6:0] ? field_byte_18 : _GEN_3627; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3724 = 7'h4a == total_offset_18[6:0] ? field_byte_18 : _GEN_3628; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3725 = 7'h4b == total_offset_18[6:0] ? field_byte_18 : _GEN_3629; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3726 = 7'h4c == total_offset_18[6:0] ? field_byte_18 : _GEN_3630; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3727 = 7'h4d == total_offset_18[6:0] ? field_byte_18 : _GEN_3631; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3728 = 7'h4e == total_offset_18[6:0] ? field_byte_18 : _GEN_3632; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3729 = 7'h4f == total_offset_18[6:0] ? field_byte_18 : _GEN_3633; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3730 = 7'h50 == total_offset_18[6:0] ? field_byte_18 : _GEN_3634; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3731 = 7'h51 == total_offset_18[6:0] ? field_byte_18 : _GEN_3635; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3732 = 7'h52 == total_offset_18[6:0] ? field_byte_18 : _GEN_3636; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3733 = 7'h53 == total_offset_18[6:0] ? field_byte_18 : _GEN_3637; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3734 = 7'h54 == total_offset_18[6:0] ? field_byte_18 : _GEN_3638; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3735 = 7'h55 == total_offset_18[6:0] ? field_byte_18 : _GEN_3639; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3736 = 7'h56 == total_offset_18[6:0] ? field_byte_18 : _GEN_3640; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3737 = 7'h57 == total_offset_18[6:0] ? field_byte_18 : _GEN_3641; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3738 = 7'h58 == total_offset_18[6:0] ? field_byte_18 : _GEN_3642; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3739 = 7'h59 == total_offset_18[6:0] ? field_byte_18 : _GEN_3643; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3740 = 7'h5a == total_offset_18[6:0] ? field_byte_18 : _GEN_3644; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3741 = 7'h5b == total_offset_18[6:0] ? field_byte_18 : _GEN_3645; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3742 = 7'h5c == total_offset_18[6:0] ? field_byte_18 : _GEN_3646; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3743 = 7'h5d == total_offset_18[6:0] ? field_byte_18 : _GEN_3647; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3744 = 7'h5e == total_offset_18[6:0] ? field_byte_18 : _GEN_3648; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3745 = 7'h5f == total_offset_18[6:0] ? field_byte_18 : _GEN_3649; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3746 = 8'h2 < length_2 ? _GEN_3650 : _GEN_3554; // @[executor.scala 290:56]
  wire [7:0] _GEN_3747 = 8'h2 < length_2 ? _GEN_3651 : _GEN_3555; // @[executor.scala 290:56]
  wire [7:0] _GEN_3748 = 8'h2 < length_2 ? _GEN_3652 : _GEN_3556; // @[executor.scala 290:56]
  wire [7:0] _GEN_3749 = 8'h2 < length_2 ? _GEN_3653 : _GEN_3557; // @[executor.scala 290:56]
  wire [7:0] _GEN_3750 = 8'h2 < length_2 ? _GEN_3654 : _GEN_3558; // @[executor.scala 290:56]
  wire [7:0] _GEN_3751 = 8'h2 < length_2 ? _GEN_3655 : _GEN_3559; // @[executor.scala 290:56]
  wire [7:0] _GEN_3752 = 8'h2 < length_2 ? _GEN_3656 : _GEN_3560; // @[executor.scala 290:56]
  wire [7:0] _GEN_3753 = 8'h2 < length_2 ? _GEN_3657 : _GEN_3561; // @[executor.scala 290:56]
  wire [7:0] _GEN_3754 = 8'h2 < length_2 ? _GEN_3658 : _GEN_3562; // @[executor.scala 290:56]
  wire [7:0] _GEN_3755 = 8'h2 < length_2 ? _GEN_3659 : _GEN_3563; // @[executor.scala 290:56]
  wire [7:0] _GEN_3756 = 8'h2 < length_2 ? _GEN_3660 : _GEN_3564; // @[executor.scala 290:56]
  wire [7:0] _GEN_3757 = 8'h2 < length_2 ? _GEN_3661 : _GEN_3565; // @[executor.scala 290:56]
  wire [7:0] _GEN_3758 = 8'h2 < length_2 ? _GEN_3662 : _GEN_3566; // @[executor.scala 290:56]
  wire [7:0] _GEN_3759 = 8'h2 < length_2 ? _GEN_3663 : _GEN_3567; // @[executor.scala 290:56]
  wire [7:0] _GEN_3760 = 8'h2 < length_2 ? _GEN_3664 : _GEN_3568; // @[executor.scala 290:56]
  wire [7:0] _GEN_3761 = 8'h2 < length_2 ? _GEN_3665 : _GEN_3569; // @[executor.scala 290:56]
  wire [7:0] _GEN_3762 = 8'h2 < length_2 ? _GEN_3666 : _GEN_3570; // @[executor.scala 290:56]
  wire [7:0] _GEN_3763 = 8'h2 < length_2 ? _GEN_3667 : _GEN_3571; // @[executor.scala 290:56]
  wire [7:0] _GEN_3764 = 8'h2 < length_2 ? _GEN_3668 : _GEN_3572; // @[executor.scala 290:56]
  wire [7:0] _GEN_3765 = 8'h2 < length_2 ? _GEN_3669 : _GEN_3573; // @[executor.scala 290:56]
  wire [7:0] _GEN_3766 = 8'h2 < length_2 ? _GEN_3670 : _GEN_3574; // @[executor.scala 290:56]
  wire [7:0] _GEN_3767 = 8'h2 < length_2 ? _GEN_3671 : _GEN_3575; // @[executor.scala 290:56]
  wire [7:0] _GEN_3768 = 8'h2 < length_2 ? _GEN_3672 : _GEN_3576; // @[executor.scala 290:56]
  wire [7:0] _GEN_3769 = 8'h2 < length_2 ? _GEN_3673 : _GEN_3577; // @[executor.scala 290:56]
  wire [7:0] _GEN_3770 = 8'h2 < length_2 ? _GEN_3674 : _GEN_3578; // @[executor.scala 290:56]
  wire [7:0] _GEN_3771 = 8'h2 < length_2 ? _GEN_3675 : _GEN_3579; // @[executor.scala 290:56]
  wire [7:0] _GEN_3772 = 8'h2 < length_2 ? _GEN_3676 : _GEN_3580; // @[executor.scala 290:56]
  wire [7:0] _GEN_3773 = 8'h2 < length_2 ? _GEN_3677 : _GEN_3581; // @[executor.scala 290:56]
  wire [7:0] _GEN_3774 = 8'h2 < length_2 ? _GEN_3678 : _GEN_3582; // @[executor.scala 290:56]
  wire [7:0] _GEN_3775 = 8'h2 < length_2 ? _GEN_3679 : _GEN_3583; // @[executor.scala 290:56]
  wire [7:0] _GEN_3776 = 8'h2 < length_2 ? _GEN_3680 : _GEN_3584; // @[executor.scala 290:56]
  wire [7:0] _GEN_3777 = 8'h2 < length_2 ? _GEN_3681 : _GEN_3585; // @[executor.scala 290:56]
  wire [7:0] _GEN_3778 = 8'h2 < length_2 ? _GEN_3682 : _GEN_3586; // @[executor.scala 290:56]
  wire [7:0] _GEN_3779 = 8'h2 < length_2 ? _GEN_3683 : _GEN_3587; // @[executor.scala 290:56]
  wire [7:0] _GEN_3780 = 8'h2 < length_2 ? _GEN_3684 : _GEN_3588; // @[executor.scala 290:56]
  wire [7:0] _GEN_3781 = 8'h2 < length_2 ? _GEN_3685 : _GEN_3589; // @[executor.scala 290:56]
  wire [7:0] _GEN_3782 = 8'h2 < length_2 ? _GEN_3686 : _GEN_3590; // @[executor.scala 290:56]
  wire [7:0] _GEN_3783 = 8'h2 < length_2 ? _GEN_3687 : _GEN_3591; // @[executor.scala 290:56]
  wire [7:0] _GEN_3784 = 8'h2 < length_2 ? _GEN_3688 : _GEN_3592; // @[executor.scala 290:56]
  wire [7:0] _GEN_3785 = 8'h2 < length_2 ? _GEN_3689 : _GEN_3593; // @[executor.scala 290:56]
  wire [7:0] _GEN_3786 = 8'h2 < length_2 ? _GEN_3690 : _GEN_3594; // @[executor.scala 290:56]
  wire [7:0] _GEN_3787 = 8'h2 < length_2 ? _GEN_3691 : _GEN_3595; // @[executor.scala 290:56]
  wire [7:0] _GEN_3788 = 8'h2 < length_2 ? _GEN_3692 : _GEN_3596; // @[executor.scala 290:56]
  wire [7:0] _GEN_3789 = 8'h2 < length_2 ? _GEN_3693 : _GEN_3597; // @[executor.scala 290:56]
  wire [7:0] _GEN_3790 = 8'h2 < length_2 ? _GEN_3694 : _GEN_3598; // @[executor.scala 290:56]
  wire [7:0] _GEN_3791 = 8'h2 < length_2 ? _GEN_3695 : _GEN_3599; // @[executor.scala 290:56]
  wire [7:0] _GEN_3792 = 8'h2 < length_2 ? _GEN_3696 : _GEN_3600; // @[executor.scala 290:56]
  wire [7:0] _GEN_3793 = 8'h2 < length_2 ? _GEN_3697 : _GEN_3601; // @[executor.scala 290:56]
  wire [7:0] _GEN_3794 = 8'h2 < length_2 ? _GEN_3698 : _GEN_3602; // @[executor.scala 290:56]
  wire [7:0] _GEN_3795 = 8'h2 < length_2 ? _GEN_3699 : _GEN_3603; // @[executor.scala 290:56]
  wire [7:0] _GEN_3796 = 8'h2 < length_2 ? _GEN_3700 : _GEN_3604; // @[executor.scala 290:56]
  wire [7:0] _GEN_3797 = 8'h2 < length_2 ? _GEN_3701 : _GEN_3605; // @[executor.scala 290:56]
  wire [7:0] _GEN_3798 = 8'h2 < length_2 ? _GEN_3702 : _GEN_3606; // @[executor.scala 290:56]
  wire [7:0] _GEN_3799 = 8'h2 < length_2 ? _GEN_3703 : _GEN_3607; // @[executor.scala 290:56]
  wire [7:0] _GEN_3800 = 8'h2 < length_2 ? _GEN_3704 : _GEN_3608; // @[executor.scala 290:56]
  wire [7:0] _GEN_3801 = 8'h2 < length_2 ? _GEN_3705 : _GEN_3609; // @[executor.scala 290:56]
  wire [7:0] _GEN_3802 = 8'h2 < length_2 ? _GEN_3706 : _GEN_3610; // @[executor.scala 290:56]
  wire [7:0] _GEN_3803 = 8'h2 < length_2 ? _GEN_3707 : _GEN_3611; // @[executor.scala 290:56]
  wire [7:0] _GEN_3804 = 8'h2 < length_2 ? _GEN_3708 : _GEN_3612; // @[executor.scala 290:56]
  wire [7:0] _GEN_3805 = 8'h2 < length_2 ? _GEN_3709 : _GEN_3613; // @[executor.scala 290:56]
  wire [7:0] _GEN_3806 = 8'h2 < length_2 ? _GEN_3710 : _GEN_3614; // @[executor.scala 290:56]
  wire [7:0] _GEN_3807 = 8'h2 < length_2 ? _GEN_3711 : _GEN_3615; // @[executor.scala 290:56]
  wire [7:0] _GEN_3808 = 8'h2 < length_2 ? _GEN_3712 : _GEN_3616; // @[executor.scala 290:56]
  wire [7:0] _GEN_3809 = 8'h2 < length_2 ? _GEN_3713 : _GEN_3617; // @[executor.scala 290:56]
  wire [7:0] _GEN_3810 = 8'h2 < length_2 ? _GEN_3714 : _GEN_3618; // @[executor.scala 290:56]
  wire [7:0] _GEN_3811 = 8'h2 < length_2 ? _GEN_3715 : _GEN_3619; // @[executor.scala 290:56]
  wire [7:0] _GEN_3812 = 8'h2 < length_2 ? _GEN_3716 : _GEN_3620; // @[executor.scala 290:56]
  wire [7:0] _GEN_3813 = 8'h2 < length_2 ? _GEN_3717 : _GEN_3621; // @[executor.scala 290:56]
  wire [7:0] _GEN_3814 = 8'h2 < length_2 ? _GEN_3718 : _GEN_3622; // @[executor.scala 290:56]
  wire [7:0] _GEN_3815 = 8'h2 < length_2 ? _GEN_3719 : _GEN_3623; // @[executor.scala 290:56]
  wire [7:0] _GEN_3816 = 8'h2 < length_2 ? _GEN_3720 : _GEN_3624; // @[executor.scala 290:56]
  wire [7:0] _GEN_3817 = 8'h2 < length_2 ? _GEN_3721 : _GEN_3625; // @[executor.scala 290:56]
  wire [7:0] _GEN_3818 = 8'h2 < length_2 ? _GEN_3722 : _GEN_3626; // @[executor.scala 290:56]
  wire [7:0] _GEN_3819 = 8'h2 < length_2 ? _GEN_3723 : _GEN_3627; // @[executor.scala 290:56]
  wire [7:0] _GEN_3820 = 8'h2 < length_2 ? _GEN_3724 : _GEN_3628; // @[executor.scala 290:56]
  wire [7:0] _GEN_3821 = 8'h2 < length_2 ? _GEN_3725 : _GEN_3629; // @[executor.scala 290:56]
  wire [7:0] _GEN_3822 = 8'h2 < length_2 ? _GEN_3726 : _GEN_3630; // @[executor.scala 290:56]
  wire [7:0] _GEN_3823 = 8'h2 < length_2 ? _GEN_3727 : _GEN_3631; // @[executor.scala 290:56]
  wire [7:0] _GEN_3824 = 8'h2 < length_2 ? _GEN_3728 : _GEN_3632; // @[executor.scala 290:56]
  wire [7:0] _GEN_3825 = 8'h2 < length_2 ? _GEN_3729 : _GEN_3633; // @[executor.scala 290:56]
  wire [7:0] _GEN_3826 = 8'h2 < length_2 ? _GEN_3730 : _GEN_3634; // @[executor.scala 290:56]
  wire [7:0] _GEN_3827 = 8'h2 < length_2 ? _GEN_3731 : _GEN_3635; // @[executor.scala 290:56]
  wire [7:0] _GEN_3828 = 8'h2 < length_2 ? _GEN_3732 : _GEN_3636; // @[executor.scala 290:56]
  wire [7:0] _GEN_3829 = 8'h2 < length_2 ? _GEN_3733 : _GEN_3637; // @[executor.scala 290:56]
  wire [7:0] _GEN_3830 = 8'h2 < length_2 ? _GEN_3734 : _GEN_3638; // @[executor.scala 290:56]
  wire [7:0] _GEN_3831 = 8'h2 < length_2 ? _GEN_3735 : _GEN_3639; // @[executor.scala 290:56]
  wire [7:0] _GEN_3832 = 8'h2 < length_2 ? _GEN_3736 : _GEN_3640; // @[executor.scala 290:56]
  wire [7:0] _GEN_3833 = 8'h2 < length_2 ? _GEN_3737 : _GEN_3641; // @[executor.scala 290:56]
  wire [7:0] _GEN_3834 = 8'h2 < length_2 ? _GEN_3738 : _GEN_3642; // @[executor.scala 290:56]
  wire [7:0] _GEN_3835 = 8'h2 < length_2 ? _GEN_3739 : _GEN_3643; // @[executor.scala 290:56]
  wire [7:0] _GEN_3836 = 8'h2 < length_2 ? _GEN_3740 : _GEN_3644; // @[executor.scala 290:56]
  wire [7:0] _GEN_3837 = 8'h2 < length_2 ? _GEN_3741 : _GEN_3645; // @[executor.scala 290:56]
  wire [7:0] _GEN_3838 = 8'h2 < length_2 ? _GEN_3742 : _GEN_3646; // @[executor.scala 290:56]
  wire [7:0] _GEN_3839 = 8'h2 < length_2 ? _GEN_3743 : _GEN_3647; // @[executor.scala 290:56]
  wire [7:0] _GEN_3840 = 8'h2 < length_2 ? _GEN_3744 : _GEN_3648; // @[executor.scala 290:56]
  wire [7:0] _GEN_3841 = 8'h2 < length_2 ? _GEN_3745 : _GEN_3649; // @[executor.scala 290:56]
  wire [7:0] field_byte_19 = field_2[39:32]; // @[executor.scala 287:53]
  wire [7:0] total_offset_19 = offset_2 + 8'h3; // @[executor.scala 289:53]
  wire [7:0] _GEN_3842 = 7'h0 == total_offset_19[6:0] ? field_byte_19 : _GEN_3746; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3843 = 7'h1 == total_offset_19[6:0] ? field_byte_19 : _GEN_3747; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3844 = 7'h2 == total_offset_19[6:0] ? field_byte_19 : _GEN_3748; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3845 = 7'h3 == total_offset_19[6:0] ? field_byte_19 : _GEN_3749; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3846 = 7'h4 == total_offset_19[6:0] ? field_byte_19 : _GEN_3750; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3847 = 7'h5 == total_offset_19[6:0] ? field_byte_19 : _GEN_3751; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3848 = 7'h6 == total_offset_19[6:0] ? field_byte_19 : _GEN_3752; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3849 = 7'h7 == total_offset_19[6:0] ? field_byte_19 : _GEN_3753; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3850 = 7'h8 == total_offset_19[6:0] ? field_byte_19 : _GEN_3754; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3851 = 7'h9 == total_offset_19[6:0] ? field_byte_19 : _GEN_3755; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3852 = 7'ha == total_offset_19[6:0] ? field_byte_19 : _GEN_3756; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3853 = 7'hb == total_offset_19[6:0] ? field_byte_19 : _GEN_3757; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3854 = 7'hc == total_offset_19[6:0] ? field_byte_19 : _GEN_3758; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3855 = 7'hd == total_offset_19[6:0] ? field_byte_19 : _GEN_3759; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3856 = 7'he == total_offset_19[6:0] ? field_byte_19 : _GEN_3760; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3857 = 7'hf == total_offset_19[6:0] ? field_byte_19 : _GEN_3761; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3858 = 7'h10 == total_offset_19[6:0] ? field_byte_19 : _GEN_3762; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3859 = 7'h11 == total_offset_19[6:0] ? field_byte_19 : _GEN_3763; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3860 = 7'h12 == total_offset_19[6:0] ? field_byte_19 : _GEN_3764; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3861 = 7'h13 == total_offset_19[6:0] ? field_byte_19 : _GEN_3765; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3862 = 7'h14 == total_offset_19[6:0] ? field_byte_19 : _GEN_3766; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3863 = 7'h15 == total_offset_19[6:0] ? field_byte_19 : _GEN_3767; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3864 = 7'h16 == total_offset_19[6:0] ? field_byte_19 : _GEN_3768; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3865 = 7'h17 == total_offset_19[6:0] ? field_byte_19 : _GEN_3769; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3866 = 7'h18 == total_offset_19[6:0] ? field_byte_19 : _GEN_3770; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3867 = 7'h19 == total_offset_19[6:0] ? field_byte_19 : _GEN_3771; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3868 = 7'h1a == total_offset_19[6:0] ? field_byte_19 : _GEN_3772; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3869 = 7'h1b == total_offset_19[6:0] ? field_byte_19 : _GEN_3773; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3870 = 7'h1c == total_offset_19[6:0] ? field_byte_19 : _GEN_3774; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3871 = 7'h1d == total_offset_19[6:0] ? field_byte_19 : _GEN_3775; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3872 = 7'h1e == total_offset_19[6:0] ? field_byte_19 : _GEN_3776; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3873 = 7'h1f == total_offset_19[6:0] ? field_byte_19 : _GEN_3777; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3874 = 7'h20 == total_offset_19[6:0] ? field_byte_19 : _GEN_3778; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3875 = 7'h21 == total_offset_19[6:0] ? field_byte_19 : _GEN_3779; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3876 = 7'h22 == total_offset_19[6:0] ? field_byte_19 : _GEN_3780; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3877 = 7'h23 == total_offset_19[6:0] ? field_byte_19 : _GEN_3781; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3878 = 7'h24 == total_offset_19[6:0] ? field_byte_19 : _GEN_3782; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3879 = 7'h25 == total_offset_19[6:0] ? field_byte_19 : _GEN_3783; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3880 = 7'h26 == total_offset_19[6:0] ? field_byte_19 : _GEN_3784; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3881 = 7'h27 == total_offset_19[6:0] ? field_byte_19 : _GEN_3785; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3882 = 7'h28 == total_offset_19[6:0] ? field_byte_19 : _GEN_3786; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3883 = 7'h29 == total_offset_19[6:0] ? field_byte_19 : _GEN_3787; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3884 = 7'h2a == total_offset_19[6:0] ? field_byte_19 : _GEN_3788; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3885 = 7'h2b == total_offset_19[6:0] ? field_byte_19 : _GEN_3789; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3886 = 7'h2c == total_offset_19[6:0] ? field_byte_19 : _GEN_3790; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3887 = 7'h2d == total_offset_19[6:0] ? field_byte_19 : _GEN_3791; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3888 = 7'h2e == total_offset_19[6:0] ? field_byte_19 : _GEN_3792; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3889 = 7'h2f == total_offset_19[6:0] ? field_byte_19 : _GEN_3793; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3890 = 7'h30 == total_offset_19[6:0] ? field_byte_19 : _GEN_3794; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3891 = 7'h31 == total_offset_19[6:0] ? field_byte_19 : _GEN_3795; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3892 = 7'h32 == total_offset_19[6:0] ? field_byte_19 : _GEN_3796; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3893 = 7'h33 == total_offset_19[6:0] ? field_byte_19 : _GEN_3797; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3894 = 7'h34 == total_offset_19[6:0] ? field_byte_19 : _GEN_3798; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3895 = 7'h35 == total_offset_19[6:0] ? field_byte_19 : _GEN_3799; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3896 = 7'h36 == total_offset_19[6:0] ? field_byte_19 : _GEN_3800; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3897 = 7'h37 == total_offset_19[6:0] ? field_byte_19 : _GEN_3801; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3898 = 7'h38 == total_offset_19[6:0] ? field_byte_19 : _GEN_3802; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3899 = 7'h39 == total_offset_19[6:0] ? field_byte_19 : _GEN_3803; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3900 = 7'h3a == total_offset_19[6:0] ? field_byte_19 : _GEN_3804; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3901 = 7'h3b == total_offset_19[6:0] ? field_byte_19 : _GEN_3805; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3902 = 7'h3c == total_offset_19[6:0] ? field_byte_19 : _GEN_3806; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3903 = 7'h3d == total_offset_19[6:0] ? field_byte_19 : _GEN_3807; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3904 = 7'h3e == total_offset_19[6:0] ? field_byte_19 : _GEN_3808; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3905 = 7'h3f == total_offset_19[6:0] ? field_byte_19 : _GEN_3809; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3906 = 7'h40 == total_offset_19[6:0] ? field_byte_19 : _GEN_3810; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3907 = 7'h41 == total_offset_19[6:0] ? field_byte_19 : _GEN_3811; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3908 = 7'h42 == total_offset_19[6:0] ? field_byte_19 : _GEN_3812; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3909 = 7'h43 == total_offset_19[6:0] ? field_byte_19 : _GEN_3813; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3910 = 7'h44 == total_offset_19[6:0] ? field_byte_19 : _GEN_3814; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3911 = 7'h45 == total_offset_19[6:0] ? field_byte_19 : _GEN_3815; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3912 = 7'h46 == total_offset_19[6:0] ? field_byte_19 : _GEN_3816; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3913 = 7'h47 == total_offset_19[6:0] ? field_byte_19 : _GEN_3817; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3914 = 7'h48 == total_offset_19[6:0] ? field_byte_19 : _GEN_3818; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3915 = 7'h49 == total_offset_19[6:0] ? field_byte_19 : _GEN_3819; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3916 = 7'h4a == total_offset_19[6:0] ? field_byte_19 : _GEN_3820; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3917 = 7'h4b == total_offset_19[6:0] ? field_byte_19 : _GEN_3821; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3918 = 7'h4c == total_offset_19[6:0] ? field_byte_19 : _GEN_3822; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3919 = 7'h4d == total_offset_19[6:0] ? field_byte_19 : _GEN_3823; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3920 = 7'h4e == total_offset_19[6:0] ? field_byte_19 : _GEN_3824; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3921 = 7'h4f == total_offset_19[6:0] ? field_byte_19 : _GEN_3825; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3922 = 7'h50 == total_offset_19[6:0] ? field_byte_19 : _GEN_3826; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3923 = 7'h51 == total_offset_19[6:0] ? field_byte_19 : _GEN_3827; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3924 = 7'h52 == total_offset_19[6:0] ? field_byte_19 : _GEN_3828; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3925 = 7'h53 == total_offset_19[6:0] ? field_byte_19 : _GEN_3829; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3926 = 7'h54 == total_offset_19[6:0] ? field_byte_19 : _GEN_3830; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3927 = 7'h55 == total_offset_19[6:0] ? field_byte_19 : _GEN_3831; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3928 = 7'h56 == total_offset_19[6:0] ? field_byte_19 : _GEN_3832; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3929 = 7'h57 == total_offset_19[6:0] ? field_byte_19 : _GEN_3833; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3930 = 7'h58 == total_offset_19[6:0] ? field_byte_19 : _GEN_3834; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3931 = 7'h59 == total_offset_19[6:0] ? field_byte_19 : _GEN_3835; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3932 = 7'h5a == total_offset_19[6:0] ? field_byte_19 : _GEN_3836; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3933 = 7'h5b == total_offset_19[6:0] ? field_byte_19 : _GEN_3837; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3934 = 7'h5c == total_offset_19[6:0] ? field_byte_19 : _GEN_3838; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3935 = 7'h5d == total_offset_19[6:0] ? field_byte_19 : _GEN_3839; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3936 = 7'h5e == total_offset_19[6:0] ? field_byte_19 : _GEN_3840; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3937 = 7'h5f == total_offset_19[6:0] ? field_byte_19 : _GEN_3841; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_3938 = 8'h3 < length_2 ? _GEN_3842 : _GEN_3746; // @[executor.scala 290:56]
  wire [7:0] _GEN_3939 = 8'h3 < length_2 ? _GEN_3843 : _GEN_3747; // @[executor.scala 290:56]
  wire [7:0] _GEN_3940 = 8'h3 < length_2 ? _GEN_3844 : _GEN_3748; // @[executor.scala 290:56]
  wire [7:0] _GEN_3941 = 8'h3 < length_2 ? _GEN_3845 : _GEN_3749; // @[executor.scala 290:56]
  wire [7:0] _GEN_3942 = 8'h3 < length_2 ? _GEN_3846 : _GEN_3750; // @[executor.scala 290:56]
  wire [7:0] _GEN_3943 = 8'h3 < length_2 ? _GEN_3847 : _GEN_3751; // @[executor.scala 290:56]
  wire [7:0] _GEN_3944 = 8'h3 < length_2 ? _GEN_3848 : _GEN_3752; // @[executor.scala 290:56]
  wire [7:0] _GEN_3945 = 8'h3 < length_2 ? _GEN_3849 : _GEN_3753; // @[executor.scala 290:56]
  wire [7:0] _GEN_3946 = 8'h3 < length_2 ? _GEN_3850 : _GEN_3754; // @[executor.scala 290:56]
  wire [7:0] _GEN_3947 = 8'h3 < length_2 ? _GEN_3851 : _GEN_3755; // @[executor.scala 290:56]
  wire [7:0] _GEN_3948 = 8'h3 < length_2 ? _GEN_3852 : _GEN_3756; // @[executor.scala 290:56]
  wire [7:0] _GEN_3949 = 8'h3 < length_2 ? _GEN_3853 : _GEN_3757; // @[executor.scala 290:56]
  wire [7:0] _GEN_3950 = 8'h3 < length_2 ? _GEN_3854 : _GEN_3758; // @[executor.scala 290:56]
  wire [7:0] _GEN_3951 = 8'h3 < length_2 ? _GEN_3855 : _GEN_3759; // @[executor.scala 290:56]
  wire [7:0] _GEN_3952 = 8'h3 < length_2 ? _GEN_3856 : _GEN_3760; // @[executor.scala 290:56]
  wire [7:0] _GEN_3953 = 8'h3 < length_2 ? _GEN_3857 : _GEN_3761; // @[executor.scala 290:56]
  wire [7:0] _GEN_3954 = 8'h3 < length_2 ? _GEN_3858 : _GEN_3762; // @[executor.scala 290:56]
  wire [7:0] _GEN_3955 = 8'h3 < length_2 ? _GEN_3859 : _GEN_3763; // @[executor.scala 290:56]
  wire [7:0] _GEN_3956 = 8'h3 < length_2 ? _GEN_3860 : _GEN_3764; // @[executor.scala 290:56]
  wire [7:0] _GEN_3957 = 8'h3 < length_2 ? _GEN_3861 : _GEN_3765; // @[executor.scala 290:56]
  wire [7:0] _GEN_3958 = 8'h3 < length_2 ? _GEN_3862 : _GEN_3766; // @[executor.scala 290:56]
  wire [7:0] _GEN_3959 = 8'h3 < length_2 ? _GEN_3863 : _GEN_3767; // @[executor.scala 290:56]
  wire [7:0] _GEN_3960 = 8'h3 < length_2 ? _GEN_3864 : _GEN_3768; // @[executor.scala 290:56]
  wire [7:0] _GEN_3961 = 8'h3 < length_2 ? _GEN_3865 : _GEN_3769; // @[executor.scala 290:56]
  wire [7:0] _GEN_3962 = 8'h3 < length_2 ? _GEN_3866 : _GEN_3770; // @[executor.scala 290:56]
  wire [7:0] _GEN_3963 = 8'h3 < length_2 ? _GEN_3867 : _GEN_3771; // @[executor.scala 290:56]
  wire [7:0] _GEN_3964 = 8'h3 < length_2 ? _GEN_3868 : _GEN_3772; // @[executor.scala 290:56]
  wire [7:0] _GEN_3965 = 8'h3 < length_2 ? _GEN_3869 : _GEN_3773; // @[executor.scala 290:56]
  wire [7:0] _GEN_3966 = 8'h3 < length_2 ? _GEN_3870 : _GEN_3774; // @[executor.scala 290:56]
  wire [7:0] _GEN_3967 = 8'h3 < length_2 ? _GEN_3871 : _GEN_3775; // @[executor.scala 290:56]
  wire [7:0] _GEN_3968 = 8'h3 < length_2 ? _GEN_3872 : _GEN_3776; // @[executor.scala 290:56]
  wire [7:0] _GEN_3969 = 8'h3 < length_2 ? _GEN_3873 : _GEN_3777; // @[executor.scala 290:56]
  wire [7:0] _GEN_3970 = 8'h3 < length_2 ? _GEN_3874 : _GEN_3778; // @[executor.scala 290:56]
  wire [7:0] _GEN_3971 = 8'h3 < length_2 ? _GEN_3875 : _GEN_3779; // @[executor.scala 290:56]
  wire [7:0] _GEN_3972 = 8'h3 < length_2 ? _GEN_3876 : _GEN_3780; // @[executor.scala 290:56]
  wire [7:0] _GEN_3973 = 8'h3 < length_2 ? _GEN_3877 : _GEN_3781; // @[executor.scala 290:56]
  wire [7:0] _GEN_3974 = 8'h3 < length_2 ? _GEN_3878 : _GEN_3782; // @[executor.scala 290:56]
  wire [7:0] _GEN_3975 = 8'h3 < length_2 ? _GEN_3879 : _GEN_3783; // @[executor.scala 290:56]
  wire [7:0] _GEN_3976 = 8'h3 < length_2 ? _GEN_3880 : _GEN_3784; // @[executor.scala 290:56]
  wire [7:0] _GEN_3977 = 8'h3 < length_2 ? _GEN_3881 : _GEN_3785; // @[executor.scala 290:56]
  wire [7:0] _GEN_3978 = 8'h3 < length_2 ? _GEN_3882 : _GEN_3786; // @[executor.scala 290:56]
  wire [7:0] _GEN_3979 = 8'h3 < length_2 ? _GEN_3883 : _GEN_3787; // @[executor.scala 290:56]
  wire [7:0] _GEN_3980 = 8'h3 < length_2 ? _GEN_3884 : _GEN_3788; // @[executor.scala 290:56]
  wire [7:0] _GEN_3981 = 8'h3 < length_2 ? _GEN_3885 : _GEN_3789; // @[executor.scala 290:56]
  wire [7:0] _GEN_3982 = 8'h3 < length_2 ? _GEN_3886 : _GEN_3790; // @[executor.scala 290:56]
  wire [7:0] _GEN_3983 = 8'h3 < length_2 ? _GEN_3887 : _GEN_3791; // @[executor.scala 290:56]
  wire [7:0] _GEN_3984 = 8'h3 < length_2 ? _GEN_3888 : _GEN_3792; // @[executor.scala 290:56]
  wire [7:0] _GEN_3985 = 8'h3 < length_2 ? _GEN_3889 : _GEN_3793; // @[executor.scala 290:56]
  wire [7:0] _GEN_3986 = 8'h3 < length_2 ? _GEN_3890 : _GEN_3794; // @[executor.scala 290:56]
  wire [7:0] _GEN_3987 = 8'h3 < length_2 ? _GEN_3891 : _GEN_3795; // @[executor.scala 290:56]
  wire [7:0] _GEN_3988 = 8'h3 < length_2 ? _GEN_3892 : _GEN_3796; // @[executor.scala 290:56]
  wire [7:0] _GEN_3989 = 8'h3 < length_2 ? _GEN_3893 : _GEN_3797; // @[executor.scala 290:56]
  wire [7:0] _GEN_3990 = 8'h3 < length_2 ? _GEN_3894 : _GEN_3798; // @[executor.scala 290:56]
  wire [7:0] _GEN_3991 = 8'h3 < length_2 ? _GEN_3895 : _GEN_3799; // @[executor.scala 290:56]
  wire [7:0] _GEN_3992 = 8'h3 < length_2 ? _GEN_3896 : _GEN_3800; // @[executor.scala 290:56]
  wire [7:0] _GEN_3993 = 8'h3 < length_2 ? _GEN_3897 : _GEN_3801; // @[executor.scala 290:56]
  wire [7:0] _GEN_3994 = 8'h3 < length_2 ? _GEN_3898 : _GEN_3802; // @[executor.scala 290:56]
  wire [7:0] _GEN_3995 = 8'h3 < length_2 ? _GEN_3899 : _GEN_3803; // @[executor.scala 290:56]
  wire [7:0] _GEN_3996 = 8'h3 < length_2 ? _GEN_3900 : _GEN_3804; // @[executor.scala 290:56]
  wire [7:0] _GEN_3997 = 8'h3 < length_2 ? _GEN_3901 : _GEN_3805; // @[executor.scala 290:56]
  wire [7:0] _GEN_3998 = 8'h3 < length_2 ? _GEN_3902 : _GEN_3806; // @[executor.scala 290:56]
  wire [7:0] _GEN_3999 = 8'h3 < length_2 ? _GEN_3903 : _GEN_3807; // @[executor.scala 290:56]
  wire [7:0] _GEN_4000 = 8'h3 < length_2 ? _GEN_3904 : _GEN_3808; // @[executor.scala 290:56]
  wire [7:0] _GEN_4001 = 8'h3 < length_2 ? _GEN_3905 : _GEN_3809; // @[executor.scala 290:56]
  wire [7:0] _GEN_4002 = 8'h3 < length_2 ? _GEN_3906 : _GEN_3810; // @[executor.scala 290:56]
  wire [7:0] _GEN_4003 = 8'h3 < length_2 ? _GEN_3907 : _GEN_3811; // @[executor.scala 290:56]
  wire [7:0] _GEN_4004 = 8'h3 < length_2 ? _GEN_3908 : _GEN_3812; // @[executor.scala 290:56]
  wire [7:0] _GEN_4005 = 8'h3 < length_2 ? _GEN_3909 : _GEN_3813; // @[executor.scala 290:56]
  wire [7:0] _GEN_4006 = 8'h3 < length_2 ? _GEN_3910 : _GEN_3814; // @[executor.scala 290:56]
  wire [7:0] _GEN_4007 = 8'h3 < length_2 ? _GEN_3911 : _GEN_3815; // @[executor.scala 290:56]
  wire [7:0] _GEN_4008 = 8'h3 < length_2 ? _GEN_3912 : _GEN_3816; // @[executor.scala 290:56]
  wire [7:0] _GEN_4009 = 8'h3 < length_2 ? _GEN_3913 : _GEN_3817; // @[executor.scala 290:56]
  wire [7:0] _GEN_4010 = 8'h3 < length_2 ? _GEN_3914 : _GEN_3818; // @[executor.scala 290:56]
  wire [7:0] _GEN_4011 = 8'h3 < length_2 ? _GEN_3915 : _GEN_3819; // @[executor.scala 290:56]
  wire [7:0] _GEN_4012 = 8'h3 < length_2 ? _GEN_3916 : _GEN_3820; // @[executor.scala 290:56]
  wire [7:0] _GEN_4013 = 8'h3 < length_2 ? _GEN_3917 : _GEN_3821; // @[executor.scala 290:56]
  wire [7:0] _GEN_4014 = 8'h3 < length_2 ? _GEN_3918 : _GEN_3822; // @[executor.scala 290:56]
  wire [7:0] _GEN_4015 = 8'h3 < length_2 ? _GEN_3919 : _GEN_3823; // @[executor.scala 290:56]
  wire [7:0] _GEN_4016 = 8'h3 < length_2 ? _GEN_3920 : _GEN_3824; // @[executor.scala 290:56]
  wire [7:0] _GEN_4017 = 8'h3 < length_2 ? _GEN_3921 : _GEN_3825; // @[executor.scala 290:56]
  wire [7:0] _GEN_4018 = 8'h3 < length_2 ? _GEN_3922 : _GEN_3826; // @[executor.scala 290:56]
  wire [7:0] _GEN_4019 = 8'h3 < length_2 ? _GEN_3923 : _GEN_3827; // @[executor.scala 290:56]
  wire [7:0] _GEN_4020 = 8'h3 < length_2 ? _GEN_3924 : _GEN_3828; // @[executor.scala 290:56]
  wire [7:0] _GEN_4021 = 8'h3 < length_2 ? _GEN_3925 : _GEN_3829; // @[executor.scala 290:56]
  wire [7:0] _GEN_4022 = 8'h3 < length_2 ? _GEN_3926 : _GEN_3830; // @[executor.scala 290:56]
  wire [7:0] _GEN_4023 = 8'h3 < length_2 ? _GEN_3927 : _GEN_3831; // @[executor.scala 290:56]
  wire [7:0] _GEN_4024 = 8'h3 < length_2 ? _GEN_3928 : _GEN_3832; // @[executor.scala 290:56]
  wire [7:0] _GEN_4025 = 8'h3 < length_2 ? _GEN_3929 : _GEN_3833; // @[executor.scala 290:56]
  wire [7:0] _GEN_4026 = 8'h3 < length_2 ? _GEN_3930 : _GEN_3834; // @[executor.scala 290:56]
  wire [7:0] _GEN_4027 = 8'h3 < length_2 ? _GEN_3931 : _GEN_3835; // @[executor.scala 290:56]
  wire [7:0] _GEN_4028 = 8'h3 < length_2 ? _GEN_3932 : _GEN_3836; // @[executor.scala 290:56]
  wire [7:0] _GEN_4029 = 8'h3 < length_2 ? _GEN_3933 : _GEN_3837; // @[executor.scala 290:56]
  wire [7:0] _GEN_4030 = 8'h3 < length_2 ? _GEN_3934 : _GEN_3838; // @[executor.scala 290:56]
  wire [7:0] _GEN_4031 = 8'h3 < length_2 ? _GEN_3935 : _GEN_3839; // @[executor.scala 290:56]
  wire [7:0] _GEN_4032 = 8'h3 < length_2 ? _GEN_3936 : _GEN_3840; // @[executor.scala 290:56]
  wire [7:0] _GEN_4033 = 8'h3 < length_2 ? _GEN_3937 : _GEN_3841; // @[executor.scala 290:56]
  wire [7:0] field_byte_20 = field_2[31:24]; // @[executor.scala 287:53]
  wire [7:0] total_offset_20 = offset_2 + 8'h4; // @[executor.scala 289:53]
  wire [7:0] _GEN_4034 = 7'h0 == total_offset_20[6:0] ? field_byte_20 : _GEN_3938; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4035 = 7'h1 == total_offset_20[6:0] ? field_byte_20 : _GEN_3939; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4036 = 7'h2 == total_offset_20[6:0] ? field_byte_20 : _GEN_3940; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4037 = 7'h3 == total_offset_20[6:0] ? field_byte_20 : _GEN_3941; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4038 = 7'h4 == total_offset_20[6:0] ? field_byte_20 : _GEN_3942; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4039 = 7'h5 == total_offset_20[6:0] ? field_byte_20 : _GEN_3943; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4040 = 7'h6 == total_offset_20[6:0] ? field_byte_20 : _GEN_3944; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4041 = 7'h7 == total_offset_20[6:0] ? field_byte_20 : _GEN_3945; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4042 = 7'h8 == total_offset_20[6:0] ? field_byte_20 : _GEN_3946; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4043 = 7'h9 == total_offset_20[6:0] ? field_byte_20 : _GEN_3947; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4044 = 7'ha == total_offset_20[6:0] ? field_byte_20 : _GEN_3948; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4045 = 7'hb == total_offset_20[6:0] ? field_byte_20 : _GEN_3949; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4046 = 7'hc == total_offset_20[6:0] ? field_byte_20 : _GEN_3950; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4047 = 7'hd == total_offset_20[6:0] ? field_byte_20 : _GEN_3951; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4048 = 7'he == total_offset_20[6:0] ? field_byte_20 : _GEN_3952; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4049 = 7'hf == total_offset_20[6:0] ? field_byte_20 : _GEN_3953; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4050 = 7'h10 == total_offset_20[6:0] ? field_byte_20 : _GEN_3954; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4051 = 7'h11 == total_offset_20[6:0] ? field_byte_20 : _GEN_3955; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4052 = 7'h12 == total_offset_20[6:0] ? field_byte_20 : _GEN_3956; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4053 = 7'h13 == total_offset_20[6:0] ? field_byte_20 : _GEN_3957; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4054 = 7'h14 == total_offset_20[6:0] ? field_byte_20 : _GEN_3958; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4055 = 7'h15 == total_offset_20[6:0] ? field_byte_20 : _GEN_3959; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4056 = 7'h16 == total_offset_20[6:0] ? field_byte_20 : _GEN_3960; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4057 = 7'h17 == total_offset_20[6:0] ? field_byte_20 : _GEN_3961; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4058 = 7'h18 == total_offset_20[6:0] ? field_byte_20 : _GEN_3962; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4059 = 7'h19 == total_offset_20[6:0] ? field_byte_20 : _GEN_3963; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4060 = 7'h1a == total_offset_20[6:0] ? field_byte_20 : _GEN_3964; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4061 = 7'h1b == total_offset_20[6:0] ? field_byte_20 : _GEN_3965; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4062 = 7'h1c == total_offset_20[6:0] ? field_byte_20 : _GEN_3966; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4063 = 7'h1d == total_offset_20[6:0] ? field_byte_20 : _GEN_3967; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4064 = 7'h1e == total_offset_20[6:0] ? field_byte_20 : _GEN_3968; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4065 = 7'h1f == total_offset_20[6:0] ? field_byte_20 : _GEN_3969; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4066 = 7'h20 == total_offset_20[6:0] ? field_byte_20 : _GEN_3970; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4067 = 7'h21 == total_offset_20[6:0] ? field_byte_20 : _GEN_3971; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4068 = 7'h22 == total_offset_20[6:0] ? field_byte_20 : _GEN_3972; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4069 = 7'h23 == total_offset_20[6:0] ? field_byte_20 : _GEN_3973; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4070 = 7'h24 == total_offset_20[6:0] ? field_byte_20 : _GEN_3974; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4071 = 7'h25 == total_offset_20[6:0] ? field_byte_20 : _GEN_3975; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4072 = 7'h26 == total_offset_20[6:0] ? field_byte_20 : _GEN_3976; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4073 = 7'h27 == total_offset_20[6:0] ? field_byte_20 : _GEN_3977; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4074 = 7'h28 == total_offset_20[6:0] ? field_byte_20 : _GEN_3978; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4075 = 7'h29 == total_offset_20[6:0] ? field_byte_20 : _GEN_3979; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4076 = 7'h2a == total_offset_20[6:0] ? field_byte_20 : _GEN_3980; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4077 = 7'h2b == total_offset_20[6:0] ? field_byte_20 : _GEN_3981; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4078 = 7'h2c == total_offset_20[6:0] ? field_byte_20 : _GEN_3982; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4079 = 7'h2d == total_offset_20[6:0] ? field_byte_20 : _GEN_3983; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4080 = 7'h2e == total_offset_20[6:0] ? field_byte_20 : _GEN_3984; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4081 = 7'h2f == total_offset_20[6:0] ? field_byte_20 : _GEN_3985; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4082 = 7'h30 == total_offset_20[6:0] ? field_byte_20 : _GEN_3986; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4083 = 7'h31 == total_offset_20[6:0] ? field_byte_20 : _GEN_3987; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4084 = 7'h32 == total_offset_20[6:0] ? field_byte_20 : _GEN_3988; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4085 = 7'h33 == total_offset_20[6:0] ? field_byte_20 : _GEN_3989; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4086 = 7'h34 == total_offset_20[6:0] ? field_byte_20 : _GEN_3990; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4087 = 7'h35 == total_offset_20[6:0] ? field_byte_20 : _GEN_3991; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4088 = 7'h36 == total_offset_20[6:0] ? field_byte_20 : _GEN_3992; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4089 = 7'h37 == total_offset_20[6:0] ? field_byte_20 : _GEN_3993; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4090 = 7'h38 == total_offset_20[6:0] ? field_byte_20 : _GEN_3994; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4091 = 7'h39 == total_offset_20[6:0] ? field_byte_20 : _GEN_3995; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4092 = 7'h3a == total_offset_20[6:0] ? field_byte_20 : _GEN_3996; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4093 = 7'h3b == total_offset_20[6:0] ? field_byte_20 : _GEN_3997; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4094 = 7'h3c == total_offset_20[6:0] ? field_byte_20 : _GEN_3998; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4095 = 7'h3d == total_offset_20[6:0] ? field_byte_20 : _GEN_3999; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4096 = 7'h3e == total_offset_20[6:0] ? field_byte_20 : _GEN_4000; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4097 = 7'h3f == total_offset_20[6:0] ? field_byte_20 : _GEN_4001; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4098 = 7'h40 == total_offset_20[6:0] ? field_byte_20 : _GEN_4002; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4099 = 7'h41 == total_offset_20[6:0] ? field_byte_20 : _GEN_4003; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4100 = 7'h42 == total_offset_20[6:0] ? field_byte_20 : _GEN_4004; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4101 = 7'h43 == total_offset_20[6:0] ? field_byte_20 : _GEN_4005; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4102 = 7'h44 == total_offset_20[6:0] ? field_byte_20 : _GEN_4006; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4103 = 7'h45 == total_offset_20[6:0] ? field_byte_20 : _GEN_4007; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4104 = 7'h46 == total_offset_20[6:0] ? field_byte_20 : _GEN_4008; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4105 = 7'h47 == total_offset_20[6:0] ? field_byte_20 : _GEN_4009; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4106 = 7'h48 == total_offset_20[6:0] ? field_byte_20 : _GEN_4010; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4107 = 7'h49 == total_offset_20[6:0] ? field_byte_20 : _GEN_4011; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4108 = 7'h4a == total_offset_20[6:0] ? field_byte_20 : _GEN_4012; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4109 = 7'h4b == total_offset_20[6:0] ? field_byte_20 : _GEN_4013; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4110 = 7'h4c == total_offset_20[6:0] ? field_byte_20 : _GEN_4014; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4111 = 7'h4d == total_offset_20[6:0] ? field_byte_20 : _GEN_4015; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4112 = 7'h4e == total_offset_20[6:0] ? field_byte_20 : _GEN_4016; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4113 = 7'h4f == total_offset_20[6:0] ? field_byte_20 : _GEN_4017; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4114 = 7'h50 == total_offset_20[6:0] ? field_byte_20 : _GEN_4018; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4115 = 7'h51 == total_offset_20[6:0] ? field_byte_20 : _GEN_4019; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4116 = 7'h52 == total_offset_20[6:0] ? field_byte_20 : _GEN_4020; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4117 = 7'h53 == total_offset_20[6:0] ? field_byte_20 : _GEN_4021; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4118 = 7'h54 == total_offset_20[6:0] ? field_byte_20 : _GEN_4022; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4119 = 7'h55 == total_offset_20[6:0] ? field_byte_20 : _GEN_4023; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4120 = 7'h56 == total_offset_20[6:0] ? field_byte_20 : _GEN_4024; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4121 = 7'h57 == total_offset_20[6:0] ? field_byte_20 : _GEN_4025; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4122 = 7'h58 == total_offset_20[6:0] ? field_byte_20 : _GEN_4026; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4123 = 7'h59 == total_offset_20[6:0] ? field_byte_20 : _GEN_4027; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4124 = 7'h5a == total_offset_20[6:0] ? field_byte_20 : _GEN_4028; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4125 = 7'h5b == total_offset_20[6:0] ? field_byte_20 : _GEN_4029; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4126 = 7'h5c == total_offset_20[6:0] ? field_byte_20 : _GEN_4030; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4127 = 7'h5d == total_offset_20[6:0] ? field_byte_20 : _GEN_4031; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4128 = 7'h5e == total_offset_20[6:0] ? field_byte_20 : _GEN_4032; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4129 = 7'h5f == total_offset_20[6:0] ? field_byte_20 : _GEN_4033; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4130 = 8'h4 < length_2 ? _GEN_4034 : _GEN_3938; // @[executor.scala 290:56]
  wire [7:0] _GEN_4131 = 8'h4 < length_2 ? _GEN_4035 : _GEN_3939; // @[executor.scala 290:56]
  wire [7:0] _GEN_4132 = 8'h4 < length_2 ? _GEN_4036 : _GEN_3940; // @[executor.scala 290:56]
  wire [7:0] _GEN_4133 = 8'h4 < length_2 ? _GEN_4037 : _GEN_3941; // @[executor.scala 290:56]
  wire [7:0] _GEN_4134 = 8'h4 < length_2 ? _GEN_4038 : _GEN_3942; // @[executor.scala 290:56]
  wire [7:0] _GEN_4135 = 8'h4 < length_2 ? _GEN_4039 : _GEN_3943; // @[executor.scala 290:56]
  wire [7:0] _GEN_4136 = 8'h4 < length_2 ? _GEN_4040 : _GEN_3944; // @[executor.scala 290:56]
  wire [7:0] _GEN_4137 = 8'h4 < length_2 ? _GEN_4041 : _GEN_3945; // @[executor.scala 290:56]
  wire [7:0] _GEN_4138 = 8'h4 < length_2 ? _GEN_4042 : _GEN_3946; // @[executor.scala 290:56]
  wire [7:0] _GEN_4139 = 8'h4 < length_2 ? _GEN_4043 : _GEN_3947; // @[executor.scala 290:56]
  wire [7:0] _GEN_4140 = 8'h4 < length_2 ? _GEN_4044 : _GEN_3948; // @[executor.scala 290:56]
  wire [7:0] _GEN_4141 = 8'h4 < length_2 ? _GEN_4045 : _GEN_3949; // @[executor.scala 290:56]
  wire [7:0] _GEN_4142 = 8'h4 < length_2 ? _GEN_4046 : _GEN_3950; // @[executor.scala 290:56]
  wire [7:0] _GEN_4143 = 8'h4 < length_2 ? _GEN_4047 : _GEN_3951; // @[executor.scala 290:56]
  wire [7:0] _GEN_4144 = 8'h4 < length_2 ? _GEN_4048 : _GEN_3952; // @[executor.scala 290:56]
  wire [7:0] _GEN_4145 = 8'h4 < length_2 ? _GEN_4049 : _GEN_3953; // @[executor.scala 290:56]
  wire [7:0] _GEN_4146 = 8'h4 < length_2 ? _GEN_4050 : _GEN_3954; // @[executor.scala 290:56]
  wire [7:0] _GEN_4147 = 8'h4 < length_2 ? _GEN_4051 : _GEN_3955; // @[executor.scala 290:56]
  wire [7:0] _GEN_4148 = 8'h4 < length_2 ? _GEN_4052 : _GEN_3956; // @[executor.scala 290:56]
  wire [7:0] _GEN_4149 = 8'h4 < length_2 ? _GEN_4053 : _GEN_3957; // @[executor.scala 290:56]
  wire [7:0] _GEN_4150 = 8'h4 < length_2 ? _GEN_4054 : _GEN_3958; // @[executor.scala 290:56]
  wire [7:0] _GEN_4151 = 8'h4 < length_2 ? _GEN_4055 : _GEN_3959; // @[executor.scala 290:56]
  wire [7:0] _GEN_4152 = 8'h4 < length_2 ? _GEN_4056 : _GEN_3960; // @[executor.scala 290:56]
  wire [7:0] _GEN_4153 = 8'h4 < length_2 ? _GEN_4057 : _GEN_3961; // @[executor.scala 290:56]
  wire [7:0] _GEN_4154 = 8'h4 < length_2 ? _GEN_4058 : _GEN_3962; // @[executor.scala 290:56]
  wire [7:0] _GEN_4155 = 8'h4 < length_2 ? _GEN_4059 : _GEN_3963; // @[executor.scala 290:56]
  wire [7:0] _GEN_4156 = 8'h4 < length_2 ? _GEN_4060 : _GEN_3964; // @[executor.scala 290:56]
  wire [7:0] _GEN_4157 = 8'h4 < length_2 ? _GEN_4061 : _GEN_3965; // @[executor.scala 290:56]
  wire [7:0] _GEN_4158 = 8'h4 < length_2 ? _GEN_4062 : _GEN_3966; // @[executor.scala 290:56]
  wire [7:0] _GEN_4159 = 8'h4 < length_2 ? _GEN_4063 : _GEN_3967; // @[executor.scala 290:56]
  wire [7:0] _GEN_4160 = 8'h4 < length_2 ? _GEN_4064 : _GEN_3968; // @[executor.scala 290:56]
  wire [7:0] _GEN_4161 = 8'h4 < length_2 ? _GEN_4065 : _GEN_3969; // @[executor.scala 290:56]
  wire [7:0] _GEN_4162 = 8'h4 < length_2 ? _GEN_4066 : _GEN_3970; // @[executor.scala 290:56]
  wire [7:0] _GEN_4163 = 8'h4 < length_2 ? _GEN_4067 : _GEN_3971; // @[executor.scala 290:56]
  wire [7:0] _GEN_4164 = 8'h4 < length_2 ? _GEN_4068 : _GEN_3972; // @[executor.scala 290:56]
  wire [7:0] _GEN_4165 = 8'h4 < length_2 ? _GEN_4069 : _GEN_3973; // @[executor.scala 290:56]
  wire [7:0] _GEN_4166 = 8'h4 < length_2 ? _GEN_4070 : _GEN_3974; // @[executor.scala 290:56]
  wire [7:0] _GEN_4167 = 8'h4 < length_2 ? _GEN_4071 : _GEN_3975; // @[executor.scala 290:56]
  wire [7:0] _GEN_4168 = 8'h4 < length_2 ? _GEN_4072 : _GEN_3976; // @[executor.scala 290:56]
  wire [7:0] _GEN_4169 = 8'h4 < length_2 ? _GEN_4073 : _GEN_3977; // @[executor.scala 290:56]
  wire [7:0] _GEN_4170 = 8'h4 < length_2 ? _GEN_4074 : _GEN_3978; // @[executor.scala 290:56]
  wire [7:0] _GEN_4171 = 8'h4 < length_2 ? _GEN_4075 : _GEN_3979; // @[executor.scala 290:56]
  wire [7:0] _GEN_4172 = 8'h4 < length_2 ? _GEN_4076 : _GEN_3980; // @[executor.scala 290:56]
  wire [7:0] _GEN_4173 = 8'h4 < length_2 ? _GEN_4077 : _GEN_3981; // @[executor.scala 290:56]
  wire [7:0] _GEN_4174 = 8'h4 < length_2 ? _GEN_4078 : _GEN_3982; // @[executor.scala 290:56]
  wire [7:0] _GEN_4175 = 8'h4 < length_2 ? _GEN_4079 : _GEN_3983; // @[executor.scala 290:56]
  wire [7:0] _GEN_4176 = 8'h4 < length_2 ? _GEN_4080 : _GEN_3984; // @[executor.scala 290:56]
  wire [7:0] _GEN_4177 = 8'h4 < length_2 ? _GEN_4081 : _GEN_3985; // @[executor.scala 290:56]
  wire [7:0] _GEN_4178 = 8'h4 < length_2 ? _GEN_4082 : _GEN_3986; // @[executor.scala 290:56]
  wire [7:0] _GEN_4179 = 8'h4 < length_2 ? _GEN_4083 : _GEN_3987; // @[executor.scala 290:56]
  wire [7:0] _GEN_4180 = 8'h4 < length_2 ? _GEN_4084 : _GEN_3988; // @[executor.scala 290:56]
  wire [7:0] _GEN_4181 = 8'h4 < length_2 ? _GEN_4085 : _GEN_3989; // @[executor.scala 290:56]
  wire [7:0] _GEN_4182 = 8'h4 < length_2 ? _GEN_4086 : _GEN_3990; // @[executor.scala 290:56]
  wire [7:0] _GEN_4183 = 8'h4 < length_2 ? _GEN_4087 : _GEN_3991; // @[executor.scala 290:56]
  wire [7:0] _GEN_4184 = 8'h4 < length_2 ? _GEN_4088 : _GEN_3992; // @[executor.scala 290:56]
  wire [7:0] _GEN_4185 = 8'h4 < length_2 ? _GEN_4089 : _GEN_3993; // @[executor.scala 290:56]
  wire [7:0] _GEN_4186 = 8'h4 < length_2 ? _GEN_4090 : _GEN_3994; // @[executor.scala 290:56]
  wire [7:0] _GEN_4187 = 8'h4 < length_2 ? _GEN_4091 : _GEN_3995; // @[executor.scala 290:56]
  wire [7:0] _GEN_4188 = 8'h4 < length_2 ? _GEN_4092 : _GEN_3996; // @[executor.scala 290:56]
  wire [7:0] _GEN_4189 = 8'h4 < length_2 ? _GEN_4093 : _GEN_3997; // @[executor.scala 290:56]
  wire [7:0] _GEN_4190 = 8'h4 < length_2 ? _GEN_4094 : _GEN_3998; // @[executor.scala 290:56]
  wire [7:0] _GEN_4191 = 8'h4 < length_2 ? _GEN_4095 : _GEN_3999; // @[executor.scala 290:56]
  wire [7:0] _GEN_4192 = 8'h4 < length_2 ? _GEN_4096 : _GEN_4000; // @[executor.scala 290:56]
  wire [7:0] _GEN_4193 = 8'h4 < length_2 ? _GEN_4097 : _GEN_4001; // @[executor.scala 290:56]
  wire [7:0] _GEN_4194 = 8'h4 < length_2 ? _GEN_4098 : _GEN_4002; // @[executor.scala 290:56]
  wire [7:0] _GEN_4195 = 8'h4 < length_2 ? _GEN_4099 : _GEN_4003; // @[executor.scala 290:56]
  wire [7:0] _GEN_4196 = 8'h4 < length_2 ? _GEN_4100 : _GEN_4004; // @[executor.scala 290:56]
  wire [7:0] _GEN_4197 = 8'h4 < length_2 ? _GEN_4101 : _GEN_4005; // @[executor.scala 290:56]
  wire [7:0] _GEN_4198 = 8'h4 < length_2 ? _GEN_4102 : _GEN_4006; // @[executor.scala 290:56]
  wire [7:0] _GEN_4199 = 8'h4 < length_2 ? _GEN_4103 : _GEN_4007; // @[executor.scala 290:56]
  wire [7:0] _GEN_4200 = 8'h4 < length_2 ? _GEN_4104 : _GEN_4008; // @[executor.scala 290:56]
  wire [7:0] _GEN_4201 = 8'h4 < length_2 ? _GEN_4105 : _GEN_4009; // @[executor.scala 290:56]
  wire [7:0] _GEN_4202 = 8'h4 < length_2 ? _GEN_4106 : _GEN_4010; // @[executor.scala 290:56]
  wire [7:0] _GEN_4203 = 8'h4 < length_2 ? _GEN_4107 : _GEN_4011; // @[executor.scala 290:56]
  wire [7:0] _GEN_4204 = 8'h4 < length_2 ? _GEN_4108 : _GEN_4012; // @[executor.scala 290:56]
  wire [7:0] _GEN_4205 = 8'h4 < length_2 ? _GEN_4109 : _GEN_4013; // @[executor.scala 290:56]
  wire [7:0] _GEN_4206 = 8'h4 < length_2 ? _GEN_4110 : _GEN_4014; // @[executor.scala 290:56]
  wire [7:0] _GEN_4207 = 8'h4 < length_2 ? _GEN_4111 : _GEN_4015; // @[executor.scala 290:56]
  wire [7:0] _GEN_4208 = 8'h4 < length_2 ? _GEN_4112 : _GEN_4016; // @[executor.scala 290:56]
  wire [7:0] _GEN_4209 = 8'h4 < length_2 ? _GEN_4113 : _GEN_4017; // @[executor.scala 290:56]
  wire [7:0] _GEN_4210 = 8'h4 < length_2 ? _GEN_4114 : _GEN_4018; // @[executor.scala 290:56]
  wire [7:0] _GEN_4211 = 8'h4 < length_2 ? _GEN_4115 : _GEN_4019; // @[executor.scala 290:56]
  wire [7:0] _GEN_4212 = 8'h4 < length_2 ? _GEN_4116 : _GEN_4020; // @[executor.scala 290:56]
  wire [7:0] _GEN_4213 = 8'h4 < length_2 ? _GEN_4117 : _GEN_4021; // @[executor.scala 290:56]
  wire [7:0] _GEN_4214 = 8'h4 < length_2 ? _GEN_4118 : _GEN_4022; // @[executor.scala 290:56]
  wire [7:0] _GEN_4215 = 8'h4 < length_2 ? _GEN_4119 : _GEN_4023; // @[executor.scala 290:56]
  wire [7:0] _GEN_4216 = 8'h4 < length_2 ? _GEN_4120 : _GEN_4024; // @[executor.scala 290:56]
  wire [7:0] _GEN_4217 = 8'h4 < length_2 ? _GEN_4121 : _GEN_4025; // @[executor.scala 290:56]
  wire [7:0] _GEN_4218 = 8'h4 < length_2 ? _GEN_4122 : _GEN_4026; // @[executor.scala 290:56]
  wire [7:0] _GEN_4219 = 8'h4 < length_2 ? _GEN_4123 : _GEN_4027; // @[executor.scala 290:56]
  wire [7:0] _GEN_4220 = 8'h4 < length_2 ? _GEN_4124 : _GEN_4028; // @[executor.scala 290:56]
  wire [7:0] _GEN_4221 = 8'h4 < length_2 ? _GEN_4125 : _GEN_4029; // @[executor.scala 290:56]
  wire [7:0] _GEN_4222 = 8'h4 < length_2 ? _GEN_4126 : _GEN_4030; // @[executor.scala 290:56]
  wire [7:0] _GEN_4223 = 8'h4 < length_2 ? _GEN_4127 : _GEN_4031; // @[executor.scala 290:56]
  wire [7:0] _GEN_4224 = 8'h4 < length_2 ? _GEN_4128 : _GEN_4032; // @[executor.scala 290:56]
  wire [7:0] _GEN_4225 = 8'h4 < length_2 ? _GEN_4129 : _GEN_4033; // @[executor.scala 290:56]
  wire [7:0] field_byte_21 = field_2[23:16]; // @[executor.scala 287:53]
  wire [7:0] total_offset_21 = offset_2 + 8'h5; // @[executor.scala 289:53]
  wire [7:0] _GEN_4226 = 7'h0 == total_offset_21[6:0] ? field_byte_21 : _GEN_4130; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4227 = 7'h1 == total_offset_21[6:0] ? field_byte_21 : _GEN_4131; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4228 = 7'h2 == total_offset_21[6:0] ? field_byte_21 : _GEN_4132; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4229 = 7'h3 == total_offset_21[6:0] ? field_byte_21 : _GEN_4133; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4230 = 7'h4 == total_offset_21[6:0] ? field_byte_21 : _GEN_4134; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4231 = 7'h5 == total_offset_21[6:0] ? field_byte_21 : _GEN_4135; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4232 = 7'h6 == total_offset_21[6:0] ? field_byte_21 : _GEN_4136; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4233 = 7'h7 == total_offset_21[6:0] ? field_byte_21 : _GEN_4137; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4234 = 7'h8 == total_offset_21[6:0] ? field_byte_21 : _GEN_4138; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4235 = 7'h9 == total_offset_21[6:0] ? field_byte_21 : _GEN_4139; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4236 = 7'ha == total_offset_21[6:0] ? field_byte_21 : _GEN_4140; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4237 = 7'hb == total_offset_21[6:0] ? field_byte_21 : _GEN_4141; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4238 = 7'hc == total_offset_21[6:0] ? field_byte_21 : _GEN_4142; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4239 = 7'hd == total_offset_21[6:0] ? field_byte_21 : _GEN_4143; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4240 = 7'he == total_offset_21[6:0] ? field_byte_21 : _GEN_4144; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4241 = 7'hf == total_offset_21[6:0] ? field_byte_21 : _GEN_4145; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4242 = 7'h10 == total_offset_21[6:0] ? field_byte_21 : _GEN_4146; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4243 = 7'h11 == total_offset_21[6:0] ? field_byte_21 : _GEN_4147; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4244 = 7'h12 == total_offset_21[6:0] ? field_byte_21 : _GEN_4148; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4245 = 7'h13 == total_offset_21[6:0] ? field_byte_21 : _GEN_4149; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4246 = 7'h14 == total_offset_21[6:0] ? field_byte_21 : _GEN_4150; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4247 = 7'h15 == total_offset_21[6:0] ? field_byte_21 : _GEN_4151; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4248 = 7'h16 == total_offset_21[6:0] ? field_byte_21 : _GEN_4152; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4249 = 7'h17 == total_offset_21[6:0] ? field_byte_21 : _GEN_4153; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4250 = 7'h18 == total_offset_21[6:0] ? field_byte_21 : _GEN_4154; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4251 = 7'h19 == total_offset_21[6:0] ? field_byte_21 : _GEN_4155; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4252 = 7'h1a == total_offset_21[6:0] ? field_byte_21 : _GEN_4156; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4253 = 7'h1b == total_offset_21[6:0] ? field_byte_21 : _GEN_4157; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4254 = 7'h1c == total_offset_21[6:0] ? field_byte_21 : _GEN_4158; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4255 = 7'h1d == total_offset_21[6:0] ? field_byte_21 : _GEN_4159; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4256 = 7'h1e == total_offset_21[6:0] ? field_byte_21 : _GEN_4160; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4257 = 7'h1f == total_offset_21[6:0] ? field_byte_21 : _GEN_4161; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4258 = 7'h20 == total_offset_21[6:0] ? field_byte_21 : _GEN_4162; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4259 = 7'h21 == total_offset_21[6:0] ? field_byte_21 : _GEN_4163; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4260 = 7'h22 == total_offset_21[6:0] ? field_byte_21 : _GEN_4164; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4261 = 7'h23 == total_offset_21[6:0] ? field_byte_21 : _GEN_4165; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4262 = 7'h24 == total_offset_21[6:0] ? field_byte_21 : _GEN_4166; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4263 = 7'h25 == total_offset_21[6:0] ? field_byte_21 : _GEN_4167; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4264 = 7'h26 == total_offset_21[6:0] ? field_byte_21 : _GEN_4168; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4265 = 7'h27 == total_offset_21[6:0] ? field_byte_21 : _GEN_4169; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4266 = 7'h28 == total_offset_21[6:0] ? field_byte_21 : _GEN_4170; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4267 = 7'h29 == total_offset_21[6:0] ? field_byte_21 : _GEN_4171; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4268 = 7'h2a == total_offset_21[6:0] ? field_byte_21 : _GEN_4172; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4269 = 7'h2b == total_offset_21[6:0] ? field_byte_21 : _GEN_4173; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4270 = 7'h2c == total_offset_21[6:0] ? field_byte_21 : _GEN_4174; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4271 = 7'h2d == total_offset_21[6:0] ? field_byte_21 : _GEN_4175; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4272 = 7'h2e == total_offset_21[6:0] ? field_byte_21 : _GEN_4176; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4273 = 7'h2f == total_offset_21[6:0] ? field_byte_21 : _GEN_4177; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4274 = 7'h30 == total_offset_21[6:0] ? field_byte_21 : _GEN_4178; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4275 = 7'h31 == total_offset_21[6:0] ? field_byte_21 : _GEN_4179; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4276 = 7'h32 == total_offset_21[6:0] ? field_byte_21 : _GEN_4180; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4277 = 7'h33 == total_offset_21[6:0] ? field_byte_21 : _GEN_4181; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4278 = 7'h34 == total_offset_21[6:0] ? field_byte_21 : _GEN_4182; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4279 = 7'h35 == total_offset_21[6:0] ? field_byte_21 : _GEN_4183; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4280 = 7'h36 == total_offset_21[6:0] ? field_byte_21 : _GEN_4184; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4281 = 7'h37 == total_offset_21[6:0] ? field_byte_21 : _GEN_4185; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4282 = 7'h38 == total_offset_21[6:0] ? field_byte_21 : _GEN_4186; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4283 = 7'h39 == total_offset_21[6:0] ? field_byte_21 : _GEN_4187; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4284 = 7'h3a == total_offset_21[6:0] ? field_byte_21 : _GEN_4188; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4285 = 7'h3b == total_offset_21[6:0] ? field_byte_21 : _GEN_4189; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4286 = 7'h3c == total_offset_21[6:0] ? field_byte_21 : _GEN_4190; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4287 = 7'h3d == total_offset_21[6:0] ? field_byte_21 : _GEN_4191; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4288 = 7'h3e == total_offset_21[6:0] ? field_byte_21 : _GEN_4192; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4289 = 7'h3f == total_offset_21[6:0] ? field_byte_21 : _GEN_4193; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4290 = 7'h40 == total_offset_21[6:0] ? field_byte_21 : _GEN_4194; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4291 = 7'h41 == total_offset_21[6:0] ? field_byte_21 : _GEN_4195; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4292 = 7'h42 == total_offset_21[6:0] ? field_byte_21 : _GEN_4196; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4293 = 7'h43 == total_offset_21[6:0] ? field_byte_21 : _GEN_4197; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4294 = 7'h44 == total_offset_21[6:0] ? field_byte_21 : _GEN_4198; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4295 = 7'h45 == total_offset_21[6:0] ? field_byte_21 : _GEN_4199; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4296 = 7'h46 == total_offset_21[6:0] ? field_byte_21 : _GEN_4200; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4297 = 7'h47 == total_offset_21[6:0] ? field_byte_21 : _GEN_4201; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4298 = 7'h48 == total_offset_21[6:0] ? field_byte_21 : _GEN_4202; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4299 = 7'h49 == total_offset_21[6:0] ? field_byte_21 : _GEN_4203; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4300 = 7'h4a == total_offset_21[6:0] ? field_byte_21 : _GEN_4204; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4301 = 7'h4b == total_offset_21[6:0] ? field_byte_21 : _GEN_4205; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4302 = 7'h4c == total_offset_21[6:0] ? field_byte_21 : _GEN_4206; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4303 = 7'h4d == total_offset_21[6:0] ? field_byte_21 : _GEN_4207; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4304 = 7'h4e == total_offset_21[6:0] ? field_byte_21 : _GEN_4208; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4305 = 7'h4f == total_offset_21[6:0] ? field_byte_21 : _GEN_4209; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4306 = 7'h50 == total_offset_21[6:0] ? field_byte_21 : _GEN_4210; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4307 = 7'h51 == total_offset_21[6:0] ? field_byte_21 : _GEN_4211; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4308 = 7'h52 == total_offset_21[6:0] ? field_byte_21 : _GEN_4212; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4309 = 7'h53 == total_offset_21[6:0] ? field_byte_21 : _GEN_4213; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4310 = 7'h54 == total_offset_21[6:0] ? field_byte_21 : _GEN_4214; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4311 = 7'h55 == total_offset_21[6:0] ? field_byte_21 : _GEN_4215; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4312 = 7'h56 == total_offset_21[6:0] ? field_byte_21 : _GEN_4216; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4313 = 7'h57 == total_offset_21[6:0] ? field_byte_21 : _GEN_4217; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4314 = 7'h58 == total_offset_21[6:0] ? field_byte_21 : _GEN_4218; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4315 = 7'h59 == total_offset_21[6:0] ? field_byte_21 : _GEN_4219; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4316 = 7'h5a == total_offset_21[6:0] ? field_byte_21 : _GEN_4220; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4317 = 7'h5b == total_offset_21[6:0] ? field_byte_21 : _GEN_4221; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4318 = 7'h5c == total_offset_21[6:0] ? field_byte_21 : _GEN_4222; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4319 = 7'h5d == total_offset_21[6:0] ? field_byte_21 : _GEN_4223; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4320 = 7'h5e == total_offset_21[6:0] ? field_byte_21 : _GEN_4224; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4321 = 7'h5f == total_offset_21[6:0] ? field_byte_21 : _GEN_4225; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4322 = 8'h5 < length_2 ? _GEN_4226 : _GEN_4130; // @[executor.scala 290:56]
  wire [7:0] _GEN_4323 = 8'h5 < length_2 ? _GEN_4227 : _GEN_4131; // @[executor.scala 290:56]
  wire [7:0] _GEN_4324 = 8'h5 < length_2 ? _GEN_4228 : _GEN_4132; // @[executor.scala 290:56]
  wire [7:0] _GEN_4325 = 8'h5 < length_2 ? _GEN_4229 : _GEN_4133; // @[executor.scala 290:56]
  wire [7:0] _GEN_4326 = 8'h5 < length_2 ? _GEN_4230 : _GEN_4134; // @[executor.scala 290:56]
  wire [7:0] _GEN_4327 = 8'h5 < length_2 ? _GEN_4231 : _GEN_4135; // @[executor.scala 290:56]
  wire [7:0] _GEN_4328 = 8'h5 < length_2 ? _GEN_4232 : _GEN_4136; // @[executor.scala 290:56]
  wire [7:0] _GEN_4329 = 8'h5 < length_2 ? _GEN_4233 : _GEN_4137; // @[executor.scala 290:56]
  wire [7:0] _GEN_4330 = 8'h5 < length_2 ? _GEN_4234 : _GEN_4138; // @[executor.scala 290:56]
  wire [7:0] _GEN_4331 = 8'h5 < length_2 ? _GEN_4235 : _GEN_4139; // @[executor.scala 290:56]
  wire [7:0] _GEN_4332 = 8'h5 < length_2 ? _GEN_4236 : _GEN_4140; // @[executor.scala 290:56]
  wire [7:0] _GEN_4333 = 8'h5 < length_2 ? _GEN_4237 : _GEN_4141; // @[executor.scala 290:56]
  wire [7:0] _GEN_4334 = 8'h5 < length_2 ? _GEN_4238 : _GEN_4142; // @[executor.scala 290:56]
  wire [7:0] _GEN_4335 = 8'h5 < length_2 ? _GEN_4239 : _GEN_4143; // @[executor.scala 290:56]
  wire [7:0] _GEN_4336 = 8'h5 < length_2 ? _GEN_4240 : _GEN_4144; // @[executor.scala 290:56]
  wire [7:0] _GEN_4337 = 8'h5 < length_2 ? _GEN_4241 : _GEN_4145; // @[executor.scala 290:56]
  wire [7:0] _GEN_4338 = 8'h5 < length_2 ? _GEN_4242 : _GEN_4146; // @[executor.scala 290:56]
  wire [7:0] _GEN_4339 = 8'h5 < length_2 ? _GEN_4243 : _GEN_4147; // @[executor.scala 290:56]
  wire [7:0] _GEN_4340 = 8'h5 < length_2 ? _GEN_4244 : _GEN_4148; // @[executor.scala 290:56]
  wire [7:0] _GEN_4341 = 8'h5 < length_2 ? _GEN_4245 : _GEN_4149; // @[executor.scala 290:56]
  wire [7:0] _GEN_4342 = 8'h5 < length_2 ? _GEN_4246 : _GEN_4150; // @[executor.scala 290:56]
  wire [7:0] _GEN_4343 = 8'h5 < length_2 ? _GEN_4247 : _GEN_4151; // @[executor.scala 290:56]
  wire [7:0] _GEN_4344 = 8'h5 < length_2 ? _GEN_4248 : _GEN_4152; // @[executor.scala 290:56]
  wire [7:0] _GEN_4345 = 8'h5 < length_2 ? _GEN_4249 : _GEN_4153; // @[executor.scala 290:56]
  wire [7:0] _GEN_4346 = 8'h5 < length_2 ? _GEN_4250 : _GEN_4154; // @[executor.scala 290:56]
  wire [7:0] _GEN_4347 = 8'h5 < length_2 ? _GEN_4251 : _GEN_4155; // @[executor.scala 290:56]
  wire [7:0] _GEN_4348 = 8'h5 < length_2 ? _GEN_4252 : _GEN_4156; // @[executor.scala 290:56]
  wire [7:0] _GEN_4349 = 8'h5 < length_2 ? _GEN_4253 : _GEN_4157; // @[executor.scala 290:56]
  wire [7:0] _GEN_4350 = 8'h5 < length_2 ? _GEN_4254 : _GEN_4158; // @[executor.scala 290:56]
  wire [7:0] _GEN_4351 = 8'h5 < length_2 ? _GEN_4255 : _GEN_4159; // @[executor.scala 290:56]
  wire [7:0] _GEN_4352 = 8'h5 < length_2 ? _GEN_4256 : _GEN_4160; // @[executor.scala 290:56]
  wire [7:0] _GEN_4353 = 8'h5 < length_2 ? _GEN_4257 : _GEN_4161; // @[executor.scala 290:56]
  wire [7:0] _GEN_4354 = 8'h5 < length_2 ? _GEN_4258 : _GEN_4162; // @[executor.scala 290:56]
  wire [7:0] _GEN_4355 = 8'h5 < length_2 ? _GEN_4259 : _GEN_4163; // @[executor.scala 290:56]
  wire [7:0] _GEN_4356 = 8'h5 < length_2 ? _GEN_4260 : _GEN_4164; // @[executor.scala 290:56]
  wire [7:0] _GEN_4357 = 8'h5 < length_2 ? _GEN_4261 : _GEN_4165; // @[executor.scala 290:56]
  wire [7:0] _GEN_4358 = 8'h5 < length_2 ? _GEN_4262 : _GEN_4166; // @[executor.scala 290:56]
  wire [7:0] _GEN_4359 = 8'h5 < length_2 ? _GEN_4263 : _GEN_4167; // @[executor.scala 290:56]
  wire [7:0] _GEN_4360 = 8'h5 < length_2 ? _GEN_4264 : _GEN_4168; // @[executor.scala 290:56]
  wire [7:0] _GEN_4361 = 8'h5 < length_2 ? _GEN_4265 : _GEN_4169; // @[executor.scala 290:56]
  wire [7:0] _GEN_4362 = 8'h5 < length_2 ? _GEN_4266 : _GEN_4170; // @[executor.scala 290:56]
  wire [7:0] _GEN_4363 = 8'h5 < length_2 ? _GEN_4267 : _GEN_4171; // @[executor.scala 290:56]
  wire [7:0] _GEN_4364 = 8'h5 < length_2 ? _GEN_4268 : _GEN_4172; // @[executor.scala 290:56]
  wire [7:0] _GEN_4365 = 8'h5 < length_2 ? _GEN_4269 : _GEN_4173; // @[executor.scala 290:56]
  wire [7:0] _GEN_4366 = 8'h5 < length_2 ? _GEN_4270 : _GEN_4174; // @[executor.scala 290:56]
  wire [7:0] _GEN_4367 = 8'h5 < length_2 ? _GEN_4271 : _GEN_4175; // @[executor.scala 290:56]
  wire [7:0] _GEN_4368 = 8'h5 < length_2 ? _GEN_4272 : _GEN_4176; // @[executor.scala 290:56]
  wire [7:0] _GEN_4369 = 8'h5 < length_2 ? _GEN_4273 : _GEN_4177; // @[executor.scala 290:56]
  wire [7:0] _GEN_4370 = 8'h5 < length_2 ? _GEN_4274 : _GEN_4178; // @[executor.scala 290:56]
  wire [7:0] _GEN_4371 = 8'h5 < length_2 ? _GEN_4275 : _GEN_4179; // @[executor.scala 290:56]
  wire [7:0] _GEN_4372 = 8'h5 < length_2 ? _GEN_4276 : _GEN_4180; // @[executor.scala 290:56]
  wire [7:0] _GEN_4373 = 8'h5 < length_2 ? _GEN_4277 : _GEN_4181; // @[executor.scala 290:56]
  wire [7:0] _GEN_4374 = 8'h5 < length_2 ? _GEN_4278 : _GEN_4182; // @[executor.scala 290:56]
  wire [7:0] _GEN_4375 = 8'h5 < length_2 ? _GEN_4279 : _GEN_4183; // @[executor.scala 290:56]
  wire [7:0] _GEN_4376 = 8'h5 < length_2 ? _GEN_4280 : _GEN_4184; // @[executor.scala 290:56]
  wire [7:0] _GEN_4377 = 8'h5 < length_2 ? _GEN_4281 : _GEN_4185; // @[executor.scala 290:56]
  wire [7:0] _GEN_4378 = 8'h5 < length_2 ? _GEN_4282 : _GEN_4186; // @[executor.scala 290:56]
  wire [7:0] _GEN_4379 = 8'h5 < length_2 ? _GEN_4283 : _GEN_4187; // @[executor.scala 290:56]
  wire [7:0] _GEN_4380 = 8'h5 < length_2 ? _GEN_4284 : _GEN_4188; // @[executor.scala 290:56]
  wire [7:0] _GEN_4381 = 8'h5 < length_2 ? _GEN_4285 : _GEN_4189; // @[executor.scala 290:56]
  wire [7:0] _GEN_4382 = 8'h5 < length_2 ? _GEN_4286 : _GEN_4190; // @[executor.scala 290:56]
  wire [7:0] _GEN_4383 = 8'h5 < length_2 ? _GEN_4287 : _GEN_4191; // @[executor.scala 290:56]
  wire [7:0] _GEN_4384 = 8'h5 < length_2 ? _GEN_4288 : _GEN_4192; // @[executor.scala 290:56]
  wire [7:0] _GEN_4385 = 8'h5 < length_2 ? _GEN_4289 : _GEN_4193; // @[executor.scala 290:56]
  wire [7:0] _GEN_4386 = 8'h5 < length_2 ? _GEN_4290 : _GEN_4194; // @[executor.scala 290:56]
  wire [7:0] _GEN_4387 = 8'h5 < length_2 ? _GEN_4291 : _GEN_4195; // @[executor.scala 290:56]
  wire [7:0] _GEN_4388 = 8'h5 < length_2 ? _GEN_4292 : _GEN_4196; // @[executor.scala 290:56]
  wire [7:0] _GEN_4389 = 8'h5 < length_2 ? _GEN_4293 : _GEN_4197; // @[executor.scala 290:56]
  wire [7:0] _GEN_4390 = 8'h5 < length_2 ? _GEN_4294 : _GEN_4198; // @[executor.scala 290:56]
  wire [7:0] _GEN_4391 = 8'h5 < length_2 ? _GEN_4295 : _GEN_4199; // @[executor.scala 290:56]
  wire [7:0] _GEN_4392 = 8'h5 < length_2 ? _GEN_4296 : _GEN_4200; // @[executor.scala 290:56]
  wire [7:0] _GEN_4393 = 8'h5 < length_2 ? _GEN_4297 : _GEN_4201; // @[executor.scala 290:56]
  wire [7:0] _GEN_4394 = 8'h5 < length_2 ? _GEN_4298 : _GEN_4202; // @[executor.scala 290:56]
  wire [7:0] _GEN_4395 = 8'h5 < length_2 ? _GEN_4299 : _GEN_4203; // @[executor.scala 290:56]
  wire [7:0] _GEN_4396 = 8'h5 < length_2 ? _GEN_4300 : _GEN_4204; // @[executor.scala 290:56]
  wire [7:0] _GEN_4397 = 8'h5 < length_2 ? _GEN_4301 : _GEN_4205; // @[executor.scala 290:56]
  wire [7:0] _GEN_4398 = 8'h5 < length_2 ? _GEN_4302 : _GEN_4206; // @[executor.scala 290:56]
  wire [7:0] _GEN_4399 = 8'h5 < length_2 ? _GEN_4303 : _GEN_4207; // @[executor.scala 290:56]
  wire [7:0] _GEN_4400 = 8'h5 < length_2 ? _GEN_4304 : _GEN_4208; // @[executor.scala 290:56]
  wire [7:0] _GEN_4401 = 8'h5 < length_2 ? _GEN_4305 : _GEN_4209; // @[executor.scala 290:56]
  wire [7:0] _GEN_4402 = 8'h5 < length_2 ? _GEN_4306 : _GEN_4210; // @[executor.scala 290:56]
  wire [7:0] _GEN_4403 = 8'h5 < length_2 ? _GEN_4307 : _GEN_4211; // @[executor.scala 290:56]
  wire [7:0] _GEN_4404 = 8'h5 < length_2 ? _GEN_4308 : _GEN_4212; // @[executor.scala 290:56]
  wire [7:0] _GEN_4405 = 8'h5 < length_2 ? _GEN_4309 : _GEN_4213; // @[executor.scala 290:56]
  wire [7:0] _GEN_4406 = 8'h5 < length_2 ? _GEN_4310 : _GEN_4214; // @[executor.scala 290:56]
  wire [7:0] _GEN_4407 = 8'h5 < length_2 ? _GEN_4311 : _GEN_4215; // @[executor.scala 290:56]
  wire [7:0] _GEN_4408 = 8'h5 < length_2 ? _GEN_4312 : _GEN_4216; // @[executor.scala 290:56]
  wire [7:0] _GEN_4409 = 8'h5 < length_2 ? _GEN_4313 : _GEN_4217; // @[executor.scala 290:56]
  wire [7:0] _GEN_4410 = 8'h5 < length_2 ? _GEN_4314 : _GEN_4218; // @[executor.scala 290:56]
  wire [7:0] _GEN_4411 = 8'h5 < length_2 ? _GEN_4315 : _GEN_4219; // @[executor.scala 290:56]
  wire [7:0] _GEN_4412 = 8'h5 < length_2 ? _GEN_4316 : _GEN_4220; // @[executor.scala 290:56]
  wire [7:0] _GEN_4413 = 8'h5 < length_2 ? _GEN_4317 : _GEN_4221; // @[executor.scala 290:56]
  wire [7:0] _GEN_4414 = 8'h5 < length_2 ? _GEN_4318 : _GEN_4222; // @[executor.scala 290:56]
  wire [7:0] _GEN_4415 = 8'h5 < length_2 ? _GEN_4319 : _GEN_4223; // @[executor.scala 290:56]
  wire [7:0] _GEN_4416 = 8'h5 < length_2 ? _GEN_4320 : _GEN_4224; // @[executor.scala 290:56]
  wire [7:0] _GEN_4417 = 8'h5 < length_2 ? _GEN_4321 : _GEN_4225; // @[executor.scala 290:56]
  wire [7:0] field_byte_22 = field_2[15:8]; // @[executor.scala 287:53]
  wire [7:0] total_offset_22 = offset_2 + 8'h6; // @[executor.scala 289:53]
  wire [7:0] _GEN_4418 = 7'h0 == total_offset_22[6:0] ? field_byte_22 : _GEN_4322; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4419 = 7'h1 == total_offset_22[6:0] ? field_byte_22 : _GEN_4323; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4420 = 7'h2 == total_offset_22[6:0] ? field_byte_22 : _GEN_4324; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4421 = 7'h3 == total_offset_22[6:0] ? field_byte_22 : _GEN_4325; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4422 = 7'h4 == total_offset_22[6:0] ? field_byte_22 : _GEN_4326; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4423 = 7'h5 == total_offset_22[6:0] ? field_byte_22 : _GEN_4327; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4424 = 7'h6 == total_offset_22[6:0] ? field_byte_22 : _GEN_4328; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4425 = 7'h7 == total_offset_22[6:0] ? field_byte_22 : _GEN_4329; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4426 = 7'h8 == total_offset_22[6:0] ? field_byte_22 : _GEN_4330; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4427 = 7'h9 == total_offset_22[6:0] ? field_byte_22 : _GEN_4331; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4428 = 7'ha == total_offset_22[6:0] ? field_byte_22 : _GEN_4332; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4429 = 7'hb == total_offset_22[6:0] ? field_byte_22 : _GEN_4333; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4430 = 7'hc == total_offset_22[6:0] ? field_byte_22 : _GEN_4334; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4431 = 7'hd == total_offset_22[6:0] ? field_byte_22 : _GEN_4335; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4432 = 7'he == total_offset_22[6:0] ? field_byte_22 : _GEN_4336; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4433 = 7'hf == total_offset_22[6:0] ? field_byte_22 : _GEN_4337; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4434 = 7'h10 == total_offset_22[6:0] ? field_byte_22 : _GEN_4338; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4435 = 7'h11 == total_offset_22[6:0] ? field_byte_22 : _GEN_4339; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4436 = 7'h12 == total_offset_22[6:0] ? field_byte_22 : _GEN_4340; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4437 = 7'h13 == total_offset_22[6:0] ? field_byte_22 : _GEN_4341; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4438 = 7'h14 == total_offset_22[6:0] ? field_byte_22 : _GEN_4342; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4439 = 7'h15 == total_offset_22[6:0] ? field_byte_22 : _GEN_4343; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4440 = 7'h16 == total_offset_22[6:0] ? field_byte_22 : _GEN_4344; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4441 = 7'h17 == total_offset_22[6:0] ? field_byte_22 : _GEN_4345; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4442 = 7'h18 == total_offset_22[6:0] ? field_byte_22 : _GEN_4346; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4443 = 7'h19 == total_offset_22[6:0] ? field_byte_22 : _GEN_4347; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4444 = 7'h1a == total_offset_22[6:0] ? field_byte_22 : _GEN_4348; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4445 = 7'h1b == total_offset_22[6:0] ? field_byte_22 : _GEN_4349; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4446 = 7'h1c == total_offset_22[6:0] ? field_byte_22 : _GEN_4350; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4447 = 7'h1d == total_offset_22[6:0] ? field_byte_22 : _GEN_4351; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4448 = 7'h1e == total_offset_22[6:0] ? field_byte_22 : _GEN_4352; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4449 = 7'h1f == total_offset_22[6:0] ? field_byte_22 : _GEN_4353; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4450 = 7'h20 == total_offset_22[6:0] ? field_byte_22 : _GEN_4354; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4451 = 7'h21 == total_offset_22[6:0] ? field_byte_22 : _GEN_4355; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4452 = 7'h22 == total_offset_22[6:0] ? field_byte_22 : _GEN_4356; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4453 = 7'h23 == total_offset_22[6:0] ? field_byte_22 : _GEN_4357; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4454 = 7'h24 == total_offset_22[6:0] ? field_byte_22 : _GEN_4358; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4455 = 7'h25 == total_offset_22[6:0] ? field_byte_22 : _GEN_4359; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4456 = 7'h26 == total_offset_22[6:0] ? field_byte_22 : _GEN_4360; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4457 = 7'h27 == total_offset_22[6:0] ? field_byte_22 : _GEN_4361; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4458 = 7'h28 == total_offset_22[6:0] ? field_byte_22 : _GEN_4362; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4459 = 7'h29 == total_offset_22[6:0] ? field_byte_22 : _GEN_4363; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4460 = 7'h2a == total_offset_22[6:0] ? field_byte_22 : _GEN_4364; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4461 = 7'h2b == total_offset_22[6:0] ? field_byte_22 : _GEN_4365; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4462 = 7'h2c == total_offset_22[6:0] ? field_byte_22 : _GEN_4366; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4463 = 7'h2d == total_offset_22[6:0] ? field_byte_22 : _GEN_4367; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4464 = 7'h2e == total_offset_22[6:0] ? field_byte_22 : _GEN_4368; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4465 = 7'h2f == total_offset_22[6:0] ? field_byte_22 : _GEN_4369; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4466 = 7'h30 == total_offset_22[6:0] ? field_byte_22 : _GEN_4370; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4467 = 7'h31 == total_offset_22[6:0] ? field_byte_22 : _GEN_4371; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4468 = 7'h32 == total_offset_22[6:0] ? field_byte_22 : _GEN_4372; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4469 = 7'h33 == total_offset_22[6:0] ? field_byte_22 : _GEN_4373; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4470 = 7'h34 == total_offset_22[6:0] ? field_byte_22 : _GEN_4374; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4471 = 7'h35 == total_offset_22[6:0] ? field_byte_22 : _GEN_4375; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4472 = 7'h36 == total_offset_22[6:0] ? field_byte_22 : _GEN_4376; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4473 = 7'h37 == total_offset_22[6:0] ? field_byte_22 : _GEN_4377; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4474 = 7'h38 == total_offset_22[6:0] ? field_byte_22 : _GEN_4378; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4475 = 7'h39 == total_offset_22[6:0] ? field_byte_22 : _GEN_4379; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4476 = 7'h3a == total_offset_22[6:0] ? field_byte_22 : _GEN_4380; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4477 = 7'h3b == total_offset_22[6:0] ? field_byte_22 : _GEN_4381; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4478 = 7'h3c == total_offset_22[6:0] ? field_byte_22 : _GEN_4382; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4479 = 7'h3d == total_offset_22[6:0] ? field_byte_22 : _GEN_4383; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4480 = 7'h3e == total_offset_22[6:0] ? field_byte_22 : _GEN_4384; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4481 = 7'h3f == total_offset_22[6:0] ? field_byte_22 : _GEN_4385; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4482 = 7'h40 == total_offset_22[6:0] ? field_byte_22 : _GEN_4386; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4483 = 7'h41 == total_offset_22[6:0] ? field_byte_22 : _GEN_4387; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4484 = 7'h42 == total_offset_22[6:0] ? field_byte_22 : _GEN_4388; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4485 = 7'h43 == total_offset_22[6:0] ? field_byte_22 : _GEN_4389; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4486 = 7'h44 == total_offset_22[6:0] ? field_byte_22 : _GEN_4390; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4487 = 7'h45 == total_offset_22[6:0] ? field_byte_22 : _GEN_4391; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4488 = 7'h46 == total_offset_22[6:0] ? field_byte_22 : _GEN_4392; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4489 = 7'h47 == total_offset_22[6:0] ? field_byte_22 : _GEN_4393; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4490 = 7'h48 == total_offset_22[6:0] ? field_byte_22 : _GEN_4394; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4491 = 7'h49 == total_offset_22[6:0] ? field_byte_22 : _GEN_4395; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4492 = 7'h4a == total_offset_22[6:0] ? field_byte_22 : _GEN_4396; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4493 = 7'h4b == total_offset_22[6:0] ? field_byte_22 : _GEN_4397; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4494 = 7'h4c == total_offset_22[6:0] ? field_byte_22 : _GEN_4398; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4495 = 7'h4d == total_offset_22[6:0] ? field_byte_22 : _GEN_4399; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4496 = 7'h4e == total_offset_22[6:0] ? field_byte_22 : _GEN_4400; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4497 = 7'h4f == total_offset_22[6:0] ? field_byte_22 : _GEN_4401; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4498 = 7'h50 == total_offset_22[6:0] ? field_byte_22 : _GEN_4402; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4499 = 7'h51 == total_offset_22[6:0] ? field_byte_22 : _GEN_4403; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4500 = 7'h52 == total_offset_22[6:0] ? field_byte_22 : _GEN_4404; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4501 = 7'h53 == total_offset_22[6:0] ? field_byte_22 : _GEN_4405; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4502 = 7'h54 == total_offset_22[6:0] ? field_byte_22 : _GEN_4406; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4503 = 7'h55 == total_offset_22[6:0] ? field_byte_22 : _GEN_4407; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4504 = 7'h56 == total_offset_22[6:0] ? field_byte_22 : _GEN_4408; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4505 = 7'h57 == total_offset_22[6:0] ? field_byte_22 : _GEN_4409; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4506 = 7'h58 == total_offset_22[6:0] ? field_byte_22 : _GEN_4410; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4507 = 7'h59 == total_offset_22[6:0] ? field_byte_22 : _GEN_4411; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4508 = 7'h5a == total_offset_22[6:0] ? field_byte_22 : _GEN_4412; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4509 = 7'h5b == total_offset_22[6:0] ? field_byte_22 : _GEN_4413; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4510 = 7'h5c == total_offset_22[6:0] ? field_byte_22 : _GEN_4414; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4511 = 7'h5d == total_offset_22[6:0] ? field_byte_22 : _GEN_4415; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4512 = 7'h5e == total_offset_22[6:0] ? field_byte_22 : _GEN_4416; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4513 = 7'h5f == total_offset_22[6:0] ? field_byte_22 : _GEN_4417; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4514 = 8'h6 < length_2 ? _GEN_4418 : _GEN_4322; // @[executor.scala 290:56]
  wire [7:0] _GEN_4515 = 8'h6 < length_2 ? _GEN_4419 : _GEN_4323; // @[executor.scala 290:56]
  wire [7:0] _GEN_4516 = 8'h6 < length_2 ? _GEN_4420 : _GEN_4324; // @[executor.scala 290:56]
  wire [7:0] _GEN_4517 = 8'h6 < length_2 ? _GEN_4421 : _GEN_4325; // @[executor.scala 290:56]
  wire [7:0] _GEN_4518 = 8'h6 < length_2 ? _GEN_4422 : _GEN_4326; // @[executor.scala 290:56]
  wire [7:0] _GEN_4519 = 8'h6 < length_2 ? _GEN_4423 : _GEN_4327; // @[executor.scala 290:56]
  wire [7:0] _GEN_4520 = 8'h6 < length_2 ? _GEN_4424 : _GEN_4328; // @[executor.scala 290:56]
  wire [7:0] _GEN_4521 = 8'h6 < length_2 ? _GEN_4425 : _GEN_4329; // @[executor.scala 290:56]
  wire [7:0] _GEN_4522 = 8'h6 < length_2 ? _GEN_4426 : _GEN_4330; // @[executor.scala 290:56]
  wire [7:0] _GEN_4523 = 8'h6 < length_2 ? _GEN_4427 : _GEN_4331; // @[executor.scala 290:56]
  wire [7:0] _GEN_4524 = 8'h6 < length_2 ? _GEN_4428 : _GEN_4332; // @[executor.scala 290:56]
  wire [7:0] _GEN_4525 = 8'h6 < length_2 ? _GEN_4429 : _GEN_4333; // @[executor.scala 290:56]
  wire [7:0] _GEN_4526 = 8'h6 < length_2 ? _GEN_4430 : _GEN_4334; // @[executor.scala 290:56]
  wire [7:0] _GEN_4527 = 8'h6 < length_2 ? _GEN_4431 : _GEN_4335; // @[executor.scala 290:56]
  wire [7:0] _GEN_4528 = 8'h6 < length_2 ? _GEN_4432 : _GEN_4336; // @[executor.scala 290:56]
  wire [7:0] _GEN_4529 = 8'h6 < length_2 ? _GEN_4433 : _GEN_4337; // @[executor.scala 290:56]
  wire [7:0] _GEN_4530 = 8'h6 < length_2 ? _GEN_4434 : _GEN_4338; // @[executor.scala 290:56]
  wire [7:0] _GEN_4531 = 8'h6 < length_2 ? _GEN_4435 : _GEN_4339; // @[executor.scala 290:56]
  wire [7:0] _GEN_4532 = 8'h6 < length_2 ? _GEN_4436 : _GEN_4340; // @[executor.scala 290:56]
  wire [7:0] _GEN_4533 = 8'h6 < length_2 ? _GEN_4437 : _GEN_4341; // @[executor.scala 290:56]
  wire [7:0] _GEN_4534 = 8'h6 < length_2 ? _GEN_4438 : _GEN_4342; // @[executor.scala 290:56]
  wire [7:0] _GEN_4535 = 8'h6 < length_2 ? _GEN_4439 : _GEN_4343; // @[executor.scala 290:56]
  wire [7:0] _GEN_4536 = 8'h6 < length_2 ? _GEN_4440 : _GEN_4344; // @[executor.scala 290:56]
  wire [7:0] _GEN_4537 = 8'h6 < length_2 ? _GEN_4441 : _GEN_4345; // @[executor.scala 290:56]
  wire [7:0] _GEN_4538 = 8'h6 < length_2 ? _GEN_4442 : _GEN_4346; // @[executor.scala 290:56]
  wire [7:0] _GEN_4539 = 8'h6 < length_2 ? _GEN_4443 : _GEN_4347; // @[executor.scala 290:56]
  wire [7:0] _GEN_4540 = 8'h6 < length_2 ? _GEN_4444 : _GEN_4348; // @[executor.scala 290:56]
  wire [7:0] _GEN_4541 = 8'h6 < length_2 ? _GEN_4445 : _GEN_4349; // @[executor.scala 290:56]
  wire [7:0] _GEN_4542 = 8'h6 < length_2 ? _GEN_4446 : _GEN_4350; // @[executor.scala 290:56]
  wire [7:0] _GEN_4543 = 8'h6 < length_2 ? _GEN_4447 : _GEN_4351; // @[executor.scala 290:56]
  wire [7:0] _GEN_4544 = 8'h6 < length_2 ? _GEN_4448 : _GEN_4352; // @[executor.scala 290:56]
  wire [7:0] _GEN_4545 = 8'h6 < length_2 ? _GEN_4449 : _GEN_4353; // @[executor.scala 290:56]
  wire [7:0] _GEN_4546 = 8'h6 < length_2 ? _GEN_4450 : _GEN_4354; // @[executor.scala 290:56]
  wire [7:0] _GEN_4547 = 8'h6 < length_2 ? _GEN_4451 : _GEN_4355; // @[executor.scala 290:56]
  wire [7:0] _GEN_4548 = 8'h6 < length_2 ? _GEN_4452 : _GEN_4356; // @[executor.scala 290:56]
  wire [7:0] _GEN_4549 = 8'h6 < length_2 ? _GEN_4453 : _GEN_4357; // @[executor.scala 290:56]
  wire [7:0] _GEN_4550 = 8'h6 < length_2 ? _GEN_4454 : _GEN_4358; // @[executor.scala 290:56]
  wire [7:0] _GEN_4551 = 8'h6 < length_2 ? _GEN_4455 : _GEN_4359; // @[executor.scala 290:56]
  wire [7:0] _GEN_4552 = 8'h6 < length_2 ? _GEN_4456 : _GEN_4360; // @[executor.scala 290:56]
  wire [7:0] _GEN_4553 = 8'h6 < length_2 ? _GEN_4457 : _GEN_4361; // @[executor.scala 290:56]
  wire [7:0] _GEN_4554 = 8'h6 < length_2 ? _GEN_4458 : _GEN_4362; // @[executor.scala 290:56]
  wire [7:0] _GEN_4555 = 8'h6 < length_2 ? _GEN_4459 : _GEN_4363; // @[executor.scala 290:56]
  wire [7:0] _GEN_4556 = 8'h6 < length_2 ? _GEN_4460 : _GEN_4364; // @[executor.scala 290:56]
  wire [7:0] _GEN_4557 = 8'h6 < length_2 ? _GEN_4461 : _GEN_4365; // @[executor.scala 290:56]
  wire [7:0] _GEN_4558 = 8'h6 < length_2 ? _GEN_4462 : _GEN_4366; // @[executor.scala 290:56]
  wire [7:0] _GEN_4559 = 8'h6 < length_2 ? _GEN_4463 : _GEN_4367; // @[executor.scala 290:56]
  wire [7:0] _GEN_4560 = 8'h6 < length_2 ? _GEN_4464 : _GEN_4368; // @[executor.scala 290:56]
  wire [7:0] _GEN_4561 = 8'h6 < length_2 ? _GEN_4465 : _GEN_4369; // @[executor.scala 290:56]
  wire [7:0] _GEN_4562 = 8'h6 < length_2 ? _GEN_4466 : _GEN_4370; // @[executor.scala 290:56]
  wire [7:0] _GEN_4563 = 8'h6 < length_2 ? _GEN_4467 : _GEN_4371; // @[executor.scala 290:56]
  wire [7:0] _GEN_4564 = 8'h6 < length_2 ? _GEN_4468 : _GEN_4372; // @[executor.scala 290:56]
  wire [7:0] _GEN_4565 = 8'h6 < length_2 ? _GEN_4469 : _GEN_4373; // @[executor.scala 290:56]
  wire [7:0] _GEN_4566 = 8'h6 < length_2 ? _GEN_4470 : _GEN_4374; // @[executor.scala 290:56]
  wire [7:0] _GEN_4567 = 8'h6 < length_2 ? _GEN_4471 : _GEN_4375; // @[executor.scala 290:56]
  wire [7:0] _GEN_4568 = 8'h6 < length_2 ? _GEN_4472 : _GEN_4376; // @[executor.scala 290:56]
  wire [7:0] _GEN_4569 = 8'h6 < length_2 ? _GEN_4473 : _GEN_4377; // @[executor.scala 290:56]
  wire [7:0] _GEN_4570 = 8'h6 < length_2 ? _GEN_4474 : _GEN_4378; // @[executor.scala 290:56]
  wire [7:0] _GEN_4571 = 8'h6 < length_2 ? _GEN_4475 : _GEN_4379; // @[executor.scala 290:56]
  wire [7:0] _GEN_4572 = 8'h6 < length_2 ? _GEN_4476 : _GEN_4380; // @[executor.scala 290:56]
  wire [7:0] _GEN_4573 = 8'h6 < length_2 ? _GEN_4477 : _GEN_4381; // @[executor.scala 290:56]
  wire [7:0] _GEN_4574 = 8'h6 < length_2 ? _GEN_4478 : _GEN_4382; // @[executor.scala 290:56]
  wire [7:0] _GEN_4575 = 8'h6 < length_2 ? _GEN_4479 : _GEN_4383; // @[executor.scala 290:56]
  wire [7:0] _GEN_4576 = 8'h6 < length_2 ? _GEN_4480 : _GEN_4384; // @[executor.scala 290:56]
  wire [7:0] _GEN_4577 = 8'h6 < length_2 ? _GEN_4481 : _GEN_4385; // @[executor.scala 290:56]
  wire [7:0] _GEN_4578 = 8'h6 < length_2 ? _GEN_4482 : _GEN_4386; // @[executor.scala 290:56]
  wire [7:0] _GEN_4579 = 8'h6 < length_2 ? _GEN_4483 : _GEN_4387; // @[executor.scala 290:56]
  wire [7:0] _GEN_4580 = 8'h6 < length_2 ? _GEN_4484 : _GEN_4388; // @[executor.scala 290:56]
  wire [7:0] _GEN_4581 = 8'h6 < length_2 ? _GEN_4485 : _GEN_4389; // @[executor.scala 290:56]
  wire [7:0] _GEN_4582 = 8'h6 < length_2 ? _GEN_4486 : _GEN_4390; // @[executor.scala 290:56]
  wire [7:0] _GEN_4583 = 8'h6 < length_2 ? _GEN_4487 : _GEN_4391; // @[executor.scala 290:56]
  wire [7:0] _GEN_4584 = 8'h6 < length_2 ? _GEN_4488 : _GEN_4392; // @[executor.scala 290:56]
  wire [7:0] _GEN_4585 = 8'h6 < length_2 ? _GEN_4489 : _GEN_4393; // @[executor.scala 290:56]
  wire [7:0] _GEN_4586 = 8'h6 < length_2 ? _GEN_4490 : _GEN_4394; // @[executor.scala 290:56]
  wire [7:0] _GEN_4587 = 8'h6 < length_2 ? _GEN_4491 : _GEN_4395; // @[executor.scala 290:56]
  wire [7:0] _GEN_4588 = 8'h6 < length_2 ? _GEN_4492 : _GEN_4396; // @[executor.scala 290:56]
  wire [7:0] _GEN_4589 = 8'h6 < length_2 ? _GEN_4493 : _GEN_4397; // @[executor.scala 290:56]
  wire [7:0] _GEN_4590 = 8'h6 < length_2 ? _GEN_4494 : _GEN_4398; // @[executor.scala 290:56]
  wire [7:0] _GEN_4591 = 8'h6 < length_2 ? _GEN_4495 : _GEN_4399; // @[executor.scala 290:56]
  wire [7:0] _GEN_4592 = 8'h6 < length_2 ? _GEN_4496 : _GEN_4400; // @[executor.scala 290:56]
  wire [7:0] _GEN_4593 = 8'h6 < length_2 ? _GEN_4497 : _GEN_4401; // @[executor.scala 290:56]
  wire [7:0] _GEN_4594 = 8'h6 < length_2 ? _GEN_4498 : _GEN_4402; // @[executor.scala 290:56]
  wire [7:0] _GEN_4595 = 8'h6 < length_2 ? _GEN_4499 : _GEN_4403; // @[executor.scala 290:56]
  wire [7:0] _GEN_4596 = 8'h6 < length_2 ? _GEN_4500 : _GEN_4404; // @[executor.scala 290:56]
  wire [7:0] _GEN_4597 = 8'h6 < length_2 ? _GEN_4501 : _GEN_4405; // @[executor.scala 290:56]
  wire [7:0] _GEN_4598 = 8'h6 < length_2 ? _GEN_4502 : _GEN_4406; // @[executor.scala 290:56]
  wire [7:0] _GEN_4599 = 8'h6 < length_2 ? _GEN_4503 : _GEN_4407; // @[executor.scala 290:56]
  wire [7:0] _GEN_4600 = 8'h6 < length_2 ? _GEN_4504 : _GEN_4408; // @[executor.scala 290:56]
  wire [7:0] _GEN_4601 = 8'h6 < length_2 ? _GEN_4505 : _GEN_4409; // @[executor.scala 290:56]
  wire [7:0] _GEN_4602 = 8'h6 < length_2 ? _GEN_4506 : _GEN_4410; // @[executor.scala 290:56]
  wire [7:0] _GEN_4603 = 8'h6 < length_2 ? _GEN_4507 : _GEN_4411; // @[executor.scala 290:56]
  wire [7:0] _GEN_4604 = 8'h6 < length_2 ? _GEN_4508 : _GEN_4412; // @[executor.scala 290:56]
  wire [7:0] _GEN_4605 = 8'h6 < length_2 ? _GEN_4509 : _GEN_4413; // @[executor.scala 290:56]
  wire [7:0] _GEN_4606 = 8'h6 < length_2 ? _GEN_4510 : _GEN_4414; // @[executor.scala 290:56]
  wire [7:0] _GEN_4607 = 8'h6 < length_2 ? _GEN_4511 : _GEN_4415; // @[executor.scala 290:56]
  wire [7:0] _GEN_4608 = 8'h6 < length_2 ? _GEN_4512 : _GEN_4416; // @[executor.scala 290:56]
  wire [7:0] _GEN_4609 = 8'h6 < length_2 ? _GEN_4513 : _GEN_4417; // @[executor.scala 290:56]
  wire [7:0] field_byte_23 = field_2[7:0]; // @[executor.scala 287:53]
  wire [7:0] total_offset_23 = offset_2 + 8'h7; // @[executor.scala 289:53]
  wire [7:0] _GEN_4610 = 7'h0 == total_offset_23[6:0] ? field_byte_23 : _GEN_4514; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4611 = 7'h1 == total_offset_23[6:0] ? field_byte_23 : _GEN_4515; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4612 = 7'h2 == total_offset_23[6:0] ? field_byte_23 : _GEN_4516; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4613 = 7'h3 == total_offset_23[6:0] ? field_byte_23 : _GEN_4517; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4614 = 7'h4 == total_offset_23[6:0] ? field_byte_23 : _GEN_4518; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4615 = 7'h5 == total_offset_23[6:0] ? field_byte_23 : _GEN_4519; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4616 = 7'h6 == total_offset_23[6:0] ? field_byte_23 : _GEN_4520; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4617 = 7'h7 == total_offset_23[6:0] ? field_byte_23 : _GEN_4521; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4618 = 7'h8 == total_offset_23[6:0] ? field_byte_23 : _GEN_4522; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4619 = 7'h9 == total_offset_23[6:0] ? field_byte_23 : _GEN_4523; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4620 = 7'ha == total_offset_23[6:0] ? field_byte_23 : _GEN_4524; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4621 = 7'hb == total_offset_23[6:0] ? field_byte_23 : _GEN_4525; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4622 = 7'hc == total_offset_23[6:0] ? field_byte_23 : _GEN_4526; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4623 = 7'hd == total_offset_23[6:0] ? field_byte_23 : _GEN_4527; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4624 = 7'he == total_offset_23[6:0] ? field_byte_23 : _GEN_4528; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4625 = 7'hf == total_offset_23[6:0] ? field_byte_23 : _GEN_4529; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4626 = 7'h10 == total_offset_23[6:0] ? field_byte_23 : _GEN_4530; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4627 = 7'h11 == total_offset_23[6:0] ? field_byte_23 : _GEN_4531; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4628 = 7'h12 == total_offset_23[6:0] ? field_byte_23 : _GEN_4532; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4629 = 7'h13 == total_offset_23[6:0] ? field_byte_23 : _GEN_4533; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4630 = 7'h14 == total_offset_23[6:0] ? field_byte_23 : _GEN_4534; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4631 = 7'h15 == total_offset_23[6:0] ? field_byte_23 : _GEN_4535; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4632 = 7'h16 == total_offset_23[6:0] ? field_byte_23 : _GEN_4536; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4633 = 7'h17 == total_offset_23[6:0] ? field_byte_23 : _GEN_4537; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4634 = 7'h18 == total_offset_23[6:0] ? field_byte_23 : _GEN_4538; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4635 = 7'h19 == total_offset_23[6:0] ? field_byte_23 : _GEN_4539; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4636 = 7'h1a == total_offset_23[6:0] ? field_byte_23 : _GEN_4540; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4637 = 7'h1b == total_offset_23[6:0] ? field_byte_23 : _GEN_4541; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4638 = 7'h1c == total_offset_23[6:0] ? field_byte_23 : _GEN_4542; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4639 = 7'h1d == total_offset_23[6:0] ? field_byte_23 : _GEN_4543; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4640 = 7'h1e == total_offset_23[6:0] ? field_byte_23 : _GEN_4544; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4641 = 7'h1f == total_offset_23[6:0] ? field_byte_23 : _GEN_4545; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4642 = 7'h20 == total_offset_23[6:0] ? field_byte_23 : _GEN_4546; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4643 = 7'h21 == total_offset_23[6:0] ? field_byte_23 : _GEN_4547; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4644 = 7'h22 == total_offset_23[6:0] ? field_byte_23 : _GEN_4548; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4645 = 7'h23 == total_offset_23[6:0] ? field_byte_23 : _GEN_4549; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4646 = 7'h24 == total_offset_23[6:0] ? field_byte_23 : _GEN_4550; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4647 = 7'h25 == total_offset_23[6:0] ? field_byte_23 : _GEN_4551; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4648 = 7'h26 == total_offset_23[6:0] ? field_byte_23 : _GEN_4552; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4649 = 7'h27 == total_offset_23[6:0] ? field_byte_23 : _GEN_4553; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4650 = 7'h28 == total_offset_23[6:0] ? field_byte_23 : _GEN_4554; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4651 = 7'h29 == total_offset_23[6:0] ? field_byte_23 : _GEN_4555; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4652 = 7'h2a == total_offset_23[6:0] ? field_byte_23 : _GEN_4556; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4653 = 7'h2b == total_offset_23[6:0] ? field_byte_23 : _GEN_4557; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4654 = 7'h2c == total_offset_23[6:0] ? field_byte_23 : _GEN_4558; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4655 = 7'h2d == total_offset_23[6:0] ? field_byte_23 : _GEN_4559; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4656 = 7'h2e == total_offset_23[6:0] ? field_byte_23 : _GEN_4560; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4657 = 7'h2f == total_offset_23[6:0] ? field_byte_23 : _GEN_4561; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4658 = 7'h30 == total_offset_23[6:0] ? field_byte_23 : _GEN_4562; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4659 = 7'h31 == total_offset_23[6:0] ? field_byte_23 : _GEN_4563; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4660 = 7'h32 == total_offset_23[6:0] ? field_byte_23 : _GEN_4564; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4661 = 7'h33 == total_offset_23[6:0] ? field_byte_23 : _GEN_4565; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4662 = 7'h34 == total_offset_23[6:0] ? field_byte_23 : _GEN_4566; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4663 = 7'h35 == total_offset_23[6:0] ? field_byte_23 : _GEN_4567; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4664 = 7'h36 == total_offset_23[6:0] ? field_byte_23 : _GEN_4568; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4665 = 7'h37 == total_offset_23[6:0] ? field_byte_23 : _GEN_4569; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4666 = 7'h38 == total_offset_23[6:0] ? field_byte_23 : _GEN_4570; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4667 = 7'h39 == total_offset_23[6:0] ? field_byte_23 : _GEN_4571; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4668 = 7'h3a == total_offset_23[6:0] ? field_byte_23 : _GEN_4572; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4669 = 7'h3b == total_offset_23[6:0] ? field_byte_23 : _GEN_4573; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4670 = 7'h3c == total_offset_23[6:0] ? field_byte_23 : _GEN_4574; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4671 = 7'h3d == total_offset_23[6:0] ? field_byte_23 : _GEN_4575; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4672 = 7'h3e == total_offset_23[6:0] ? field_byte_23 : _GEN_4576; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4673 = 7'h3f == total_offset_23[6:0] ? field_byte_23 : _GEN_4577; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4674 = 7'h40 == total_offset_23[6:0] ? field_byte_23 : _GEN_4578; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4675 = 7'h41 == total_offset_23[6:0] ? field_byte_23 : _GEN_4579; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4676 = 7'h42 == total_offset_23[6:0] ? field_byte_23 : _GEN_4580; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4677 = 7'h43 == total_offset_23[6:0] ? field_byte_23 : _GEN_4581; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4678 = 7'h44 == total_offset_23[6:0] ? field_byte_23 : _GEN_4582; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4679 = 7'h45 == total_offset_23[6:0] ? field_byte_23 : _GEN_4583; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4680 = 7'h46 == total_offset_23[6:0] ? field_byte_23 : _GEN_4584; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4681 = 7'h47 == total_offset_23[6:0] ? field_byte_23 : _GEN_4585; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4682 = 7'h48 == total_offset_23[6:0] ? field_byte_23 : _GEN_4586; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4683 = 7'h49 == total_offset_23[6:0] ? field_byte_23 : _GEN_4587; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4684 = 7'h4a == total_offset_23[6:0] ? field_byte_23 : _GEN_4588; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4685 = 7'h4b == total_offset_23[6:0] ? field_byte_23 : _GEN_4589; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4686 = 7'h4c == total_offset_23[6:0] ? field_byte_23 : _GEN_4590; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4687 = 7'h4d == total_offset_23[6:0] ? field_byte_23 : _GEN_4591; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4688 = 7'h4e == total_offset_23[6:0] ? field_byte_23 : _GEN_4592; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4689 = 7'h4f == total_offset_23[6:0] ? field_byte_23 : _GEN_4593; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4690 = 7'h50 == total_offset_23[6:0] ? field_byte_23 : _GEN_4594; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4691 = 7'h51 == total_offset_23[6:0] ? field_byte_23 : _GEN_4595; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4692 = 7'h52 == total_offset_23[6:0] ? field_byte_23 : _GEN_4596; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4693 = 7'h53 == total_offset_23[6:0] ? field_byte_23 : _GEN_4597; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4694 = 7'h54 == total_offset_23[6:0] ? field_byte_23 : _GEN_4598; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4695 = 7'h55 == total_offset_23[6:0] ? field_byte_23 : _GEN_4599; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4696 = 7'h56 == total_offset_23[6:0] ? field_byte_23 : _GEN_4600; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4697 = 7'h57 == total_offset_23[6:0] ? field_byte_23 : _GEN_4601; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4698 = 7'h58 == total_offset_23[6:0] ? field_byte_23 : _GEN_4602; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4699 = 7'h59 == total_offset_23[6:0] ? field_byte_23 : _GEN_4603; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4700 = 7'h5a == total_offset_23[6:0] ? field_byte_23 : _GEN_4604; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4701 = 7'h5b == total_offset_23[6:0] ? field_byte_23 : _GEN_4605; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4702 = 7'h5c == total_offset_23[6:0] ? field_byte_23 : _GEN_4606; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4703 = 7'h5d == total_offset_23[6:0] ? field_byte_23 : _GEN_4607; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4704 = 7'h5e == total_offset_23[6:0] ? field_byte_23 : _GEN_4608; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4705 = 7'h5f == total_offset_23[6:0] ? field_byte_23 : _GEN_4609; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4706 = 8'h7 < length_2 ? _GEN_4610 : _GEN_4514; // @[executor.scala 290:56]
  wire [7:0] _GEN_4707 = 8'h7 < length_2 ? _GEN_4611 : _GEN_4515; // @[executor.scala 290:56]
  wire [7:0] _GEN_4708 = 8'h7 < length_2 ? _GEN_4612 : _GEN_4516; // @[executor.scala 290:56]
  wire [7:0] _GEN_4709 = 8'h7 < length_2 ? _GEN_4613 : _GEN_4517; // @[executor.scala 290:56]
  wire [7:0] _GEN_4710 = 8'h7 < length_2 ? _GEN_4614 : _GEN_4518; // @[executor.scala 290:56]
  wire [7:0] _GEN_4711 = 8'h7 < length_2 ? _GEN_4615 : _GEN_4519; // @[executor.scala 290:56]
  wire [7:0] _GEN_4712 = 8'h7 < length_2 ? _GEN_4616 : _GEN_4520; // @[executor.scala 290:56]
  wire [7:0] _GEN_4713 = 8'h7 < length_2 ? _GEN_4617 : _GEN_4521; // @[executor.scala 290:56]
  wire [7:0] _GEN_4714 = 8'h7 < length_2 ? _GEN_4618 : _GEN_4522; // @[executor.scala 290:56]
  wire [7:0] _GEN_4715 = 8'h7 < length_2 ? _GEN_4619 : _GEN_4523; // @[executor.scala 290:56]
  wire [7:0] _GEN_4716 = 8'h7 < length_2 ? _GEN_4620 : _GEN_4524; // @[executor.scala 290:56]
  wire [7:0] _GEN_4717 = 8'h7 < length_2 ? _GEN_4621 : _GEN_4525; // @[executor.scala 290:56]
  wire [7:0] _GEN_4718 = 8'h7 < length_2 ? _GEN_4622 : _GEN_4526; // @[executor.scala 290:56]
  wire [7:0] _GEN_4719 = 8'h7 < length_2 ? _GEN_4623 : _GEN_4527; // @[executor.scala 290:56]
  wire [7:0] _GEN_4720 = 8'h7 < length_2 ? _GEN_4624 : _GEN_4528; // @[executor.scala 290:56]
  wire [7:0] _GEN_4721 = 8'h7 < length_2 ? _GEN_4625 : _GEN_4529; // @[executor.scala 290:56]
  wire [7:0] _GEN_4722 = 8'h7 < length_2 ? _GEN_4626 : _GEN_4530; // @[executor.scala 290:56]
  wire [7:0] _GEN_4723 = 8'h7 < length_2 ? _GEN_4627 : _GEN_4531; // @[executor.scala 290:56]
  wire [7:0] _GEN_4724 = 8'h7 < length_2 ? _GEN_4628 : _GEN_4532; // @[executor.scala 290:56]
  wire [7:0] _GEN_4725 = 8'h7 < length_2 ? _GEN_4629 : _GEN_4533; // @[executor.scala 290:56]
  wire [7:0] _GEN_4726 = 8'h7 < length_2 ? _GEN_4630 : _GEN_4534; // @[executor.scala 290:56]
  wire [7:0] _GEN_4727 = 8'h7 < length_2 ? _GEN_4631 : _GEN_4535; // @[executor.scala 290:56]
  wire [7:0] _GEN_4728 = 8'h7 < length_2 ? _GEN_4632 : _GEN_4536; // @[executor.scala 290:56]
  wire [7:0] _GEN_4729 = 8'h7 < length_2 ? _GEN_4633 : _GEN_4537; // @[executor.scala 290:56]
  wire [7:0] _GEN_4730 = 8'h7 < length_2 ? _GEN_4634 : _GEN_4538; // @[executor.scala 290:56]
  wire [7:0] _GEN_4731 = 8'h7 < length_2 ? _GEN_4635 : _GEN_4539; // @[executor.scala 290:56]
  wire [7:0] _GEN_4732 = 8'h7 < length_2 ? _GEN_4636 : _GEN_4540; // @[executor.scala 290:56]
  wire [7:0] _GEN_4733 = 8'h7 < length_2 ? _GEN_4637 : _GEN_4541; // @[executor.scala 290:56]
  wire [7:0] _GEN_4734 = 8'h7 < length_2 ? _GEN_4638 : _GEN_4542; // @[executor.scala 290:56]
  wire [7:0] _GEN_4735 = 8'h7 < length_2 ? _GEN_4639 : _GEN_4543; // @[executor.scala 290:56]
  wire [7:0] _GEN_4736 = 8'h7 < length_2 ? _GEN_4640 : _GEN_4544; // @[executor.scala 290:56]
  wire [7:0] _GEN_4737 = 8'h7 < length_2 ? _GEN_4641 : _GEN_4545; // @[executor.scala 290:56]
  wire [7:0] _GEN_4738 = 8'h7 < length_2 ? _GEN_4642 : _GEN_4546; // @[executor.scala 290:56]
  wire [7:0] _GEN_4739 = 8'h7 < length_2 ? _GEN_4643 : _GEN_4547; // @[executor.scala 290:56]
  wire [7:0] _GEN_4740 = 8'h7 < length_2 ? _GEN_4644 : _GEN_4548; // @[executor.scala 290:56]
  wire [7:0] _GEN_4741 = 8'h7 < length_2 ? _GEN_4645 : _GEN_4549; // @[executor.scala 290:56]
  wire [7:0] _GEN_4742 = 8'h7 < length_2 ? _GEN_4646 : _GEN_4550; // @[executor.scala 290:56]
  wire [7:0] _GEN_4743 = 8'h7 < length_2 ? _GEN_4647 : _GEN_4551; // @[executor.scala 290:56]
  wire [7:0] _GEN_4744 = 8'h7 < length_2 ? _GEN_4648 : _GEN_4552; // @[executor.scala 290:56]
  wire [7:0] _GEN_4745 = 8'h7 < length_2 ? _GEN_4649 : _GEN_4553; // @[executor.scala 290:56]
  wire [7:0] _GEN_4746 = 8'h7 < length_2 ? _GEN_4650 : _GEN_4554; // @[executor.scala 290:56]
  wire [7:0] _GEN_4747 = 8'h7 < length_2 ? _GEN_4651 : _GEN_4555; // @[executor.scala 290:56]
  wire [7:0] _GEN_4748 = 8'h7 < length_2 ? _GEN_4652 : _GEN_4556; // @[executor.scala 290:56]
  wire [7:0] _GEN_4749 = 8'h7 < length_2 ? _GEN_4653 : _GEN_4557; // @[executor.scala 290:56]
  wire [7:0] _GEN_4750 = 8'h7 < length_2 ? _GEN_4654 : _GEN_4558; // @[executor.scala 290:56]
  wire [7:0] _GEN_4751 = 8'h7 < length_2 ? _GEN_4655 : _GEN_4559; // @[executor.scala 290:56]
  wire [7:0] _GEN_4752 = 8'h7 < length_2 ? _GEN_4656 : _GEN_4560; // @[executor.scala 290:56]
  wire [7:0] _GEN_4753 = 8'h7 < length_2 ? _GEN_4657 : _GEN_4561; // @[executor.scala 290:56]
  wire [7:0] _GEN_4754 = 8'h7 < length_2 ? _GEN_4658 : _GEN_4562; // @[executor.scala 290:56]
  wire [7:0] _GEN_4755 = 8'h7 < length_2 ? _GEN_4659 : _GEN_4563; // @[executor.scala 290:56]
  wire [7:0] _GEN_4756 = 8'h7 < length_2 ? _GEN_4660 : _GEN_4564; // @[executor.scala 290:56]
  wire [7:0] _GEN_4757 = 8'h7 < length_2 ? _GEN_4661 : _GEN_4565; // @[executor.scala 290:56]
  wire [7:0] _GEN_4758 = 8'h7 < length_2 ? _GEN_4662 : _GEN_4566; // @[executor.scala 290:56]
  wire [7:0] _GEN_4759 = 8'h7 < length_2 ? _GEN_4663 : _GEN_4567; // @[executor.scala 290:56]
  wire [7:0] _GEN_4760 = 8'h7 < length_2 ? _GEN_4664 : _GEN_4568; // @[executor.scala 290:56]
  wire [7:0] _GEN_4761 = 8'h7 < length_2 ? _GEN_4665 : _GEN_4569; // @[executor.scala 290:56]
  wire [7:0] _GEN_4762 = 8'h7 < length_2 ? _GEN_4666 : _GEN_4570; // @[executor.scala 290:56]
  wire [7:0] _GEN_4763 = 8'h7 < length_2 ? _GEN_4667 : _GEN_4571; // @[executor.scala 290:56]
  wire [7:0] _GEN_4764 = 8'h7 < length_2 ? _GEN_4668 : _GEN_4572; // @[executor.scala 290:56]
  wire [7:0] _GEN_4765 = 8'h7 < length_2 ? _GEN_4669 : _GEN_4573; // @[executor.scala 290:56]
  wire [7:0] _GEN_4766 = 8'h7 < length_2 ? _GEN_4670 : _GEN_4574; // @[executor.scala 290:56]
  wire [7:0] _GEN_4767 = 8'h7 < length_2 ? _GEN_4671 : _GEN_4575; // @[executor.scala 290:56]
  wire [7:0] _GEN_4768 = 8'h7 < length_2 ? _GEN_4672 : _GEN_4576; // @[executor.scala 290:56]
  wire [7:0] _GEN_4769 = 8'h7 < length_2 ? _GEN_4673 : _GEN_4577; // @[executor.scala 290:56]
  wire [7:0] _GEN_4770 = 8'h7 < length_2 ? _GEN_4674 : _GEN_4578; // @[executor.scala 290:56]
  wire [7:0] _GEN_4771 = 8'h7 < length_2 ? _GEN_4675 : _GEN_4579; // @[executor.scala 290:56]
  wire [7:0] _GEN_4772 = 8'h7 < length_2 ? _GEN_4676 : _GEN_4580; // @[executor.scala 290:56]
  wire [7:0] _GEN_4773 = 8'h7 < length_2 ? _GEN_4677 : _GEN_4581; // @[executor.scala 290:56]
  wire [7:0] _GEN_4774 = 8'h7 < length_2 ? _GEN_4678 : _GEN_4582; // @[executor.scala 290:56]
  wire [7:0] _GEN_4775 = 8'h7 < length_2 ? _GEN_4679 : _GEN_4583; // @[executor.scala 290:56]
  wire [7:0] _GEN_4776 = 8'h7 < length_2 ? _GEN_4680 : _GEN_4584; // @[executor.scala 290:56]
  wire [7:0] _GEN_4777 = 8'h7 < length_2 ? _GEN_4681 : _GEN_4585; // @[executor.scala 290:56]
  wire [7:0] _GEN_4778 = 8'h7 < length_2 ? _GEN_4682 : _GEN_4586; // @[executor.scala 290:56]
  wire [7:0] _GEN_4779 = 8'h7 < length_2 ? _GEN_4683 : _GEN_4587; // @[executor.scala 290:56]
  wire [7:0] _GEN_4780 = 8'h7 < length_2 ? _GEN_4684 : _GEN_4588; // @[executor.scala 290:56]
  wire [7:0] _GEN_4781 = 8'h7 < length_2 ? _GEN_4685 : _GEN_4589; // @[executor.scala 290:56]
  wire [7:0] _GEN_4782 = 8'h7 < length_2 ? _GEN_4686 : _GEN_4590; // @[executor.scala 290:56]
  wire [7:0] _GEN_4783 = 8'h7 < length_2 ? _GEN_4687 : _GEN_4591; // @[executor.scala 290:56]
  wire [7:0] _GEN_4784 = 8'h7 < length_2 ? _GEN_4688 : _GEN_4592; // @[executor.scala 290:56]
  wire [7:0] _GEN_4785 = 8'h7 < length_2 ? _GEN_4689 : _GEN_4593; // @[executor.scala 290:56]
  wire [7:0] _GEN_4786 = 8'h7 < length_2 ? _GEN_4690 : _GEN_4594; // @[executor.scala 290:56]
  wire [7:0] _GEN_4787 = 8'h7 < length_2 ? _GEN_4691 : _GEN_4595; // @[executor.scala 290:56]
  wire [7:0] _GEN_4788 = 8'h7 < length_2 ? _GEN_4692 : _GEN_4596; // @[executor.scala 290:56]
  wire [7:0] _GEN_4789 = 8'h7 < length_2 ? _GEN_4693 : _GEN_4597; // @[executor.scala 290:56]
  wire [7:0] _GEN_4790 = 8'h7 < length_2 ? _GEN_4694 : _GEN_4598; // @[executor.scala 290:56]
  wire [7:0] _GEN_4791 = 8'h7 < length_2 ? _GEN_4695 : _GEN_4599; // @[executor.scala 290:56]
  wire [7:0] _GEN_4792 = 8'h7 < length_2 ? _GEN_4696 : _GEN_4600; // @[executor.scala 290:56]
  wire [7:0] _GEN_4793 = 8'h7 < length_2 ? _GEN_4697 : _GEN_4601; // @[executor.scala 290:56]
  wire [7:0] _GEN_4794 = 8'h7 < length_2 ? _GEN_4698 : _GEN_4602; // @[executor.scala 290:56]
  wire [7:0] _GEN_4795 = 8'h7 < length_2 ? _GEN_4699 : _GEN_4603; // @[executor.scala 290:56]
  wire [7:0] _GEN_4796 = 8'h7 < length_2 ? _GEN_4700 : _GEN_4604; // @[executor.scala 290:56]
  wire [7:0] _GEN_4797 = 8'h7 < length_2 ? _GEN_4701 : _GEN_4605; // @[executor.scala 290:56]
  wire [7:0] _GEN_4798 = 8'h7 < length_2 ? _GEN_4702 : _GEN_4606; // @[executor.scala 290:56]
  wire [7:0] _GEN_4799 = 8'h7 < length_2 ? _GEN_4703 : _GEN_4607; // @[executor.scala 290:56]
  wire [7:0] _GEN_4800 = 8'h7 < length_2 ? _GEN_4704 : _GEN_4608; // @[executor.scala 290:56]
  wire [7:0] _GEN_4801 = 8'h7 < length_2 ? _GEN_4705 : _GEN_4609; // @[executor.scala 290:56]
  wire [63:0] _GEN_4802 = length_2 == 8'h0 ? field_2 : _GEN_3169; // @[executor.scala 283:67 executor.scala 284:51]
  wire [7:0] _GEN_4803 = length_2 == 8'h0 ? _GEN_3170 : _GEN_4706; // @[executor.scala 283:67]
  wire [7:0] _GEN_4804 = length_2 == 8'h0 ? _GEN_3171 : _GEN_4707; // @[executor.scala 283:67]
  wire [7:0] _GEN_4805 = length_2 == 8'h0 ? _GEN_3172 : _GEN_4708; // @[executor.scala 283:67]
  wire [7:0] _GEN_4806 = length_2 == 8'h0 ? _GEN_3173 : _GEN_4709; // @[executor.scala 283:67]
  wire [7:0] _GEN_4807 = length_2 == 8'h0 ? _GEN_3174 : _GEN_4710; // @[executor.scala 283:67]
  wire [7:0] _GEN_4808 = length_2 == 8'h0 ? _GEN_3175 : _GEN_4711; // @[executor.scala 283:67]
  wire [7:0] _GEN_4809 = length_2 == 8'h0 ? _GEN_3176 : _GEN_4712; // @[executor.scala 283:67]
  wire [7:0] _GEN_4810 = length_2 == 8'h0 ? _GEN_3177 : _GEN_4713; // @[executor.scala 283:67]
  wire [7:0] _GEN_4811 = length_2 == 8'h0 ? _GEN_3178 : _GEN_4714; // @[executor.scala 283:67]
  wire [7:0] _GEN_4812 = length_2 == 8'h0 ? _GEN_3179 : _GEN_4715; // @[executor.scala 283:67]
  wire [7:0] _GEN_4813 = length_2 == 8'h0 ? _GEN_3180 : _GEN_4716; // @[executor.scala 283:67]
  wire [7:0] _GEN_4814 = length_2 == 8'h0 ? _GEN_3181 : _GEN_4717; // @[executor.scala 283:67]
  wire [7:0] _GEN_4815 = length_2 == 8'h0 ? _GEN_3182 : _GEN_4718; // @[executor.scala 283:67]
  wire [7:0] _GEN_4816 = length_2 == 8'h0 ? _GEN_3183 : _GEN_4719; // @[executor.scala 283:67]
  wire [7:0] _GEN_4817 = length_2 == 8'h0 ? _GEN_3184 : _GEN_4720; // @[executor.scala 283:67]
  wire [7:0] _GEN_4818 = length_2 == 8'h0 ? _GEN_3185 : _GEN_4721; // @[executor.scala 283:67]
  wire [7:0] _GEN_4819 = length_2 == 8'h0 ? _GEN_3186 : _GEN_4722; // @[executor.scala 283:67]
  wire [7:0] _GEN_4820 = length_2 == 8'h0 ? _GEN_3187 : _GEN_4723; // @[executor.scala 283:67]
  wire [7:0] _GEN_4821 = length_2 == 8'h0 ? _GEN_3188 : _GEN_4724; // @[executor.scala 283:67]
  wire [7:0] _GEN_4822 = length_2 == 8'h0 ? _GEN_3189 : _GEN_4725; // @[executor.scala 283:67]
  wire [7:0] _GEN_4823 = length_2 == 8'h0 ? _GEN_3190 : _GEN_4726; // @[executor.scala 283:67]
  wire [7:0] _GEN_4824 = length_2 == 8'h0 ? _GEN_3191 : _GEN_4727; // @[executor.scala 283:67]
  wire [7:0] _GEN_4825 = length_2 == 8'h0 ? _GEN_3192 : _GEN_4728; // @[executor.scala 283:67]
  wire [7:0] _GEN_4826 = length_2 == 8'h0 ? _GEN_3193 : _GEN_4729; // @[executor.scala 283:67]
  wire [7:0] _GEN_4827 = length_2 == 8'h0 ? _GEN_3194 : _GEN_4730; // @[executor.scala 283:67]
  wire [7:0] _GEN_4828 = length_2 == 8'h0 ? _GEN_3195 : _GEN_4731; // @[executor.scala 283:67]
  wire [7:0] _GEN_4829 = length_2 == 8'h0 ? _GEN_3196 : _GEN_4732; // @[executor.scala 283:67]
  wire [7:0] _GEN_4830 = length_2 == 8'h0 ? _GEN_3197 : _GEN_4733; // @[executor.scala 283:67]
  wire [7:0] _GEN_4831 = length_2 == 8'h0 ? _GEN_3198 : _GEN_4734; // @[executor.scala 283:67]
  wire [7:0] _GEN_4832 = length_2 == 8'h0 ? _GEN_3199 : _GEN_4735; // @[executor.scala 283:67]
  wire [7:0] _GEN_4833 = length_2 == 8'h0 ? _GEN_3200 : _GEN_4736; // @[executor.scala 283:67]
  wire [7:0] _GEN_4834 = length_2 == 8'h0 ? _GEN_3201 : _GEN_4737; // @[executor.scala 283:67]
  wire [7:0] _GEN_4835 = length_2 == 8'h0 ? _GEN_3202 : _GEN_4738; // @[executor.scala 283:67]
  wire [7:0] _GEN_4836 = length_2 == 8'h0 ? _GEN_3203 : _GEN_4739; // @[executor.scala 283:67]
  wire [7:0] _GEN_4837 = length_2 == 8'h0 ? _GEN_3204 : _GEN_4740; // @[executor.scala 283:67]
  wire [7:0] _GEN_4838 = length_2 == 8'h0 ? _GEN_3205 : _GEN_4741; // @[executor.scala 283:67]
  wire [7:0] _GEN_4839 = length_2 == 8'h0 ? _GEN_3206 : _GEN_4742; // @[executor.scala 283:67]
  wire [7:0] _GEN_4840 = length_2 == 8'h0 ? _GEN_3207 : _GEN_4743; // @[executor.scala 283:67]
  wire [7:0] _GEN_4841 = length_2 == 8'h0 ? _GEN_3208 : _GEN_4744; // @[executor.scala 283:67]
  wire [7:0] _GEN_4842 = length_2 == 8'h0 ? _GEN_3209 : _GEN_4745; // @[executor.scala 283:67]
  wire [7:0] _GEN_4843 = length_2 == 8'h0 ? _GEN_3210 : _GEN_4746; // @[executor.scala 283:67]
  wire [7:0] _GEN_4844 = length_2 == 8'h0 ? _GEN_3211 : _GEN_4747; // @[executor.scala 283:67]
  wire [7:0] _GEN_4845 = length_2 == 8'h0 ? _GEN_3212 : _GEN_4748; // @[executor.scala 283:67]
  wire [7:0] _GEN_4846 = length_2 == 8'h0 ? _GEN_3213 : _GEN_4749; // @[executor.scala 283:67]
  wire [7:0] _GEN_4847 = length_2 == 8'h0 ? _GEN_3214 : _GEN_4750; // @[executor.scala 283:67]
  wire [7:0] _GEN_4848 = length_2 == 8'h0 ? _GEN_3215 : _GEN_4751; // @[executor.scala 283:67]
  wire [7:0] _GEN_4849 = length_2 == 8'h0 ? _GEN_3216 : _GEN_4752; // @[executor.scala 283:67]
  wire [7:0] _GEN_4850 = length_2 == 8'h0 ? _GEN_3217 : _GEN_4753; // @[executor.scala 283:67]
  wire [7:0] _GEN_4851 = length_2 == 8'h0 ? _GEN_3218 : _GEN_4754; // @[executor.scala 283:67]
  wire [7:0] _GEN_4852 = length_2 == 8'h0 ? _GEN_3219 : _GEN_4755; // @[executor.scala 283:67]
  wire [7:0] _GEN_4853 = length_2 == 8'h0 ? _GEN_3220 : _GEN_4756; // @[executor.scala 283:67]
  wire [7:0] _GEN_4854 = length_2 == 8'h0 ? _GEN_3221 : _GEN_4757; // @[executor.scala 283:67]
  wire [7:0] _GEN_4855 = length_2 == 8'h0 ? _GEN_3222 : _GEN_4758; // @[executor.scala 283:67]
  wire [7:0] _GEN_4856 = length_2 == 8'h0 ? _GEN_3223 : _GEN_4759; // @[executor.scala 283:67]
  wire [7:0] _GEN_4857 = length_2 == 8'h0 ? _GEN_3224 : _GEN_4760; // @[executor.scala 283:67]
  wire [7:0] _GEN_4858 = length_2 == 8'h0 ? _GEN_3225 : _GEN_4761; // @[executor.scala 283:67]
  wire [7:0] _GEN_4859 = length_2 == 8'h0 ? _GEN_3226 : _GEN_4762; // @[executor.scala 283:67]
  wire [7:0] _GEN_4860 = length_2 == 8'h0 ? _GEN_3227 : _GEN_4763; // @[executor.scala 283:67]
  wire [7:0] _GEN_4861 = length_2 == 8'h0 ? _GEN_3228 : _GEN_4764; // @[executor.scala 283:67]
  wire [7:0] _GEN_4862 = length_2 == 8'h0 ? _GEN_3229 : _GEN_4765; // @[executor.scala 283:67]
  wire [7:0] _GEN_4863 = length_2 == 8'h0 ? _GEN_3230 : _GEN_4766; // @[executor.scala 283:67]
  wire [7:0] _GEN_4864 = length_2 == 8'h0 ? _GEN_3231 : _GEN_4767; // @[executor.scala 283:67]
  wire [7:0] _GEN_4865 = length_2 == 8'h0 ? _GEN_3232 : _GEN_4768; // @[executor.scala 283:67]
  wire [7:0] _GEN_4866 = length_2 == 8'h0 ? _GEN_3233 : _GEN_4769; // @[executor.scala 283:67]
  wire [7:0] _GEN_4867 = length_2 == 8'h0 ? _GEN_3234 : _GEN_4770; // @[executor.scala 283:67]
  wire [7:0] _GEN_4868 = length_2 == 8'h0 ? _GEN_3235 : _GEN_4771; // @[executor.scala 283:67]
  wire [7:0] _GEN_4869 = length_2 == 8'h0 ? _GEN_3236 : _GEN_4772; // @[executor.scala 283:67]
  wire [7:0] _GEN_4870 = length_2 == 8'h0 ? _GEN_3237 : _GEN_4773; // @[executor.scala 283:67]
  wire [7:0] _GEN_4871 = length_2 == 8'h0 ? _GEN_3238 : _GEN_4774; // @[executor.scala 283:67]
  wire [7:0] _GEN_4872 = length_2 == 8'h0 ? _GEN_3239 : _GEN_4775; // @[executor.scala 283:67]
  wire [7:0] _GEN_4873 = length_2 == 8'h0 ? _GEN_3240 : _GEN_4776; // @[executor.scala 283:67]
  wire [7:0] _GEN_4874 = length_2 == 8'h0 ? _GEN_3241 : _GEN_4777; // @[executor.scala 283:67]
  wire [7:0] _GEN_4875 = length_2 == 8'h0 ? _GEN_3242 : _GEN_4778; // @[executor.scala 283:67]
  wire [7:0] _GEN_4876 = length_2 == 8'h0 ? _GEN_3243 : _GEN_4779; // @[executor.scala 283:67]
  wire [7:0] _GEN_4877 = length_2 == 8'h0 ? _GEN_3244 : _GEN_4780; // @[executor.scala 283:67]
  wire [7:0] _GEN_4878 = length_2 == 8'h0 ? _GEN_3245 : _GEN_4781; // @[executor.scala 283:67]
  wire [7:0] _GEN_4879 = length_2 == 8'h0 ? _GEN_3246 : _GEN_4782; // @[executor.scala 283:67]
  wire [7:0] _GEN_4880 = length_2 == 8'h0 ? _GEN_3247 : _GEN_4783; // @[executor.scala 283:67]
  wire [7:0] _GEN_4881 = length_2 == 8'h0 ? _GEN_3248 : _GEN_4784; // @[executor.scala 283:67]
  wire [7:0] _GEN_4882 = length_2 == 8'h0 ? _GEN_3249 : _GEN_4785; // @[executor.scala 283:67]
  wire [7:0] _GEN_4883 = length_2 == 8'h0 ? _GEN_3250 : _GEN_4786; // @[executor.scala 283:67]
  wire [7:0] _GEN_4884 = length_2 == 8'h0 ? _GEN_3251 : _GEN_4787; // @[executor.scala 283:67]
  wire [7:0] _GEN_4885 = length_2 == 8'h0 ? _GEN_3252 : _GEN_4788; // @[executor.scala 283:67]
  wire [7:0] _GEN_4886 = length_2 == 8'h0 ? _GEN_3253 : _GEN_4789; // @[executor.scala 283:67]
  wire [7:0] _GEN_4887 = length_2 == 8'h0 ? _GEN_3254 : _GEN_4790; // @[executor.scala 283:67]
  wire [7:0] _GEN_4888 = length_2 == 8'h0 ? _GEN_3255 : _GEN_4791; // @[executor.scala 283:67]
  wire [7:0] _GEN_4889 = length_2 == 8'h0 ? _GEN_3256 : _GEN_4792; // @[executor.scala 283:67]
  wire [7:0] _GEN_4890 = length_2 == 8'h0 ? _GEN_3257 : _GEN_4793; // @[executor.scala 283:67]
  wire [7:0] _GEN_4891 = length_2 == 8'h0 ? _GEN_3258 : _GEN_4794; // @[executor.scala 283:67]
  wire [7:0] _GEN_4892 = length_2 == 8'h0 ? _GEN_3259 : _GEN_4795; // @[executor.scala 283:67]
  wire [7:0] _GEN_4893 = length_2 == 8'h0 ? _GEN_3260 : _GEN_4796; // @[executor.scala 283:67]
  wire [7:0] _GEN_4894 = length_2 == 8'h0 ? _GEN_3261 : _GEN_4797; // @[executor.scala 283:67]
  wire [7:0] _GEN_4895 = length_2 == 8'h0 ? _GEN_3262 : _GEN_4798; // @[executor.scala 283:67]
  wire [7:0] _GEN_4896 = length_2 == 8'h0 ? _GEN_3263 : _GEN_4799; // @[executor.scala 283:67]
  wire [7:0] _GEN_4897 = length_2 == 8'h0 ? _GEN_3264 : _GEN_4800; // @[executor.scala 283:67]
  wire [7:0] _GEN_4898 = length_2 == 8'h0 ? _GEN_3265 : _GEN_4801; // @[executor.scala 283:67]
  wire [7:0] field_byte_24 = field_3[63:56]; // @[executor.scala 287:53]
  wire [8:0] _total_offset_T_24 = {{1'd0}, offset_3}; // @[executor.scala 289:53]
  wire [7:0] total_offset_24 = _total_offset_T_24[7:0]; // @[executor.scala 289:53]
  wire [7:0] _GEN_4899 = 7'h0 == total_offset_24[6:0] ? field_byte_24 : _GEN_4803; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4900 = 7'h1 == total_offset_24[6:0] ? field_byte_24 : _GEN_4804; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4901 = 7'h2 == total_offset_24[6:0] ? field_byte_24 : _GEN_4805; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4902 = 7'h3 == total_offset_24[6:0] ? field_byte_24 : _GEN_4806; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4903 = 7'h4 == total_offset_24[6:0] ? field_byte_24 : _GEN_4807; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4904 = 7'h5 == total_offset_24[6:0] ? field_byte_24 : _GEN_4808; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4905 = 7'h6 == total_offset_24[6:0] ? field_byte_24 : _GEN_4809; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4906 = 7'h7 == total_offset_24[6:0] ? field_byte_24 : _GEN_4810; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4907 = 7'h8 == total_offset_24[6:0] ? field_byte_24 : _GEN_4811; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4908 = 7'h9 == total_offset_24[6:0] ? field_byte_24 : _GEN_4812; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4909 = 7'ha == total_offset_24[6:0] ? field_byte_24 : _GEN_4813; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4910 = 7'hb == total_offset_24[6:0] ? field_byte_24 : _GEN_4814; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4911 = 7'hc == total_offset_24[6:0] ? field_byte_24 : _GEN_4815; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4912 = 7'hd == total_offset_24[6:0] ? field_byte_24 : _GEN_4816; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4913 = 7'he == total_offset_24[6:0] ? field_byte_24 : _GEN_4817; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4914 = 7'hf == total_offset_24[6:0] ? field_byte_24 : _GEN_4818; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4915 = 7'h10 == total_offset_24[6:0] ? field_byte_24 : _GEN_4819; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4916 = 7'h11 == total_offset_24[6:0] ? field_byte_24 : _GEN_4820; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4917 = 7'h12 == total_offset_24[6:0] ? field_byte_24 : _GEN_4821; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4918 = 7'h13 == total_offset_24[6:0] ? field_byte_24 : _GEN_4822; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4919 = 7'h14 == total_offset_24[6:0] ? field_byte_24 : _GEN_4823; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4920 = 7'h15 == total_offset_24[6:0] ? field_byte_24 : _GEN_4824; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4921 = 7'h16 == total_offset_24[6:0] ? field_byte_24 : _GEN_4825; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4922 = 7'h17 == total_offset_24[6:0] ? field_byte_24 : _GEN_4826; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4923 = 7'h18 == total_offset_24[6:0] ? field_byte_24 : _GEN_4827; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4924 = 7'h19 == total_offset_24[6:0] ? field_byte_24 : _GEN_4828; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4925 = 7'h1a == total_offset_24[6:0] ? field_byte_24 : _GEN_4829; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4926 = 7'h1b == total_offset_24[6:0] ? field_byte_24 : _GEN_4830; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4927 = 7'h1c == total_offset_24[6:0] ? field_byte_24 : _GEN_4831; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4928 = 7'h1d == total_offset_24[6:0] ? field_byte_24 : _GEN_4832; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4929 = 7'h1e == total_offset_24[6:0] ? field_byte_24 : _GEN_4833; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4930 = 7'h1f == total_offset_24[6:0] ? field_byte_24 : _GEN_4834; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4931 = 7'h20 == total_offset_24[6:0] ? field_byte_24 : _GEN_4835; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4932 = 7'h21 == total_offset_24[6:0] ? field_byte_24 : _GEN_4836; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4933 = 7'h22 == total_offset_24[6:0] ? field_byte_24 : _GEN_4837; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4934 = 7'h23 == total_offset_24[6:0] ? field_byte_24 : _GEN_4838; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4935 = 7'h24 == total_offset_24[6:0] ? field_byte_24 : _GEN_4839; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4936 = 7'h25 == total_offset_24[6:0] ? field_byte_24 : _GEN_4840; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4937 = 7'h26 == total_offset_24[6:0] ? field_byte_24 : _GEN_4841; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4938 = 7'h27 == total_offset_24[6:0] ? field_byte_24 : _GEN_4842; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4939 = 7'h28 == total_offset_24[6:0] ? field_byte_24 : _GEN_4843; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4940 = 7'h29 == total_offset_24[6:0] ? field_byte_24 : _GEN_4844; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4941 = 7'h2a == total_offset_24[6:0] ? field_byte_24 : _GEN_4845; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4942 = 7'h2b == total_offset_24[6:0] ? field_byte_24 : _GEN_4846; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4943 = 7'h2c == total_offset_24[6:0] ? field_byte_24 : _GEN_4847; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4944 = 7'h2d == total_offset_24[6:0] ? field_byte_24 : _GEN_4848; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4945 = 7'h2e == total_offset_24[6:0] ? field_byte_24 : _GEN_4849; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4946 = 7'h2f == total_offset_24[6:0] ? field_byte_24 : _GEN_4850; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4947 = 7'h30 == total_offset_24[6:0] ? field_byte_24 : _GEN_4851; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4948 = 7'h31 == total_offset_24[6:0] ? field_byte_24 : _GEN_4852; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4949 = 7'h32 == total_offset_24[6:0] ? field_byte_24 : _GEN_4853; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4950 = 7'h33 == total_offset_24[6:0] ? field_byte_24 : _GEN_4854; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4951 = 7'h34 == total_offset_24[6:0] ? field_byte_24 : _GEN_4855; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4952 = 7'h35 == total_offset_24[6:0] ? field_byte_24 : _GEN_4856; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4953 = 7'h36 == total_offset_24[6:0] ? field_byte_24 : _GEN_4857; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4954 = 7'h37 == total_offset_24[6:0] ? field_byte_24 : _GEN_4858; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4955 = 7'h38 == total_offset_24[6:0] ? field_byte_24 : _GEN_4859; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4956 = 7'h39 == total_offset_24[6:0] ? field_byte_24 : _GEN_4860; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4957 = 7'h3a == total_offset_24[6:0] ? field_byte_24 : _GEN_4861; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4958 = 7'h3b == total_offset_24[6:0] ? field_byte_24 : _GEN_4862; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4959 = 7'h3c == total_offset_24[6:0] ? field_byte_24 : _GEN_4863; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4960 = 7'h3d == total_offset_24[6:0] ? field_byte_24 : _GEN_4864; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4961 = 7'h3e == total_offset_24[6:0] ? field_byte_24 : _GEN_4865; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4962 = 7'h3f == total_offset_24[6:0] ? field_byte_24 : _GEN_4866; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4963 = 7'h40 == total_offset_24[6:0] ? field_byte_24 : _GEN_4867; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4964 = 7'h41 == total_offset_24[6:0] ? field_byte_24 : _GEN_4868; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4965 = 7'h42 == total_offset_24[6:0] ? field_byte_24 : _GEN_4869; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4966 = 7'h43 == total_offset_24[6:0] ? field_byte_24 : _GEN_4870; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4967 = 7'h44 == total_offset_24[6:0] ? field_byte_24 : _GEN_4871; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4968 = 7'h45 == total_offset_24[6:0] ? field_byte_24 : _GEN_4872; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4969 = 7'h46 == total_offset_24[6:0] ? field_byte_24 : _GEN_4873; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4970 = 7'h47 == total_offset_24[6:0] ? field_byte_24 : _GEN_4874; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4971 = 7'h48 == total_offset_24[6:0] ? field_byte_24 : _GEN_4875; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4972 = 7'h49 == total_offset_24[6:0] ? field_byte_24 : _GEN_4876; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4973 = 7'h4a == total_offset_24[6:0] ? field_byte_24 : _GEN_4877; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4974 = 7'h4b == total_offset_24[6:0] ? field_byte_24 : _GEN_4878; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4975 = 7'h4c == total_offset_24[6:0] ? field_byte_24 : _GEN_4879; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4976 = 7'h4d == total_offset_24[6:0] ? field_byte_24 : _GEN_4880; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4977 = 7'h4e == total_offset_24[6:0] ? field_byte_24 : _GEN_4881; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4978 = 7'h4f == total_offset_24[6:0] ? field_byte_24 : _GEN_4882; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4979 = 7'h50 == total_offset_24[6:0] ? field_byte_24 : _GEN_4883; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4980 = 7'h51 == total_offset_24[6:0] ? field_byte_24 : _GEN_4884; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4981 = 7'h52 == total_offset_24[6:0] ? field_byte_24 : _GEN_4885; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4982 = 7'h53 == total_offset_24[6:0] ? field_byte_24 : _GEN_4886; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4983 = 7'h54 == total_offset_24[6:0] ? field_byte_24 : _GEN_4887; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4984 = 7'h55 == total_offset_24[6:0] ? field_byte_24 : _GEN_4888; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4985 = 7'h56 == total_offset_24[6:0] ? field_byte_24 : _GEN_4889; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4986 = 7'h57 == total_offset_24[6:0] ? field_byte_24 : _GEN_4890; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4987 = 7'h58 == total_offset_24[6:0] ? field_byte_24 : _GEN_4891; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4988 = 7'h59 == total_offset_24[6:0] ? field_byte_24 : _GEN_4892; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4989 = 7'h5a == total_offset_24[6:0] ? field_byte_24 : _GEN_4893; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4990 = 7'h5b == total_offset_24[6:0] ? field_byte_24 : _GEN_4894; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4991 = 7'h5c == total_offset_24[6:0] ? field_byte_24 : _GEN_4895; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4992 = 7'h5d == total_offset_24[6:0] ? field_byte_24 : _GEN_4896; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4993 = 7'h5e == total_offset_24[6:0] ? field_byte_24 : _GEN_4897; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4994 = 7'h5f == total_offset_24[6:0] ? field_byte_24 : _GEN_4898; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_4995 = 8'h0 < length_3 ? _GEN_4899 : _GEN_4803; // @[executor.scala 290:56]
  wire [7:0] _GEN_4996 = 8'h0 < length_3 ? _GEN_4900 : _GEN_4804; // @[executor.scala 290:56]
  wire [7:0] _GEN_4997 = 8'h0 < length_3 ? _GEN_4901 : _GEN_4805; // @[executor.scala 290:56]
  wire [7:0] _GEN_4998 = 8'h0 < length_3 ? _GEN_4902 : _GEN_4806; // @[executor.scala 290:56]
  wire [7:0] _GEN_4999 = 8'h0 < length_3 ? _GEN_4903 : _GEN_4807; // @[executor.scala 290:56]
  wire [7:0] _GEN_5000 = 8'h0 < length_3 ? _GEN_4904 : _GEN_4808; // @[executor.scala 290:56]
  wire [7:0] _GEN_5001 = 8'h0 < length_3 ? _GEN_4905 : _GEN_4809; // @[executor.scala 290:56]
  wire [7:0] _GEN_5002 = 8'h0 < length_3 ? _GEN_4906 : _GEN_4810; // @[executor.scala 290:56]
  wire [7:0] _GEN_5003 = 8'h0 < length_3 ? _GEN_4907 : _GEN_4811; // @[executor.scala 290:56]
  wire [7:0] _GEN_5004 = 8'h0 < length_3 ? _GEN_4908 : _GEN_4812; // @[executor.scala 290:56]
  wire [7:0] _GEN_5005 = 8'h0 < length_3 ? _GEN_4909 : _GEN_4813; // @[executor.scala 290:56]
  wire [7:0] _GEN_5006 = 8'h0 < length_3 ? _GEN_4910 : _GEN_4814; // @[executor.scala 290:56]
  wire [7:0] _GEN_5007 = 8'h0 < length_3 ? _GEN_4911 : _GEN_4815; // @[executor.scala 290:56]
  wire [7:0] _GEN_5008 = 8'h0 < length_3 ? _GEN_4912 : _GEN_4816; // @[executor.scala 290:56]
  wire [7:0] _GEN_5009 = 8'h0 < length_3 ? _GEN_4913 : _GEN_4817; // @[executor.scala 290:56]
  wire [7:0] _GEN_5010 = 8'h0 < length_3 ? _GEN_4914 : _GEN_4818; // @[executor.scala 290:56]
  wire [7:0] _GEN_5011 = 8'h0 < length_3 ? _GEN_4915 : _GEN_4819; // @[executor.scala 290:56]
  wire [7:0] _GEN_5012 = 8'h0 < length_3 ? _GEN_4916 : _GEN_4820; // @[executor.scala 290:56]
  wire [7:0] _GEN_5013 = 8'h0 < length_3 ? _GEN_4917 : _GEN_4821; // @[executor.scala 290:56]
  wire [7:0] _GEN_5014 = 8'h0 < length_3 ? _GEN_4918 : _GEN_4822; // @[executor.scala 290:56]
  wire [7:0] _GEN_5015 = 8'h0 < length_3 ? _GEN_4919 : _GEN_4823; // @[executor.scala 290:56]
  wire [7:0] _GEN_5016 = 8'h0 < length_3 ? _GEN_4920 : _GEN_4824; // @[executor.scala 290:56]
  wire [7:0] _GEN_5017 = 8'h0 < length_3 ? _GEN_4921 : _GEN_4825; // @[executor.scala 290:56]
  wire [7:0] _GEN_5018 = 8'h0 < length_3 ? _GEN_4922 : _GEN_4826; // @[executor.scala 290:56]
  wire [7:0] _GEN_5019 = 8'h0 < length_3 ? _GEN_4923 : _GEN_4827; // @[executor.scala 290:56]
  wire [7:0] _GEN_5020 = 8'h0 < length_3 ? _GEN_4924 : _GEN_4828; // @[executor.scala 290:56]
  wire [7:0] _GEN_5021 = 8'h0 < length_3 ? _GEN_4925 : _GEN_4829; // @[executor.scala 290:56]
  wire [7:0] _GEN_5022 = 8'h0 < length_3 ? _GEN_4926 : _GEN_4830; // @[executor.scala 290:56]
  wire [7:0] _GEN_5023 = 8'h0 < length_3 ? _GEN_4927 : _GEN_4831; // @[executor.scala 290:56]
  wire [7:0] _GEN_5024 = 8'h0 < length_3 ? _GEN_4928 : _GEN_4832; // @[executor.scala 290:56]
  wire [7:0] _GEN_5025 = 8'h0 < length_3 ? _GEN_4929 : _GEN_4833; // @[executor.scala 290:56]
  wire [7:0] _GEN_5026 = 8'h0 < length_3 ? _GEN_4930 : _GEN_4834; // @[executor.scala 290:56]
  wire [7:0] _GEN_5027 = 8'h0 < length_3 ? _GEN_4931 : _GEN_4835; // @[executor.scala 290:56]
  wire [7:0] _GEN_5028 = 8'h0 < length_3 ? _GEN_4932 : _GEN_4836; // @[executor.scala 290:56]
  wire [7:0] _GEN_5029 = 8'h0 < length_3 ? _GEN_4933 : _GEN_4837; // @[executor.scala 290:56]
  wire [7:0] _GEN_5030 = 8'h0 < length_3 ? _GEN_4934 : _GEN_4838; // @[executor.scala 290:56]
  wire [7:0] _GEN_5031 = 8'h0 < length_3 ? _GEN_4935 : _GEN_4839; // @[executor.scala 290:56]
  wire [7:0] _GEN_5032 = 8'h0 < length_3 ? _GEN_4936 : _GEN_4840; // @[executor.scala 290:56]
  wire [7:0] _GEN_5033 = 8'h0 < length_3 ? _GEN_4937 : _GEN_4841; // @[executor.scala 290:56]
  wire [7:0] _GEN_5034 = 8'h0 < length_3 ? _GEN_4938 : _GEN_4842; // @[executor.scala 290:56]
  wire [7:0] _GEN_5035 = 8'h0 < length_3 ? _GEN_4939 : _GEN_4843; // @[executor.scala 290:56]
  wire [7:0] _GEN_5036 = 8'h0 < length_3 ? _GEN_4940 : _GEN_4844; // @[executor.scala 290:56]
  wire [7:0] _GEN_5037 = 8'h0 < length_3 ? _GEN_4941 : _GEN_4845; // @[executor.scala 290:56]
  wire [7:0] _GEN_5038 = 8'h0 < length_3 ? _GEN_4942 : _GEN_4846; // @[executor.scala 290:56]
  wire [7:0] _GEN_5039 = 8'h0 < length_3 ? _GEN_4943 : _GEN_4847; // @[executor.scala 290:56]
  wire [7:0] _GEN_5040 = 8'h0 < length_3 ? _GEN_4944 : _GEN_4848; // @[executor.scala 290:56]
  wire [7:0] _GEN_5041 = 8'h0 < length_3 ? _GEN_4945 : _GEN_4849; // @[executor.scala 290:56]
  wire [7:0] _GEN_5042 = 8'h0 < length_3 ? _GEN_4946 : _GEN_4850; // @[executor.scala 290:56]
  wire [7:0] _GEN_5043 = 8'h0 < length_3 ? _GEN_4947 : _GEN_4851; // @[executor.scala 290:56]
  wire [7:0] _GEN_5044 = 8'h0 < length_3 ? _GEN_4948 : _GEN_4852; // @[executor.scala 290:56]
  wire [7:0] _GEN_5045 = 8'h0 < length_3 ? _GEN_4949 : _GEN_4853; // @[executor.scala 290:56]
  wire [7:0] _GEN_5046 = 8'h0 < length_3 ? _GEN_4950 : _GEN_4854; // @[executor.scala 290:56]
  wire [7:0] _GEN_5047 = 8'h0 < length_3 ? _GEN_4951 : _GEN_4855; // @[executor.scala 290:56]
  wire [7:0] _GEN_5048 = 8'h0 < length_3 ? _GEN_4952 : _GEN_4856; // @[executor.scala 290:56]
  wire [7:0] _GEN_5049 = 8'h0 < length_3 ? _GEN_4953 : _GEN_4857; // @[executor.scala 290:56]
  wire [7:0] _GEN_5050 = 8'h0 < length_3 ? _GEN_4954 : _GEN_4858; // @[executor.scala 290:56]
  wire [7:0] _GEN_5051 = 8'h0 < length_3 ? _GEN_4955 : _GEN_4859; // @[executor.scala 290:56]
  wire [7:0] _GEN_5052 = 8'h0 < length_3 ? _GEN_4956 : _GEN_4860; // @[executor.scala 290:56]
  wire [7:0] _GEN_5053 = 8'h0 < length_3 ? _GEN_4957 : _GEN_4861; // @[executor.scala 290:56]
  wire [7:0] _GEN_5054 = 8'h0 < length_3 ? _GEN_4958 : _GEN_4862; // @[executor.scala 290:56]
  wire [7:0] _GEN_5055 = 8'h0 < length_3 ? _GEN_4959 : _GEN_4863; // @[executor.scala 290:56]
  wire [7:0] _GEN_5056 = 8'h0 < length_3 ? _GEN_4960 : _GEN_4864; // @[executor.scala 290:56]
  wire [7:0] _GEN_5057 = 8'h0 < length_3 ? _GEN_4961 : _GEN_4865; // @[executor.scala 290:56]
  wire [7:0] _GEN_5058 = 8'h0 < length_3 ? _GEN_4962 : _GEN_4866; // @[executor.scala 290:56]
  wire [7:0] _GEN_5059 = 8'h0 < length_3 ? _GEN_4963 : _GEN_4867; // @[executor.scala 290:56]
  wire [7:0] _GEN_5060 = 8'h0 < length_3 ? _GEN_4964 : _GEN_4868; // @[executor.scala 290:56]
  wire [7:0] _GEN_5061 = 8'h0 < length_3 ? _GEN_4965 : _GEN_4869; // @[executor.scala 290:56]
  wire [7:0] _GEN_5062 = 8'h0 < length_3 ? _GEN_4966 : _GEN_4870; // @[executor.scala 290:56]
  wire [7:0] _GEN_5063 = 8'h0 < length_3 ? _GEN_4967 : _GEN_4871; // @[executor.scala 290:56]
  wire [7:0] _GEN_5064 = 8'h0 < length_3 ? _GEN_4968 : _GEN_4872; // @[executor.scala 290:56]
  wire [7:0] _GEN_5065 = 8'h0 < length_3 ? _GEN_4969 : _GEN_4873; // @[executor.scala 290:56]
  wire [7:0] _GEN_5066 = 8'h0 < length_3 ? _GEN_4970 : _GEN_4874; // @[executor.scala 290:56]
  wire [7:0] _GEN_5067 = 8'h0 < length_3 ? _GEN_4971 : _GEN_4875; // @[executor.scala 290:56]
  wire [7:0] _GEN_5068 = 8'h0 < length_3 ? _GEN_4972 : _GEN_4876; // @[executor.scala 290:56]
  wire [7:0] _GEN_5069 = 8'h0 < length_3 ? _GEN_4973 : _GEN_4877; // @[executor.scala 290:56]
  wire [7:0] _GEN_5070 = 8'h0 < length_3 ? _GEN_4974 : _GEN_4878; // @[executor.scala 290:56]
  wire [7:0] _GEN_5071 = 8'h0 < length_3 ? _GEN_4975 : _GEN_4879; // @[executor.scala 290:56]
  wire [7:0] _GEN_5072 = 8'h0 < length_3 ? _GEN_4976 : _GEN_4880; // @[executor.scala 290:56]
  wire [7:0] _GEN_5073 = 8'h0 < length_3 ? _GEN_4977 : _GEN_4881; // @[executor.scala 290:56]
  wire [7:0] _GEN_5074 = 8'h0 < length_3 ? _GEN_4978 : _GEN_4882; // @[executor.scala 290:56]
  wire [7:0] _GEN_5075 = 8'h0 < length_3 ? _GEN_4979 : _GEN_4883; // @[executor.scala 290:56]
  wire [7:0] _GEN_5076 = 8'h0 < length_3 ? _GEN_4980 : _GEN_4884; // @[executor.scala 290:56]
  wire [7:0] _GEN_5077 = 8'h0 < length_3 ? _GEN_4981 : _GEN_4885; // @[executor.scala 290:56]
  wire [7:0] _GEN_5078 = 8'h0 < length_3 ? _GEN_4982 : _GEN_4886; // @[executor.scala 290:56]
  wire [7:0] _GEN_5079 = 8'h0 < length_3 ? _GEN_4983 : _GEN_4887; // @[executor.scala 290:56]
  wire [7:0] _GEN_5080 = 8'h0 < length_3 ? _GEN_4984 : _GEN_4888; // @[executor.scala 290:56]
  wire [7:0] _GEN_5081 = 8'h0 < length_3 ? _GEN_4985 : _GEN_4889; // @[executor.scala 290:56]
  wire [7:0] _GEN_5082 = 8'h0 < length_3 ? _GEN_4986 : _GEN_4890; // @[executor.scala 290:56]
  wire [7:0] _GEN_5083 = 8'h0 < length_3 ? _GEN_4987 : _GEN_4891; // @[executor.scala 290:56]
  wire [7:0] _GEN_5084 = 8'h0 < length_3 ? _GEN_4988 : _GEN_4892; // @[executor.scala 290:56]
  wire [7:0] _GEN_5085 = 8'h0 < length_3 ? _GEN_4989 : _GEN_4893; // @[executor.scala 290:56]
  wire [7:0] _GEN_5086 = 8'h0 < length_3 ? _GEN_4990 : _GEN_4894; // @[executor.scala 290:56]
  wire [7:0] _GEN_5087 = 8'h0 < length_3 ? _GEN_4991 : _GEN_4895; // @[executor.scala 290:56]
  wire [7:0] _GEN_5088 = 8'h0 < length_3 ? _GEN_4992 : _GEN_4896; // @[executor.scala 290:56]
  wire [7:0] _GEN_5089 = 8'h0 < length_3 ? _GEN_4993 : _GEN_4897; // @[executor.scala 290:56]
  wire [7:0] _GEN_5090 = 8'h0 < length_3 ? _GEN_4994 : _GEN_4898; // @[executor.scala 290:56]
  wire [7:0] field_byte_25 = field_3[55:48]; // @[executor.scala 287:53]
  wire [7:0] total_offset_25 = offset_3 + 8'h1; // @[executor.scala 289:53]
  wire [7:0] _GEN_5091 = 7'h0 == total_offset_25[6:0] ? field_byte_25 : _GEN_4995; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5092 = 7'h1 == total_offset_25[6:0] ? field_byte_25 : _GEN_4996; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5093 = 7'h2 == total_offset_25[6:0] ? field_byte_25 : _GEN_4997; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5094 = 7'h3 == total_offset_25[6:0] ? field_byte_25 : _GEN_4998; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5095 = 7'h4 == total_offset_25[6:0] ? field_byte_25 : _GEN_4999; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5096 = 7'h5 == total_offset_25[6:0] ? field_byte_25 : _GEN_5000; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5097 = 7'h6 == total_offset_25[6:0] ? field_byte_25 : _GEN_5001; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5098 = 7'h7 == total_offset_25[6:0] ? field_byte_25 : _GEN_5002; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5099 = 7'h8 == total_offset_25[6:0] ? field_byte_25 : _GEN_5003; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5100 = 7'h9 == total_offset_25[6:0] ? field_byte_25 : _GEN_5004; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5101 = 7'ha == total_offset_25[6:0] ? field_byte_25 : _GEN_5005; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5102 = 7'hb == total_offset_25[6:0] ? field_byte_25 : _GEN_5006; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5103 = 7'hc == total_offset_25[6:0] ? field_byte_25 : _GEN_5007; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5104 = 7'hd == total_offset_25[6:0] ? field_byte_25 : _GEN_5008; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5105 = 7'he == total_offset_25[6:0] ? field_byte_25 : _GEN_5009; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5106 = 7'hf == total_offset_25[6:0] ? field_byte_25 : _GEN_5010; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5107 = 7'h10 == total_offset_25[6:0] ? field_byte_25 : _GEN_5011; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5108 = 7'h11 == total_offset_25[6:0] ? field_byte_25 : _GEN_5012; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5109 = 7'h12 == total_offset_25[6:0] ? field_byte_25 : _GEN_5013; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5110 = 7'h13 == total_offset_25[6:0] ? field_byte_25 : _GEN_5014; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5111 = 7'h14 == total_offset_25[6:0] ? field_byte_25 : _GEN_5015; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5112 = 7'h15 == total_offset_25[6:0] ? field_byte_25 : _GEN_5016; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5113 = 7'h16 == total_offset_25[6:0] ? field_byte_25 : _GEN_5017; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5114 = 7'h17 == total_offset_25[6:0] ? field_byte_25 : _GEN_5018; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5115 = 7'h18 == total_offset_25[6:0] ? field_byte_25 : _GEN_5019; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5116 = 7'h19 == total_offset_25[6:0] ? field_byte_25 : _GEN_5020; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5117 = 7'h1a == total_offset_25[6:0] ? field_byte_25 : _GEN_5021; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5118 = 7'h1b == total_offset_25[6:0] ? field_byte_25 : _GEN_5022; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5119 = 7'h1c == total_offset_25[6:0] ? field_byte_25 : _GEN_5023; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5120 = 7'h1d == total_offset_25[6:0] ? field_byte_25 : _GEN_5024; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5121 = 7'h1e == total_offset_25[6:0] ? field_byte_25 : _GEN_5025; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5122 = 7'h1f == total_offset_25[6:0] ? field_byte_25 : _GEN_5026; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5123 = 7'h20 == total_offset_25[6:0] ? field_byte_25 : _GEN_5027; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5124 = 7'h21 == total_offset_25[6:0] ? field_byte_25 : _GEN_5028; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5125 = 7'h22 == total_offset_25[6:0] ? field_byte_25 : _GEN_5029; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5126 = 7'h23 == total_offset_25[6:0] ? field_byte_25 : _GEN_5030; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5127 = 7'h24 == total_offset_25[6:0] ? field_byte_25 : _GEN_5031; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5128 = 7'h25 == total_offset_25[6:0] ? field_byte_25 : _GEN_5032; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5129 = 7'h26 == total_offset_25[6:0] ? field_byte_25 : _GEN_5033; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5130 = 7'h27 == total_offset_25[6:0] ? field_byte_25 : _GEN_5034; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5131 = 7'h28 == total_offset_25[6:0] ? field_byte_25 : _GEN_5035; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5132 = 7'h29 == total_offset_25[6:0] ? field_byte_25 : _GEN_5036; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5133 = 7'h2a == total_offset_25[6:0] ? field_byte_25 : _GEN_5037; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5134 = 7'h2b == total_offset_25[6:0] ? field_byte_25 : _GEN_5038; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5135 = 7'h2c == total_offset_25[6:0] ? field_byte_25 : _GEN_5039; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5136 = 7'h2d == total_offset_25[6:0] ? field_byte_25 : _GEN_5040; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5137 = 7'h2e == total_offset_25[6:0] ? field_byte_25 : _GEN_5041; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5138 = 7'h2f == total_offset_25[6:0] ? field_byte_25 : _GEN_5042; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5139 = 7'h30 == total_offset_25[6:0] ? field_byte_25 : _GEN_5043; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5140 = 7'h31 == total_offset_25[6:0] ? field_byte_25 : _GEN_5044; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5141 = 7'h32 == total_offset_25[6:0] ? field_byte_25 : _GEN_5045; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5142 = 7'h33 == total_offset_25[6:0] ? field_byte_25 : _GEN_5046; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5143 = 7'h34 == total_offset_25[6:0] ? field_byte_25 : _GEN_5047; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5144 = 7'h35 == total_offset_25[6:0] ? field_byte_25 : _GEN_5048; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5145 = 7'h36 == total_offset_25[6:0] ? field_byte_25 : _GEN_5049; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5146 = 7'h37 == total_offset_25[6:0] ? field_byte_25 : _GEN_5050; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5147 = 7'h38 == total_offset_25[6:0] ? field_byte_25 : _GEN_5051; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5148 = 7'h39 == total_offset_25[6:0] ? field_byte_25 : _GEN_5052; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5149 = 7'h3a == total_offset_25[6:0] ? field_byte_25 : _GEN_5053; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5150 = 7'h3b == total_offset_25[6:0] ? field_byte_25 : _GEN_5054; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5151 = 7'h3c == total_offset_25[6:0] ? field_byte_25 : _GEN_5055; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5152 = 7'h3d == total_offset_25[6:0] ? field_byte_25 : _GEN_5056; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5153 = 7'h3e == total_offset_25[6:0] ? field_byte_25 : _GEN_5057; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5154 = 7'h3f == total_offset_25[6:0] ? field_byte_25 : _GEN_5058; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5155 = 7'h40 == total_offset_25[6:0] ? field_byte_25 : _GEN_5059; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5156 = 7'h41 == total_offset_25[6:0] ? field_byte_25 : _GEN_5060; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5157 = 7'h42 == total_offset_25[6:0] ? field_byte_25 : _GEN_5061; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5158 = 7'h43 == total_offset_25[6:0] ? field_byte_25 : _GEN_5062; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5159 = 7'h44 == total_offset_25[6:0] ? field_byte_25 : _GEN_5063; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5160 = 7'h45 == total_offset_25[6:0] ? field_byte_25 : _GEN_5064; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5161 = 7'h46 == total_offset_25[6:0] ? field_byte_25 : _GEN_5065; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5162 = 7'h47 == total_offset_25[6:0] ? field_byte_25 : _GEN_5066; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5163 = 7'h48 == total_offset_25[6:0] ? field_byte_25 : _GEN_5067; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5164 = 7'h49 == total_offset_25[6:0] ? field_byte_25 : _GEN_5068; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5165 = 7'h4a == total_offset_25[6:0] ? field_byte_25 : _GEN_5069; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5166 = 7'h4b == total_offset_25[6:0] ? field_byte_25 : _GEN_5070; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5167 = 7'h4c == total_offset_25[6:0] ? field_byte_25 : _GEN_5071; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5168 = 7'h4d == total_offset_25[6:0] ? field_byte_25 : _GEN_5072; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5169 = 7'h4e == total_offset_25[6:0] ? field_byte_25 : _GEN_5073; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5170 = 7'h4f == total_offset_25[6:0] ? field_byte_25 : _GEN_5074; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5171 = 7'h50 == total_offset_25[6:0] ? field_byte_25 : _GEN_5075; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5172 = 7'h51 == total_offset_25[6:0] ? field_byte_25 : _GEN_5076; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5173 = 7'h52 == total_offset_25[6:0] ? field_byte_25 : _GEN_5077; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5174 = 7'h53 == total_offset_25[6:0] ? field_byte_25 : _GEN_5078; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5175 = 7'h54 == total_offset_25[6:0] ? field_byte_25 : _GEN_5079; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5176 = 7'h55 == total_offset_25[6:0] ? field_byte_25 : _GEN_5080; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5177 = 7'h56 == total_offset_25[6:0] ? field_byte_25 : _GEN_5081; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5178 = 7'h57 == total_offset_25[6:0] ? field_byte_25 : _GEN_5082; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5179 = 7'h58 == total_offset_25[6:0] ? field_byte_25 : _GEN_5083; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5180 = 7'h59 == total_offset_25[6:0] ? field_byte_25 : _GEN_5084; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5181 = 7'h5a == total_offset_25[6:0] ? field_byte_25 : _GEN_5085; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5182 = 7'h5b == total_offset_25[6:0] ? field_byte_25 : _GEN_5086; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5183 = 7'h5c == total_offset_25[6:0] ? field_byte_25 : _GEN_5087; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5184 = 7'h5d == total_offset_25[6:0] ? field_byte_25 : _GEN_5088; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5185 = 7'h5e == total_offset_25[6:0] ? field_byte_25 : _GEN_5089; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5186 = 7'h5f == total_offset_25[6:0] ? field_byte_25 : _GEN_5090; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5187 = 8'h1 < length_3 ? _GEN_5091 : _GEN_4995; // @[executor.scala 290:56]
  wire [7:0] _GEN_5188 = 8'h1 < length_3 ? _GEN_5092 : _GEN_4996; // @[executor.scala 290:56]
  wire [7:0] _GEN_5189 = 8'h1 < length_3 ? _GEN_5093 : _GEN_4997; // @[executor.scala 290:56]
  wire [7:0] _GEN_5190 = 8'h1 < length_3 ? _GEN_5094 : _GEN_4998; // @[executor.scala 290:56]
  wire [7:0] _GEN_5191 = 8'h1 < length_3 ? _GEN_5095 : _GEN_4999; // @[executor.scala 290:56]
  wire [7:0] _GEN_5192 = 8'h1 < length_3 ? _GEN_5096 : _GEN_5000; // @[executor.scala 290:56]
  wire [7:0] _GEN_5193 = 8'h1 < length_3 ? _GEN_5097 : _GEN_5001; // @[executor.scala 290:56]
  wire [7:0] _GEN_5194 = 8'h1 < length_3 ? _GEN_5098 : _GEN_5002; // @[executor.scala 290:56]
  wire [7:0] _GEN_5195 = 8'h1 < length_3 ? _GEN_5099 : _GEN_5003; // @[executor.scala 290:56]
  wire [7:0] _GEN_5196 = 8'h1 < length_3 ? _GEN_5100 : _GEN_5004; // @[executor.scala 290:56]
  wire [7:0] _GEN_5197 = 8'h1 < length_3 ? _GEN_5101 : _GEN_5005; // @[executor.scala 290:56]
  wire [7:0] _GEN_5198 = 8'h1 < length_3 ? _GEN_5102 : _GEN_5006; // @[executor.scala 290:56]
  wire [7:0] _GEN_5199 = 8'h1 < length_3 ? _GEN_5103 : _GEN_5007; // @[executor.scala 290:56]
  wire [7:0] _GEN_5200 = 8'h1 < length_3 ? _GEN_5104 : _GEN_5008; // @[executor.scala 290:56]
  wire [7:0] _GEN_5201 = 8'h1 < length_3 ? _GEN_5105 : _GEN_5009; // @[executor.scala 290:56]
  wire [7:0] _GEN_5202 = 8'h1 < length_3 ? _GEN_5106 : _GEN_5010; // @[executor.scala 290:56]
  wire [7:0] _GEN_5203 = 8'h1 < length_3 ? _GEN_5107 : _GEN_5011; // @[executor.scala 290:56]
  wire [7:0] _GEN_5204 = 8'h1 < length_3 ? _GEN_5108 : _GEN_5012; // @[executor.scala 290:56]
  wire [7:0] _GEN_5205 = 8'h1 < length_3 ? _GEN_5109 : _GEN_5013; // @[executor.scala 290:56]
  wire [7:0] _GEN_5206 = 8'h1 < length_3 ? _GEN_5110 : _GEN_5014; // @[executor.scala 290:56]
  wire [7:0] _GEN_5207 = 8'h1 < length_3 ? _GEN_5111 : _GEN_5015; // @[executor.scala 290:56]
  wire [7:0] _GEN_5208 = 8'h1 < length_3 ? _GEN_5112 : _GEN_5016; // @[executor.scala 290:56]
  wire [7:0] _GEN_5209 = 8'h1 < length_3 ? _GEN_5113 : _GEN_5017; // @[executor.scala 290:56]
  wire [7:0] _GEN_5210 = 8'h1 < length_3 ? _GEN_5114 : _GEN_5018; // @[executor.scala 290:56]
  wire [7:0] _GEN_5211 = 8'h1 < length_3 ? _GEN_5115 : _GEN_5019; // @[executor.scala 290:56]
  wire [7:0] _GEN_5212 = 8'h1 < length_3 ? _GEN_5116 : _GEN_5020; // @[executor.scala 290:56]
  wire [7:0] _GEN_5213 = 8'h1 < length_3 ? _GEN_5117 : _GEN_5021; // @[executor.scala 290:56]
  wire [7:0] _GEN_5214 = 8'h1 < length_3 ? _GEN_5118 : _GEN_5022; // @[executor.scala 290:56]
  wire [7:0] _GEN_5215 = 8'h1 < length_3 ? _GEN_5119 : _GEN_5023; // @[executor.scala 290:56]
  wire [7:0] _GEN_5216 = 8'h1 < length_3 ? _GEN_5120 : _GEN_5024; // @[executor.scala 290:56]
  wire [7:0] _GEN_5217 = 8'h1 < length_3 ? _GEN_5121 : _GEN_5025; // @[executor.scala 290:56]
  wire [7:0] _GEN_5218 = 8'h1 < length_3 ? _GEN_5122 : _GEN_5026; // @[executor.scala 290:56]
  wire [7:0] _GEN_5219 = 8'h1 < length_3 ? _GEN_5123 : _GEN_5027; // @[executor.scala 290:56]
  wire [7:0] _GEN_5220 = 8'h1 < length_3 ? _GEN_5124 : _GEN_5028; // @[executor.scala 290:56]
  wire [7:0] _GEN_5221 = 8'h1 < length_3 ? _GEN_5125 : _GEN_5029; // @[executor.scala 290:56]
  wire [7:0] _GEN_5222 = 8'h1 < length_3 ? _GEN_5126 : _GEN_5030; // @[executor.scala 290:56]
  wire [7:0] _GEN_5223 = 8'h1 < length_3 ? _GEN_5127 : _GEN_5031; // @[executor.scala 290:56]
  wire [7:0] _GEN_5224 = 8'h1 < length_3 ? _GEN_5128 : _GEN_5032; // @[executor.scala 290:56]
  wire [7:0] _GEN_5225 = 8'h1 < length_3 ? _GEN_5129 : _GEN_5033; // @[executor.scala 290:56]
  wire [7:0] _GEN_5226 = 8'h1 < length_3 ? _GEN_5130 : _GEN_5034; // @[executor.scala 290:56]
  wire [7:0] _GEN_5227 = 8'h1 < length_3 ? _GEN_5131 : _GEN_5035; // @[executor.scala 290:56]
  wire [7:0] _GEN_5228 = 8'h1 < length_3 ? _GEN_5132 : _GEN_5036; // @[executor.scala 290:56]
  wire [7:0] _GEN_5229 = 8'h1 < length_3 ? _GEN_5133 : _GEN_5037; // @[executor.scala 290:56]
  wire [7:0] _GEN_5230 = 8'h1 < length_3 ? _GEN_5134 : _GEN_5038; // @[executor.scala 290:56]
  wire [7:0] _GEN_5231 = 8'h1 < length_3 ? _GEN_5135 : _GEN_5039; // @[executor.scala 290:56]
  wire [7:0] _GEN_5232 = 8'h1 < length_3 ? _GEN_5136 : _GEN_5040; // @[executor.scala 290:56]
  wire [7:0] _GEN_5233 = 8'h1 < length_3 ? _GEN_5137 : _GEN_5041; // @[executor.scala 290:56]
  wire [7:0] _GEN_5234 = 8'h1 < length_3 ? _GEN_5138 : _GEN_5042; // @[executor.scala 290:56]
  wire [7:0] _GEN_5235 = 8'h1 < length_3 ? _GEN_5139 : _GEN_5043; // @[executor.scala 290:56]
  wire [7:0] _GEN_5236 = 8'h1 < length_3 ? _GEN_5140 : _GEN_5044; // @[executor.scala 290:56]
  wire [7:0] _GEN_5237 = 8'h1 < length_3 ? _GEN_5141 : _GEN_5045; // @[executor.scala 290:56]
  wire [7:0] _GEN_5238 = 8'h1 < length_3 ? _GEN_5142 : _GEN_5046; // @[executor.scala 290:56]
  wire [7:0] _GEN_5239 = 8'h1 < length_3 ? _GEN_5143 : _GEN_5047; // @[executor.scala 290:56]
  wire [7:0] _GEN_5240 = 8'h1 < length_3 ? _GEN_5144 : _GEN_5048; // @[executor.scala 290:56]
  wire [7:0] _GEN_5241 = 8'h1 < length_3 ? _GEN_5145 : _GEN_5049; // @[executor.scala 290:56]
  wire [7:0] _GEN_5242 = 8'h1 < length_3 ? _GEN_5146 : _GEN_5050; // @[executor.scala 290:56]
  wire [7:0] _GEN_5243 = 8'h1 < length_3 ? _GEN_5147 : _GEN_5051; // @[executor.scala 290:56]
  wire [7:0] _GEN_5244 = 8'h1 < length_3 ? _GEN_5148 : _GEN_5052; // @[executor.scala 290:56]
  wire [7:0] _GEN_5245 = 8'h1 < length_3 ? _GEN_5149 : _GEN_5053; // @[executor.scala 290:56]
  wire [7:0] _GEN_5246 = 8'h1 < length_3 ? _GEN_5150 : _GEN_5054; // @[executor.scala 290:56]
  wire [7:0] _GEN_5247 = 8'h1 < length_3 ? _GEN_5151 : _GEN_5055; // @[executor.scala 290:56]
  wire [7:0] _GEN_5248 = 8'h1 < length_3 ? _GEN_5152 : _GEN_5056; // @[executor.scala 290:56]
  wire [7:0] _GEN_5249 = 8'h1 < length_3 ? _GEN_5153 : _GEN_5057; // @[executor.scala 290:56]
  wire [7:0] _GEN_5250 = 8'h1 < length_3 ? _GEN_5154 : _GEN_5058; // @[executor.scala 290:56]
  wire [7:0] _GEN_5251 = 8'h1 < length_3 ? _GEN_5155 : _GEN_5059; // @[executor.scala 290:56]
  wire [7:0] _GEN_5252 = 8'h1 < length_3 ? _GEN_5156 : _GEN_5060; // @[executor.scala 290:56]
  wire [7:0] _GEN_5253 = 8'h1 < length_3 ? _GEN_5157 : _GEN_5061; // @[executor.scala 290:56]
  wire [7:0] _GEN_5254 = 8'h1 < length_3 ? _GEN_5158 : _GEN_5062; // @[executor.scala 290:56]
  wire [7:0] _GEN_5255 = 8'h1 < length_3 ? _GEN_5159 : _GEN_5063; // @[executor.scala 290:56]
  wire [7:0] _GEN_5256 = 8'h1 < length_3 ? _GEN_5160 : _GEN_5064; // @[executor.scala 290:56]
  wire [7:0] _GEN_5257 = 8'h1 < length_3 ? _GEN_5161 : _GEN_5065; // @[executor.scala 290:56]
  wire [7:0] _GEN_5258 = 8'h1 < length_3 ? _GEN_5162 : _GEN_5066; // @[executor.scala 290:56]
  wire [7:0] _GEN_5259 = 8'h1 < length_3 ? _GEN_5163 : _GEN_5067; // @[executor.scala 290:56]
  wire [7:0] _GEN_5260 = 8'h1 < length_3 ? _GEN_5164 : _GEN_5068; // @[executor.scala 290:56]
  wire [7:0] _GEN_5261 = 8'h1 < length_3 ? _GEN_5165 : _GEN_5069; // @[executor.scala 290:56]
  wire [7:0] _GEN_5262 = 8'h1 < length_3 ? _GEN_5166 : _GEN_5070; // @[executor.scala 290:56]
  wire [7:0] _GEN_5263 = 8'h1 < length_3 ? _GEN_5167 : _GEN_5071; // @[executor.scala 290:56]
  wire [7:0] _GEN_5264 = 8'h1 < length_3 ? _GEN_5168 : _GEN_5072; // @[executor.scala 290:56]
  wire [7:0] _GEN_5265 = 8'h1 < length_3 ? _GEN_5169 : _GEN_5073; // @[executor.scala 290:56]
  wire [7:0] _GEN_5266 = 8'h1 < length_3 ? _GEN_5170 : _GEN_5074; // @[executor.scala 290:56]
  wire [7:0] _GEN_5267 = 8'h1 < length_3 ? _GEN_5171 : _GEN_5075; // @[executor.scala 290:56]
  wire [7:0] _GEN_5268 = 8'h1 < length_3 ? _GEN_5172 : _GEN_5076; // @[executor.scala 290:56]
  wire [7:0] _GEN_5269 = 8'h1 < length_3 ? _GEN_5173 : _GEN_5077; // @[executor.scala 290:56]
  wire [7:0] _GEN_5270 = 8'h1 < length_3 ? _GEN_5174 : _GEN_5078; // @[executor.scala 290:56]
  wire [7:0] _GEN_5271 = 8'h1 < length_3 ? _GEN_5175 : _GEN_5079; // @[executor.scala 290:56]
  wire [7:0] _GEN_5272 = 8'h1 < length_3 ? _GEN_5176 : _GEN_5080; // @[executor.scala 290:56]
  wire [7:0] _GEN_5273 = 8'h1 < length_3 ? _GEN_5177 : _GEN_5081; // @[executor.scala 290:56]
  wire [7:0] _GEN_5274 = 8'h1 < length_3 ? _GEN_5178 : _GEN_5082; // @[executor.scala 290:56]
  wire [7:0] _GEN_5275 = 8'h1 < length_3 ? _GEN_5179 : _GEN_5083; // @[executor.scala 290:56]
  wire [7:0] _GEN_5276 = 8'h1 < length_3 ? _GEN_5180 : _GEN_5084; // @[executor.scala 290:56]
  wire [7:0] _GEN_5277 = 8'h1 < length_3 ? _GEN_5181 : _GEN_5085; // @[executor.scala 290:56]
  wire [7:0] _GEN_5278 = 8'h1 < length_3 ? _GEN_5182 : _GEN_5086; // @[executor.scala 290:56]
  wire [7:0] _GEN_5279 = 8'h1 < length_3 ? _GEN_5183 : _GEN_5087; // @[executor.scala 290:56]
  wire [7:0] _GEN_5280 = 8'h1 < length_3 ? _GEN_5184 : _GEN_5088; // @[executor.scala 290:56]
  wire [7:0] _GEN_5281 = 8'h1 < length_3 ? _GEN_5185 : _GEN_5089; // @[executor.scala 290:56]
  wire [7:0] _GEN_5282 = 8'h1 < length_3 ? _GEN_5186 : _GEN_5090; // @[executor.scala 290:56]
  wire [7:0] field_byte_26 = field_3[47:40]; // @[executor.scala 287:53]
  wire [7:0] total_offset_26 = offset_3 + 8'h2; // @[executor.scala 289:53]
  wire [7:0] _GEN_5283 = 7'h0 == total_offset_26[6:0] ? field_byte_26 : _GEN_5187; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5284 = 7'h1 == total_offset_26[6:0] ? field_byte_26 : _GEN_5188; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5285 = 7'h2 == total_offset_26[6:0] ? field_byte_26 : _GEN_5189; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5286 = 7'h3 == total_offset_26[6:0] ? field_byte_26 : _GEN_5190; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5287 = 7'h4 == total_offset_26[6:0] ? field_byte_26 : _GEN_5191; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5288 = 7'h5 == total_offset_26[6:0] ? field_byte_26 : _GEN_5192; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5289 = 7'h6 == total_offset_26[6:0] ? field_byte_26 : _GEN_5193; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5290 = 7'h7 == total_offset_26[6:0] ? field_byte_26 : _GEN_5194; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5291 = 7'h8 == total_offset_26[6:0] ? field_byte_26 : _GEN_5195; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5292 = 7'h9 == total_offset_26[6:0] ? field_byte_26 : _GEN_5196; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5293 = 7'ha == total_offset_26[6:0] ? field_byte_26 : _GEN_5197; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5294 = 7'hb == total_offset_26[6:0] ? field_byte_26 : _GEN_5198; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5295 = 7'hc == total_offset_26[6:0] ? field_byte_26 : _GEN_5199; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5296 = 7'hd == total_offset_26[6:0] ? field_byte_26 : _GEN_5200; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5297 = 7'he == total_offset_26[6:0] ? field_byte_26 : _GEN_5201; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5298 = 7'hf == total_offset_26[6:0] ? field_byte_26 : _GEN_5202; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5299 = 7'h10 == total_offset_26[6:0] ? field_byte_26 : _GEN_5203; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5300 = 7'h11 == total_offset_26[6:0] ? field_byte_26 : _GEN_5204; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5301 = 7'h12 == total_offset_26[6:0] ? field_byte_26 : _GEN_5205; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5302 = 7'h13 == total_offset_26[6:0] ? field_byte_26 : _GEN_5206; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5303 = 7'h14 == total_offset_26[6:0] ? field_byte_26 : _GEN_5207; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5304 = 7'h15 == total_offset_26[6:0] ? field_byte_26 : _GEN_5208; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5305 = 7'h16 == total_offset_26[6:0] ? field_byte_26 : _GEN_5209; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5306 = 7'h17 == total_offset_26[6:0] ? field_byte_26 : _GEN_5210; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5307 = 7'h18 == total_offset_26[6:0] ? field_byte_26 : _GEN_5211; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5308 = 7'h19 == total_offset_26[6:0] ? field_byte_26 : _GEN_5212; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5309 = 7'h1a == total_offset_26[6:0] ? field_byte_26 : _GEN_5213; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5310 = 7'h1b == total_offset_26[6:0] ? field_byte_26 : _GEN_5214; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5311 = 7'h1c == total_offset_26[6:0] ? field_byte_26 : _GEN_5215; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5312 = 7'h1d == total_offset_26[6:0] ? field_byte_26 : _GEN_5216; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5313 = 7'h1e == total_offset_26[6:0] ? field_byte_26 : _GEN_5217; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5314 = 7'h1f == total_offset_26[6:0] ? field_byte_26 : _GEN_5218; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5315 = 7'h20 == total_offset_26[6:0] ? field_byte_26 : _GEN_5219; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5316 = 7'h21 == total_offset_26[6:0] ? field_byte_26 : _GEN_5220; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5317 = 7'h22 == total_offset_26[6:0] ? field_byte_26 : _GEN_5221; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5318 = 7'h23 == total_offset_26[6:0] ? field_byte_26 : _GEN_5222; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5319 = 7'h24 == total_offset_26[6:0] ? field_byte_26 : _GEN_5223; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5320 = 7'h25 == total_offset_26[6:0] ? field_byte_26 : _GEN_5224; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5321 = 7'h26 == total_offset_26[6:0] ? field_byte_26 : _GEN_5225; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5322 = 7'h27 == total_offset_26[6:0] ? field_byte_26 : _GEN_5226; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5323 = 7'h28 == total_offset_26[6:0] ? field_byte_26 : _GEN_5227; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5324 = 7'h29 == total_offset_26[6:0] ? field_byte_26 : _GEN_5228; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5325 = 7'h2a == total_offset_26[6:0] ? field_byte_26 : _GEN_5229; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5326 = 7'h2b == total_offset_26[6:0] ? field_byte_26 : _GEN_5230; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5327 = 7'h2c == total_offset_26[6:0] ? field_byte_26 : _GEN_5231; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5328 = 7'h2d == total_offset_26[6:0] ? field_byte_26 : _GEN_5232; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5329 = 7'h2e == total_offset_26[6:0] ? field_byte_26 : _GEN_5233; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5330 = 7'h2f == total_offset_26[6:0] ? field_byte_26 : _GEN_5234; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5331 = 7'h30 == total_offset_26[6:0] ? field_byte_26 : _GEN_5235; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5332 = 7'h31 == total_offset_26[6:0] ? field_byte_26 : _GEN_5236; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5333 = 7'h32 == total_offset_26[6:0] ? field_byte_26 : _GEN_5237; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5334 = 7'h33 == total_offset_26[6:0] ? field_byte_26 : _GEN_5238; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5335 = 7'h34 == total_offset_26[6:0] ? field_byte_26 : _GEN_5239; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5336 = 7'h35 == total_offset_26[6:0] ? field_byte_26 : _GEN_5240; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5337 = 7'h36 == total_offset_26[6:0] ? field_byte_26 : _GEN_5241; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5338 = 7'h37 == total_offset_26[6:0] ? field_byte_26 : _GEN_5242; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5339 = 7'h38 == total_offset_26[6:0] ? field_byte_26 : _GEN_5243; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5340 = 7'h39 == total_offset_26[6:0] ? field_byte_26 : _GEN_5244; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5341 = 7'h3a == total_offset_26[6:0] ? field_byte_26 : _GEN_5245; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5342 = 7'h3b == total_offset_26[6:0] ? field_byte_26 : _GEN_5246; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5343 = 7'h3c == total_offset_26[6:0] ? field_byte_26 : _GEN_5247; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5344 = 7'h3d == total_offset_26[6:0] ? field_byte_26 : _GEN_5248; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5345 = 7'h3e == total_offset_26[6:0] ? field_byte_26 : _GEN_5249; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5346 = 7'h3f == total_offset_26[6:0] ? field_byte_26 : _GEN_5250; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5347 = 7'h40 == total_offset_26[6:0] ? field_byte_26 : _GEN_5251; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5348 = 7'h41 == total_offset_26[6:0] ? field_byte_26 : _GEN_5252; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5349 = 7'h42 == total_offset_26[6:0] ? field_byte_26 : _GEN_5253; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5350 = 7'h43 == total_offset_26[6:0] ? field_byte_26 : _GEN_5254; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5351 = 7'h44 == total_offset_26[6:0] ? field_byte_26 : _GEN_5255; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5352 = 7'h45 == total_offset_26[6:0] ? field_byte_26 : _GEN_5256; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5353 = 7'h46 == total_offset_26[6:0] ? field_byte_26 : _GEN_5257; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5354 = 7'h47 == total_offset_26[6:0] ? field_byte_26 : _GEN_5258; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5355 = 7'h48 == total_offset_26[6:0] ? field_byte_26 : _GEN_5259; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5356 = 7'h49 == total_offset_26[6:0] ? field_byte_26 : _GEN_5260; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5357 = 7'h4a == total_offset_26[6:0] ? field_byte_26 : _GEN_5261; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5358 = 7'h4b == total_offset_26[6:0] ? field_byte_26 : _GEN_5262; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5359 = 7'h4c == total_offset_26[6:0] ? field_byte_26 : _GEN_5263; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5360 = 7'h4d == total_offset_26[6:0] ? field_byte_26 : _GEN_5264; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5361 = 7'h4e == total_offset_26[6:0] ? field_byte_26 : _GEN_5265; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5362 = 7'h4f == total_offset_26[6:0] ? field_byte_26 : _GEN_5266; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5363 = 7'h50 == total_offset_26[6:0] ? field_byte_26 : _GEN_5267; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5364 = 7'h51 == total_offset_26[6:0] ? field_byte_26 : _GEN_5268; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5365 = 7'h52 == total_offset_26[6:0] ? field_byte_26 : _GEN_5269; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5366 = 7'h53 == total_offset_26[6:0] ? field_byte_26 : _GEN_5270; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5367 = 7'h54 == total_offset_26[6:0] ? field_byte_26 : _GEN_5271; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5368 = 7'h55 == total_offset_26[6:0] ? field_byte_26 : _GEN_5272; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5369 = 7'h56 == total_offset_26[6:0] ? field_byte_26 : _GEN_5273; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5370 = 7'h57 == total_offset_26[6:0] ? field_byte_26 : _GEN_5274; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5371 = 7'h58 == total_offset_26[6:0] ? field_byte_26 : _GEN_5275; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5372 = 7'h59 == total_offset_26[6:0] ? field_byte_26 : _GEN_5276; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5373 = 7'h5a == total_offset_26[6:0] ? field_byte_26 : _GEN_5277; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5374 = 7'h5b == total_offset_26[6:0] ? field_byte_26 : _GEN_5278; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5375 = 7'h5c == total_offset_26[6:0] ? field_byte_26 : _GEN_5279; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5376 = 7'h5d == total_offset_26[6:0] ? field_byte_26 : _GEN_5280; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5377 = 7'h5e == total_offset_26[6:0] ? field_byte_26 : _GEN_5281; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5378 = 7'h5f == total_offset_26[6:0] ? field_byte_26 : _GEN_5282; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5379 = 8'h2 < length_3 ? _GEN_5283 : _GEN_5187; // @[executor.scala 290:56]
  wire [7:0] _GEN_5380 = 8'h2 < length_3 ? _GEN_5284 : _GEN_5188; // @[executor.scala 290:56]
  wire [7:0] _GEN_5381 = 8'h2 < length_3 ? _GEN_5285 : _GEN_5189; // @[executor.scala 290:56]
  wire [7:0] _GEN_5382 = 8'h2 < length_3 ? _GEN_5286 : _GEN_5190; // @[executor.scala 290:56]
  wire [7:0] _GEN_5383 = 8'h2 < length_3 ? _GEN_5287 : _GEN_5191; // @[executor.scala 290:56]
  wire [7:0] _GEN_5384 = 8'h2 < length_3 ? _GEN_5288 : _GEN_5192; // @[executor.scala 290:56]
  wire [7:0] _GEN_5385 = 8'h2 < length_3 ? _GEN_5289 : _GEN_5193; // @[executor.scala 290:56]
  wire [7:0] _GEN_5386 = 8'h2 < length_3 ? _GEN_5290 : _GEN_5194; // @[executor.scala 290:56]
  wire [7:0] _GEN_5387 = 8'h2 < length_3 ? _GEN_5291 : _GEN_5195; // @[executor.scala 290:56]
  wire [7:0] _GEN_5388 = 8'h2 < length_3 ? _GEN_5292 : _GEN_5196; // @[executor.scala 290:56]
  wire [7:0] _GEN_5389 = 8'h2 < length_3 ? _GEN_5293 : _GEN_5197; // @[executor.scala 290:56]
  wire [7:0] _GEN_5390 = 8'h2 < length_3 ? _GEN_5294 : _GEN_5198; // @[executor.scala 290:56]
  wire [7:0] _GEN_5391 = 8'h2 < length_3 ? _GEN_5295 : _GEN_5199; // @[executor.scala 290:56]
  wire [7:0] _GEN_5392 = 8'h2 < length_3 ? _GEN_5296 : _GEN_5200; // @[executor.scala 290:56]
  wire [7:0] _GEN_5393 = 8'h2 < length_3 ? _GEN_5297 : _GEN_5201; // @[executor.scala 290:56]
  wire [7:0] _GEN_5394 = 8'h2 < length_3 ? _GEN_5298 : _GEN_5202; // @[executor.scala 290:56]
  wire [7:0] _GEN_5395 = 8'h2 < length_3 ? _GEN_5299 : _GEN_5203; // @[executor.scala 290:56]
  wire [7:0] _GEN_5396 = 8'h2 < length_3 ? _GEN_5300 : _GEN_5204; // @[executor.scala 290:56]
  wire [7:0] _GEN_5397 = 8'h2 < length_3 ? _GEN_5301 : _GEN_5205; // @[executor.scala 290:56]
  wire [7:0] _GEN_5398 = 8'h2 < length_3 ? _GEN_5302 : _GEN_5206; // @[executor.scala 290:56]
  wire [7:0] _GEN_5399 = 8'h2 < length_3 ? _GEN_5303 : _GEN_5207; // @[executor.scala 290:56]
  wire [7:0] _GEN_5400 = 8'h2 < length_3 ? _GEN_5304 : _GEN_5208; // @[executor.scala 290:56]
  wire [7:0] _GEN_5401 = 8'h2 < length_3 ? _GEN_5305 : _GEN_5209; // @[executor.scala 290:56]
  wire [7:0] _GEN_5402 = 8'h2 < length_3 ? _GEN_5306 : _GEN_5210; // @[executor.scala 290:56]
  wire [7:0] _GEN_5403 = 8'h2 < length_3 ? _GEN_5307 : _GEN_5211; // @[executor.scala 290:56]
  wire [7:0] _GEN_5404 = 8'h2 < length_3 ? _GEN_5308 : _GEN_5212; // @[executor.scala 290:56]
  wire [7:0] _GEN_5405 = 8'h2 < length_3 ? _GEN_5309 : _GEN_5213; // @[executor.scala 290:56]
  wire [7:0] _GEN_5406 = 8'h2 < length_3 ? _GEN_5310 : _GEN_5214; // @[executor.scala 290:56]
  wire [7:0] _GEN_5407 = 8'h2 < length_3 ? _GEN_5311 : _GEN_5215; // @[executor.scala 290:56]
  wire [7:0] _GEN_5408 = 8'h2 < length_3 ? _GEN_5312 : _GEN_5216; // @[executor.scala 290:56]
  wire [7:0] _GEN_5409 = 8'h2 < length_3 ? _GEN_5313 : _GEN_5217; // @[executor.scala 290:56]
  wire [7:0] _GEN_5410 = 8'h2 < length_3 ? _GEN_5314 : _GEN_5218; // @[executor.scala 290:56]
  wire [7:0] _GEN_5411 = 8'h2 < length_3 ? _GEN_5315 : _GEN_5219; // @[executor.scala 290:56]
  wire [7:0] _GEN_5412 = 8'h2 < length_3 ? _GEN_5316 : _GEN_5220; // @[executor.scala 290:56]
  wire [7:0] _GEN_5413 = 8'h2 < length_3 ? _GEN_5317 : _GEN_5221; // @[executor.scala 290:56]
  wire [7:0] _GEN_5414 = 8'h2 < length_3 ? _GEN_5318 : _GEN_5222; // @[executor.scala 290:56]
  wire [7:0] _GEN_5415 = 8'h2 < length_3 ? _GEN_5319 : _GEN_5223; // @[executor.scala 290:56]
  wire [7:0] _GEN_5416 = 8'h2 < length_3 ? _GEN_5320 : _GEN_5224; // @[executor.scala 290:56]
  wire [7:0] _GEN_5417 = 8'h2 < length_3 ? _GEN_5321 : _GEN_5225; // @[executor.scala 290:56]
  wire [7:0] _GEN_5418 = 8'h2 < length_3 ? _GEN_5322 : _GEN_5226; // @[executor.scala 290:56]
  wire [7:0] _GEN_5419 = 8'h2 < length_3 ? _GEN_5323 : _GEN_5227; // @[executor.scala 290:56]
  wire [7:0] _GEN_5420 = 8'h2 < length_3 ? _GEN_5324 : _GEN_5228; // @[executor.scala 290:56]
  wire [7:0] _GEN_5421 = 8'h2 < length_3 ? _GEN_5325 : _GEN_5229; // @[executor.scala 290:56]
  wire [7:0] _GEN_5422 = 8'h2 < length_3 ? _GEN_5326 : _GEN_5230; // @[executor.scala 290:56]
  wire [7:0] _GEN_5423 = 8'h2 < length_3 ? _GEN_5327 : _GEN_5231; // @[executor.scala 290:56]
  wire [7:0] _GEN_5424 = 8'h2 < length_3 ? _GEN_5328 : _GEN_5232; // @[executor.scala 290:56]
  wire [7:0] _GEN_5425 = 8'h2 < length_3 ? _GEN_5329 : _GEN_5233; // @[executor.scala 290:56]
  wire [7:0] _GEN_5426 = 8'h2 < length_3 ? _GEN_5330 : _GEN_5234; // @[executor.scala 290:56]
  wire [7:0] _GEN_5427 = 8'h2 < length_3 ? _GEN_5331 : _GEN_5235; // @[executor.scala 290:56]
  wire [7:0] _GEN_5428 = 8'h2 < length_3 ? _GEN_5332 : _GEN_5236; // @[executor.scala 290:56]
  wire [7:0] _GEN_5429 = 8'h2 < length_3 ? _GEN_5333 : _GEN_5237; // @[executor.scala 290:56]
  wire [7:0] _GEN_5430 = 8'h2 < length_3 ? _GEN_5334 : _GEN_5238; // @[executor.scala 290:56]
  wire [7:0] _GEN_5431 = 8'h2 < length_3 ? _GEN_5335 : _GEN_5239; // @[executor.scala 290:56]
  wire [7:0] _GEN_5432 = 8'h2 < length_3 ? _GEN_5336 : _GEN_5240; // @[executor.scala 290:56]
  wire [7:0] _GEN_5433 = 8'h2 < length_3 ? _GEN_5337 : _GEN_5241; // @[executor.scala 290:56]
  wire [7:0] _GEN_5434 = 8'h2 < length_3 ? _GEN_5338 : _GEN_5242; // @[executor.scala 290:56]
  wire [7:0] _GEN_5435 = 8'h2 < length_3 ? _GEN_5339 : _GEN_5243; // @[executor.scala 290:56]
  wire [7:0] _GEN_5436 = 8'h2 < length_3 ? _GEN_5340 : _GEN_5244; // @[executor.scala 290:56]
  wire [7:0] _GEN_5437 = 8'h2 < length_3 ? _GEN_5341 : _GEN_5245; // @[executor.scala 290:56]
  wire [7:0] _GEN_5438 = 8'h2 < length_3 ? _GEN_5342 : _GEN_5246; // @[executor.scala 290:56]
  wire [7:0] _GEN_5439 = 8'h2 < length_3 ? _GEN_5343 : _GEN_5247; // @[executor.scala 290:56]
  wire [7:0] _GEN_5440 = 8'h2 < length_3 ? _GEN_5344 : _GEN_5248; // @[executor.scala 290:56]
  wire [7:0] _GEN_5441 = 8'h2 < length_3 ? _GEN_5345 : _GEN_5249; // @[executor.scala 290:56]
  wire [7:0] _GEN_5442 = 8'h2 < length_3 ? _GEN_5346 : _GEN_5250; // @[executor.scala 290:56]
  wire [7:0] _GEN_5443 = 8'h2 < length_3 ? _GEN_5347 : _GEN_5251; // @[executor.scala 290:56]
  wire [7:0] _GEN_5444 = 8'h2 < length_3 ? _GEN_5348 : _GEN_5252; // @[executor.scala 290:56]
  wire [7:0] _GEN_5445 = 8'h2 < length_3 ? _GEN_5349 : _GEN_5253; // @[executor.scala 290:56]
  wire [7:0] _GEN_5446 = 8'h2 < length_3 ? _GEN_5350 : _GEN_5254; // @[executor.scala 290:56]
  wire [7:0] _GEN_5447 = 8'h2 < length_3 ? _GEN_5351 : _GEN_5255; // @[executor.scala 290:56]
  wire [7:0] _GEN_5448 = 8'h2 < length_3 ? _GEN_5352 : _GEN_5256; // @[executor.scala 290:56]
  wire [7:0] _GEN_5449 = 8'h2 < length_3 ? _GEN_5353 : _GEN_5257; // @[executor.scala 290:56]
  wire [7:0] _GEN_5450 = 8'h2 < length_3 ? _GEN_5354 : _GEN_5258; // @[executor.scala 290:56]
  wire [7:0] _GEN_5451 = 8'h2 < length_3 ? _GEN_5355 : _GEN_5259; // @[executor.scala 290:56]
  wire [7:0] _GEN_5452 = 8'h2 < length_3 ? _GEN_5356 : _GEN_5260; // @[executor.scala 290:56]
  wire [7:0] _GEN_5453 = 8'h2 < length_3 ? _GEN_5357 : _GEN_5261; // @[executor.scala 290:56]
  wire [7:0] _GEN_5454 = 8'h2 < length_3 ? _GEN_5358 : _GEN_5262; // @[executor.scala 290:56]
  wire [7:0] _GEN_5455 = 8'h2 < length_3 ? _GEN_5359 : _GEN_5263; // @[executor.scala 290:56]
  wire [7:0] _GEN_5456 = 8'h2 < length_3 ? _GEN_5360 : _GEN_5264; // @[executor.scala 290:56]
  wire [7:0] _GEN_5457 = 8'h2 < length_3 ? _GEN_5361 : _GEN_5265; // @[executor.scala 290:56]
  wire [7:0] _GEN_5458 = 8'h2 < length_3 ? _GEN_5362 : _GEN_5266; // @[executor.scala 290:56]
  wire [7:0] _GEN_5459 = 8'h2 < length_3 ? _GEN_5363 : _GEN_5267; // @[executor.scala 290:56]
  wire [7:0] _GEN_5460 = 8'h2 < length_3 ? _GEN_5364 : _GEN_5268; // @[executor.scala 290:56]
  wire [7:0] _GEN_5461 = 8'h2 < length_3 ? _GEN_5365 : _GEN_5269; // @[executor.scala 290:56]
  wire [7:0] _GEN_5462 = 8'h2 < length_3 ? _GEN_5366 : _GEN_5270; // @[executor.scala 290:56]
  wire [7:0] _GEN_5463 = 8'h2 < length_3 ? _GEN_5367 : _GEN_5271; // @[executor.scala 290:56]
  wire [7:0] _GEN_5464 = 8'h2 < length_3 ? _GEN_5368 : _GEN_5272; // @[executor.scala 290:56]
  wire [7:0] _GEN_5465 = 8'h2 < length_3 ? _GEN_5369 : _GEN_5273; // @[executor.scala 290:56]
  wire [7:0] _GEN_5466 = 8'h2 < length_3 ? _GEN_5370 : _GEN_5274; // @[executor.scala 290:56]
  wire [7:0] _GEN_5467 = 8'h2 < length_3 ? _GEN_5371 : _GEN_5275; // @[executor.scala 290:56]
  wire [7:0] _GEN_5468 = 8'h2 < length_3 ? _GEN_5372 : _GEN_5276; // @[executor.scala 290:56]
  wire [7:0] _GEN_5469 = 8'h2 < length_3 ? _GEN_5373 : _GEN_5277; // @[executor.scala 290:56]
  wire [7:0] _GEN_5470 = 8'h2 < length_3 ? _GEN_5374 : _GEN_5278; // @[executor.scala 290:56]
  wire [7:0] _GEN_5471 = 8'h2 < length_3 ? _GEN_5375 : _GEN_5279; // @[executor.scala 290:56]
  wire [7:0] _GEN_5472 = 8'h2 < length_3 ? _GEN_5376 : _GEN_5280; // @[executor.scala 290:56]
  wire [7:0] _GEN_5473 = 8'h2 < length_3 ? _GEN_5377 : _GEN_5281; // @[executor.scala 290:56]
  wire [7:0] _GEN_5474 = 8'h2 < length_3 ? _GEN_5378 : _GEN_5282; // @[executor.scala 290:56]
  wire [7:0] field_byte_27 = field_3[39:32]; // @[executor.scala 287:53]
  wire [7:0] total_offset_27 = offset_3 + 8'h3; // @[executor.scala 289:53]
  wire [7:0] _GEN_5475 = 7'h0 == total_offset_27[6:0] ? field_byte_27 : _GEN_5379; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5476 = 7'h1 == total_offset_27[6:0] ? field_byte_27 : _GEN_5380; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5477 = 7'h2 == total_offset_27[6:0] ? field_byte_27 : _GEN_5381; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5478 = 7'h3 == total_offset_27[6:0] ? field_byte_27 : _GEN_5382; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5479 = 7'h4 == total_offset_27[6:0] ? field_byte_27 : _GEN_5383; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5480 = 7'h5 == total_offset_27[6:0] ? field_byte_27 : _GEN_5384; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5481 = 7'h6 == total_offset_27[6:0] ? field_byte_27 : _GEN_5385; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5482 = 7'h7 == total_offset_27[6:0] ? field_byte_27 : _GEN_5386; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5483 = 7'h8 == total_offset_27[6:0] ? field_byte_27 : _GEN_5387; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5484 = 7'h9 == total_offset_27[6:0] ? field_byte_27 : _GEN_5388; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5485 = 7'ha == total_offset_27[6:0] ? field_byte_27 : _GEN_5389; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5486 = 7'hb == total_offset_27[6:0] ? field_byte_27 : _GEN_5390; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5487 = 7'hc == total_offset_27[6:0] ? field_byte_27 : _GEN_5391; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5488 = 7'hd == total_offset_27[6:0] ? field_byte_27 : _GEN_5392; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5489 = 7'he == total_offset_27[6:0] ? field_byte_27 : _GEN_5393; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5490 = 7'hf == total_offset_27[6:0] ? field_byte_27 : _GEN_5394; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5491 = 7'h10 == total_offset_27[6:0] ? field_byte_27 : _GEN_5395; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5492 = 7'h11 == total_offset_27[6:0] ? field_byte_27 : _GEN_5396; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5493 = 7'h12 == total_offset_27[6:0] ? field_byte_27 : _GEN_5397; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5494 = 7'h13 == total_offset_27[6:0] ? field_byte_27 : _GEN_5398; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5495 = 7'h14 == total_offset_27[6:0] ? field_byte_27 : _GEN_5399; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5496 = 7'h15 == total_offset_27[6:0] ? field_byte_27 : _GEN_5400; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5497 = 7'h16 == total_offset_27[6:0] ? field_byte_27 : _GEN_5401; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5498 = 7'h17 == total_offset_27[6:0] ? field_byte_27 : _GEN_5402; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5499 = 7'h18 == total_offset_27[6:0] ? field_byte_27 : _GEN_5403; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5500 = 7'h19 == total_offset_27[6:0] ? field_byte_27 : _GEN_5404; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5501 = 7'h1a == total_offset_27[6:0] ? field_byte_27 : _GEN_5405; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5502 = 7'h1b == total_offset_27[6:0] ? field_byte_27 : _GEN_5406; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5503 = 7'h1c == total_offset_27[6:0] ? field_byte_27 : _GEN_5407; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5504 = 7'h1d == total_offset_27[6:0] ? field_byte_27 : _GEN_5408; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5505 = 7'h1e == total_offset_27[6:0] ? field_byte_27 : _GEN_5409; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5506 = 7'h1f == total_offset_27[6:0] ? field_byte_27 : _GEN_5410; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5507 = 7'h20 == total_offset_27[6:0] ? field_byte_27 : _GEN_5411; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5508 = 7'h21 == total_offset_27[6:0] ? field_byte_27 : _GEN_5412; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5509 = 7'h22 == total_offset_27[6:0] ? field_byte_27 : _GEN_5413; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5510 = 7'h23 == total_offset_27[6:0] ? field_byte_27 : _GEN_5414; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5511 = 7'h24 == total_offset_27[6:0] ? field_byte_27 : _GEN_5415; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5512 = 7'h25 == total_offset_27[6:0] ? field_byte_27 : _GEN_5416; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5513 = 7'h26 == total_offset_27[6:0] ? field_byte_27 : _GEN_5417; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5514 = 7'h27 == total_offset_27[6:0] ? field_byte_27 : _GEN_5418; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5515 = 7'h28 == total_offset_27[6:0] ? field_byte_27 : _GEN_5419; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5516 = 7'h29 == total_offset_27[6:0] ? field_byte_27 : _GEN_5420; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5517 = 7'h2a == total_offset_27[6:0] ? field_byte_27 : _GEN_5421; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5518 = 7'h2b == total_offset_27[6:0] ? field_byte_27 : _GEN_5422; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5519 = 7'h2c == total_offset_27[6:0] ? field_byte_27 : _GEN_5423; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5520 = 7'h2d == total_offset_27[6:0] ? field_byte_27 : _GEN_5424; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5521 = 7'h2e == total_offset_27[6:0] ? field_byte_27 : _GEN_5425; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5522 = 7'h2f == total_offset_27[6:0] ? field_byte_27 : _GEN_5426; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5523 = 7'h30 == total_offset_27[6:0] ? field_byte_27 : _GEN_5427; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5524 = 7'h31 == total_offset_27[6:0] ? field_byte_27 : _GEN_5428; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5525 = 7'h32 == total_offset_27[6:0] ? field_byte_27 : _GEN_5429; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5526 = 7'h33 == total_offset_27[6:0] ? field_byte_27 : _GEN_5430; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5527 = 7'h34 == total_offset_27[6:0] ? field_byte_27 : _GEN_5431; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5528 = 7'h35 == total_offset_27[6:0] ? field_byte_27 : _GEN_5432; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5529 = 7'h36 == total_offset_27[6:0] ? field_byte_27 : _GEN_5433; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5530 = 7'h37 == total_offset_27[6:0] ? field_byte_27 : _GEN_5434; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5531 = 7'h38 == total_offset_27[6:0] ? field_byte_27 : _GEN_5435; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5532 = 7'h39 == total_offset_27[6:0] ? field_byte_27 : _GEN_5436; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5533 = 7'h3a == total_offset_27[6:0] ? field_byte_27 : _GEN_5437; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5534 = 7'h3b == total_offset_27[6:0] ? field_byte_27 : _GEN_5438; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5535 = 7'h3c == total_offset_27[6:0] ? field_byte_27 : _GEN_5439; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5536 = 7'h3d == total_offset_27[6:0] ? field_byte_27 : _GEN_5440; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5537 = 7'h3e == total_offset_27[6:0] ? field_byte_27 : _GEN_5441; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5538 = 7'h3f == total_offset_27[6:0] ? field_byte_27 : _GEN_5442; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5539 = 7'h40 == total_offset_27[6:0] ? field_byte_27 : _GEN_5443; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5540 = 7'h41 == total_offset_27[6:0] ? field_byte_27 : _GEN_5444; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5541 = 7'h42 == total_offset_27[6:0] ? field_byte_27 : _GEN_5445; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5542 = 7'h43 == total_offset_27[6:0] ? field_byte_27 : _GEN_5446; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5543 = 7'h44 == total_offset_27[6:0] ? field_byte_27 : _GEN_5447; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5544 = 7'h45 == total_offset_27[6:0] ? field_byte_27 : _GEN_5448; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5545 = 7'h46 == total_offset_27[6:0] ? field_byte_27 : _GEN_5449; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5546 = 7'h47 == total_offset_27[6:0] ? field_byte_27 : _GEN_5450; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5547 = 7'h48 == total_offset_27[6:0] ? field_byte_27 : _GEN_5451; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5548 = 7'h49 == total_offset_27[6:0] ? field_byte_27 : _GEN_5452; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5549 = 7'h4a == total_offset_27[6:0] ? field_byte_27 : _GEN_5453; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5550 = 7'h4b == total_offset_27[6:0] ? field_byte_27 : _GEN_5454; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5551 = 7'h4c == total_offset_27[6:0] ? field_byte_27 : _GEN_5455; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5552 = 7'h4d == total_offset_27[6:0] ? field_byte_27 : _GEN_5456; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5553 = 7'h4e == total_offset_27[6:0] ? field_byte_27 : _GEN_5457; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5554 = 7'h4f == total_offset_27[6:0] ? field_byte_27 : _GEN_5458; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5555 = 7'h50 == total_offset_27[6:0] ? field_byte_27 : _GEN_5459; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5556 = 7'h51 == total_offset_27[6:0] ? field_byte_27 : _GEN_5460; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5557 = 7'h52 == total_offset_27[6:0] ? field_byte_27 : _GEN_5461; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5558 = 7'h53 == total_offset_27[6:0] ? field_byte_27 : _GEN_5462; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5559 = 7'h54 == total_offset_27[6:0] ? field_byte_27 : _GEN_5463; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5560 = 7'h55 == total_offset_27[6:0] ? field_byte_27 : _GEN_5464; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5561 = 7'h56 == total_offset_27[6:0] ? field_byte_27 : _GEN_5465; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5562 = 7'h57 == total_offset_27[6:0] ? field_byte_27 : _GEN_5466; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5563 = 7'h58 == total_offset_27[6:0] ? field_byte_27 : _GEN_5467; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5564 = 7'h59 == total_offset_27[6:0] ? field_byte_27 : _GEN_5468; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5565 = 7'h5a == total_offset_27[6:0] ? field_byte_27 : _GEN_5469; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5566 = 7'h5b == total_offset_27[6:0] ? field_byte_27 : _GEN_5470; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5567 = 7'h5c == total_offset_27[6:0] ? field_byte_27 : _GEN_5471; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5568 = 7'h5d == total_offset_27[6:0] ? field_byte_27 : _GEN_5472; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5569 = 7'h5e == total_offset_27[6:0] ? field_byte_27 : _GEN_5473; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5570 = 7'h5f == total_offset_27[6:0] ? field_byte_27 : _GEN_5474; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5571 = 8'h3 < length_3 ? _GEN_5475 : _GEN_5379; // @[executor.scala 290:56]
  wire [7:0] _GEN_5572 = 8'h3 < length_3 ? _GEN_5476 : _GEN_5380; // @[executor.scala 290:56]
  wire [7:0] _GEN_5573 = 8'h3 < length_3 ? _GEN_5477 : _GEN_5381; // @[executor.scala 290:56]
  wire [7:0] _GEN_5574 = 8'h3 < length_3 ? _GEN_5478 : _GEN_5382; // @[executor.scala 290:56]
  wire [7:0] _GEN_5575 = 8'h3 < length_3 ? _GEN_5479 : _GEN_5383; // @[executor.scala 290:56]
  wire [7:0] _GEN_5576 = 8'h3 < length_3 ? _GEN_5480 : _GEN_5384; // @[executor.scala 290:56]
  wire [7:0] _GEN_5577 = 8'h3 < length_3 ? _GEN_5481 : _GEN_5385; // @[executor.scala 290:56]
  wire [7:0] _GEN_5578 = 8'h3 < length_3 ? _GEN_5482 : _GEN_5386; // @[executor.scala 290:56]
  wire [7:0] _GEN_5579 = 8'h3 < length_3 ? _GEN_5483 : _GEN_5387; // @[executor.scala 290:56]
  wire [7:0] _GEN_5580 = 8'h3 < length_3 ? _GEN_5484 : _GEN_5388; // @[executor.scala 290:56]
  wire [7:0] _GEN_5581 = 8'h3 < length_3 ? _GEN_5485 : _GEN_5389; // @[executor.scala 290:56]
  wire [7:0] _GEN_5582 = 8'h3 < length_3 ? _GEN_5486 : _GEN_5390; // @[executor.scala 290:56]
  wire [7:0] _GEN_5583 = 8'h3 < length_3 ? _GEN_5487 : _GEN_5391; // @[executor.scala 290:56]
  wire [7:0] _GEN_5584 = 8'h3 < length_3 ? _GEN_5488 : _GEN_5392; // @[executor.scala 290:56]
  wire [7:0] _GEN_5585 = 8'h3 < length_3 ? _GEN_5489 : _GEN_5393; // @[executor.scala 290:56]
  wire [7:0] _GEN_5586 = 8'h3 < length_3 ? _GEN_5490 : _GEN_5394; // @[executor.scala 290:56]
  wire [7:0] _GEN_5587 = 8'h3 < length_3 ? _GEN_5491 : _GEN_5395; // @[executor.scala 290:56]
  wire [7:0] _GEN_5588 = 8'h3 < length_3 ? _GEN_5492 : _GEN_5396; // @[executor.scala 290:56]
  wire [7:0] _GEN_5589 = 8'h3 < length_3 ? _GEN_5493 : _GEN_5397; // @[executor.scala 290:56]
  wire [7:0] _GEN_5590 = 8'h3 < length_3 ? _GEN_5494 : _GEN_5398; // @[executor.scala 290:56]
  wire [7:0] _GEN_5591 = 8'h3 < length_3 ? _GEN_5495 : _GEN_5399; // @[executor.scala 290:56]
  wire [7:0] _GEN_5592 = 8'h3 < length_3 ? _GEN_5496 : _GEN_5400; // @[executor.scala 290:56]
  wire [7:0] _GEN_5593 = 8'h3 < length_3 ? _GEN_5497 : _GEN_5401; // @[executor.scala 290:56]
  wire [7:0] _GEN_5594 = 8'h3 < length_3 ? _GEN_5498 : _GEN_5402; // @[executor.scala 290:56]
  wire [7:0] _GEN_5595 = 8'h3 < length_3 ? _GEN_5499 : _GEN_5403; // @[executor.scala 290:56]
  wire [7:0] _GEN_5596 = 8'h3 < length_3 ? _GEN_5500 : _GEN_5404; // @[executor.scala 290:56]
  wire [7:0] _GEN_5597 = 8'h3 < length_3 ? _GEN_5501 : _GEN_5405; // @[executor.scala 290:56]
  wire [7:0] _GEN_5598 = 8'h3 < length_3 ? _GEN_5502 : _GEN_5406; // @[executor.scala 290:56]
  wire [7:0] _GEN_5599 = 8'h3 < length_3 ? _GEN_5503 : _GEN_5407; // @[executor.scala 290:56]
  wire [7:0] _GEN_5600 = 8'h3 < length_3 ? _GEN_5504 : _GEN_5408; // @[executor.scala 290:56]
  wire [7:0] _GEN_5601 = 8'h3 < length_3 ? _GEN_5505 : _GEN_5409; // @[executor.scala 290:56]
  wire [7:0] _GEN_5602 = 8'h3 < length_3 ? _GEN_5506 : _GEN_5410; // @[executor.scala 290:56]
  wire [7:0] _GEN_5603 = 8'h3 < length_3 ? _GEN_5507 : _GEN_5411; // @[executor.scala 290:56]
  wire [7:0] _GEN_5604 = 8'h3 < length_3 ? _GEN_5508 : _GEN_5412; // @[executor.scala 290:56]
  wire [7:0] _GEN_5605 = 8'h3 < length_3 ? _GEN_5509 : _GEN_5413; // @[executor.scala 290:56]
  wire [7:0] _GEN_5606 = 8'h3 < length_3 ? _GEN_5510 : _GEN_5414; // @[executor.scala 290:56]
  wire [7:0] _GEN_5607 = 8'h3 < length_3 ? _GEN_5511 : _GEN_5415; // @[executor.scala 290:56]
  wire [7:0] _GEN_5608 = 8'h3 < length_3 ? _GEN_5512 : _GEN_5416; // @[executor.scala 290:56]
  wire [7:0] _GEN_5609 = 8'h3 < length_3 ? _GEN_5513 : _GEN_5417; // @[executor.scala 290:56]
  wire [7:0] _GEN_5610 = 8'h3 < length_3 ? _GEN_5514 : _GEN_5418; // @[executor.scala 290:56]
  wire [7:0] _GEN_5611 = 8'h3 < length_3 ? _GEN_5515 : _GEN_5419; // @[executor.scala 290:56]
  wire [7:0] _GEN_5612 = 8'h3 < length_3 ? _GEN_5516 : _GEN_5420; // @[executor.scala 290:56]
  wire [7:0] _GEN_5613 = 8'h3 < length_3 ? _GEN_5517 : _GEN_5421; // @[executor.scala 290:56]
  wire [7:0] _GEN_5614 = 8'h3 < length_3 ? _GEN_5518 : _GEN_5422; // @[executor.scala 290:56]
  wire [7:0] _GEN_5615 = 8'h3 < length_3 ? _GEN_5519 : _GEN_5423; // @[executor.scala 290:56]
  wire [7:0] _GEN_5616 = 8'h3 < length_3 ? _GEN_5520 : _GEN_5424; // @[executor.scala 290:56]
  wire [7:0] _GEN_5617 = 8'h3 < length_3 ? _GEN_5521 : _GEN_5425; // @[executor.scala 290:56]
  wire [7:0] _GEN_5618 = 8'h3 < length_3 ? _GEN_5522 : _GEN_5426; // @[executor.scala 290:56]
  wire [7:0] _GEN_5619 = 8'h3 < length_3 ? _GEN_5523 : _GEN_5427; // @[executor.scala 290:56]
  wire [7:0] _GEN_5620 = 8'h3 < length_3 ? _GEN_5524 : _GEN_5428; // @[executor.scala 290:56]
  wire [7:0] _GEN_5621 = 8'h3 < length_3 ? _GEN_5525 : _GEN_5429; // @[executor.scala 290:56]
  wire [7:0] _GEN_5622 = 8'h3 < length_3 ? _GEN_5526 : _GEN_5430; // @[executor.scala 290:56]
  wire [7:0] _GEN_5623 = 8'h3 < length_3 ? _GEN_5527 : _GEN_5431; // @[executor.scala 290:56]
  wire [7:0] _GEN_5624 = 8'h3 < length_3 ? _GEN_5528 : _GEN_5432; // @[executor.scala 290:56]
  wire [7:0] _GEN_5625 = 8'h3 < length_3 ? _GEN_5529 : _GEN_5433; // @[executor.scala 290:56]
  wire [7:0] _GEN_5626 = 8'h3 < length_3 ? _GEN_5530 : _GEN_5434; // @[executor.scala 290:56]
  wire [7:0] _GEN_5627 = 8'h3 < length_3 ? _GEN_5531 : _GEN_5435; // @[executor.scala 290:56]
  wire [7:0] _GEN_5628 = 8'h3 < length_3 ? _GEN_5532 : _GEN_5436; // @[executor.scala 290:56]
  wire [7:0] _GEN_5629 = 8'h3 < length_3 ? _GEN_5533 : _GEN_5437; // @[executor.scala 290:56]
  wire [7:0] _GEN_5630 = 8'h3 < length_3 ? _GEN_5534 : _GEN_5438; // @[executor.scala 290:56]
  wire [7:0] _GEN_5631 = 8'h3 < length_3 ? _GEN_5535 : _GEN_5439; // @[executor.scala 290:56]
  wire [7:0] _GEN_5632 = 8'h3 < length_3 ? _GEN_5536 : _GEN_5440; // @[executor.scala 290:56]
  wire [7:0] _GEN_5633 = 8'h3 < length_3 ? _GEN_5537 : _GEN_5441; // @[executor.scala 290:56]
  wire [7:0] _GEN_5634 = 8'h3 < length_3 ? _GEN_5538 : _GEN_5442; // @[executor.scala 290:56]
  wire [7:0] _GEN_5635 = 8'h3 < length_3 ? _GEN_5539 : _GEN_5443; // @[executor.scala 290:56]
  wire [7:0] _GEN_5636 = 8'h3 < length_3 ? _GEN_5540 : _GEN_5444; // @[executor.scala 290:56]
  wire [7:0] _GEN_5637 = 8'h3 < length_3 ? _GEN_5541 : _GEN_5445; // @[executor.scala 290:56]
  wire [7:0] _GEN_5638 = 8'h3 < length_3 ? _GEN_5542 : _GEN_5446; // @[executor.scala 290:56]
  wire [7:0] _GEN_5639 = 8'h3 < length_3 ? _GEN_5543 : _GEN_5447; // @[executor.scala 290:56]
  wire [7:0] _GEN_5640 = 8'h3 < length_3 ? _GEN_5544 : _GEN_5448; // @[executor.scala 290:56]
  wire [7:0] _GEN_5641 = 8'h3 < length_3 ? _GEN_5545 : _GEN_5449; // @[executor.scala 290:56]
  wire [7:0] _GEN_5642 = 8'h3 < length_3 ? _GEN_5546 : _GEN_5450; // @[executor.scala 290:56]
  wire [7:0] _GEN_5643 = 8'h3 < length_3 ? _GEN_5547 : _GEN_5451; // @[executor.scala 290:56]
  wire [7:0] _GEN_5644 = 8'h3 < length_3 ? _GEN_5548 : _GEN_5452; // @[executor.scala 290:56]
  wire [7:0] _GEN_5645 = 8'h3 < length_3 ? _GEN_5549 : _GEN_5453; // @[executor.scala 290:56]
  wire [7:0] _GEN_5646 = 8'h3 < length_3 ? _GEN_5550 : _GEN_5454; // @[executor.scala 290:56]
  wire [7:0] _GEN_5647 = 8'h3 < length_3 ? _GEN_5551 : _GEN_5455; // @[executor.scala 290:56]
  wire [7:0] _GEN_5648 = 8'h3 < length_3 ? _GEN_5552 : _GEN_5456; // @[executor.scala 290:56]
  wire [7:0] _GEN_5649 = 8'h3 < length_3 ? _GEN_5553 : _GEN_5457; // @[executor.scala 290:56]
  wire [7:0] _GEN_5650 = 8'h3 < length_3 ? _GEN_5554 : _GEN_5458; // @[executor.scala 290:56]
  wire [7:0] _GEN_5651 = 8'h3 < length_3 ? _GEN_5555 : _GEN_5459; // @[executor.scala 290:56]
  wire [7:0] _GEN_5652 = 8'h3 < length_3 ? _GEN_5556 : _GEN_5460; // @[executor.scala 290:56]
  wire [7:0] _GEN_5653 = 8'h3 < length_3 ? _GEN_5557 : _GEN_5461; // @[executor.scala 290:56]
  wire [7:0] _GEN_5654 = 8'h3 < length_3 ? _GEN_5558 : _GEN_5462; // @[executor.scala 290:56]
  wire [7:0] _GEN_5655 = 8'h3 < length_3 ? _GEN_5559 : _GEN_5463; // @[executor.scala 290:56]
  wire [7:0] _GEN_5656 = 8'h3 < length_3 ? _GEN_5560 : _GEN_5464; // @[executor.scala 290:56]
  wire [7:0] _GEN_5657 = 8'h3 < length_3 ? _GEN_5561 : _GEN_5465; // @[executor.scala 290:56]
  wire [7:0] _GEN_5658 = 8'h3 < length_3 ? _GEN_5562 : _GEN_5466; // @[executor.scala 290:56]
  wire [7:0] _GEN_5659 = 8'h3 < length_3 ? _GEN_5563 : _GEN_5467; // @[executor.scala 290:56]
  wire [7:0] _GEN_5660 = 8'h3 < length_3 ? _GEN_5564 : _GEN_5468; // @[executor.scala 290:56]
  wire [7:0] _GEN_5661 = 8'h3 < length_3 ? _GEN_5565 : _GEN_5469; // @[executor.scala 290:56]
  wire [7:0] _GEN_5662 = 8'h3 < length_3 ? _GEN_5566 : _GEN_5470; // @[executor.scala 290:56]
  wire [7:0] _GEN_5663 = 8'h3 < length_3 ? _GEN_5567 : _GEN_5471; // @[executor.scala 290:56]
  wire [7:0] _GEN_5664 = 8'h3 < length_3 ? _GEN_5568 : _GEN_5472; // @[executor.scala 290:56]
  wire [7:0] _GEN_5665 = 8'h3 < length_3 ? _GEN_5569 : _GEN_5473; // @[executor.scala 290:56]
  wire [7:0] _GEN_5666 = 8'h3 < length_3 ? _GEN_5570 : _GEN_5474; // @[executor.scala 290:56]
  wire [7:0] field_byte_28 = field_3[31:24]; // @[executor.scala 287:53]
  wire [7:0] total_offset_28 = offset_3 + 8'h4; // @[executor.scala 289:53]
  wire [7:0] _GEN_5667 = 7'h0 == total_offset_28[6:0] ? field_byte_28 : _GEN_5571; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5668 = 7'h1 == total_offset_28[6:0] ? field_byte_28 : _GEN_5572; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5669 = 7'h2 == total_offset_28[6:0] ? field_byte_28 : _GEN_5573; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5670 = 7'h3 == total_offset_28[6:0] ? field_byte_28 : _GEN_5574; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5671 = 7'h4 == total_offset_28[6:0] ? field_byte_28 : _GEN_5575; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5672 = 7'h5 == total_offset_28[6:0] ? field_byte_28 : _GEN_5576; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5673 = 7'h6 == total_offset_28[6:0] ? field_byte_28 : _GEN_5577; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5674 = 7'h7 == total_offset_28[6:0] ? field_byte_28 : _GEN_5578; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5675 = 7'h8 == total_offset_28[6:0] ? field_byte_28 : _GEN_5579; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5676 = 7'h9 == total_offset_28[6:0] ? field_byte_28 : _GEN_5580; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5677 = 7'ha == total_offset_28[6:0] ? field_byte_28 : _GEN_5581; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5678 = 7'hb == total_offset_28[6:0] ? field_byte_28 : _GEN_5582; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5679 = 7'hc == total_offset_28[6:0] ? field_byte_28 : _GEN_5583; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5680 = 7'hd == total_offset_28[6:0] ? field_byte_28 : _GEN_5584; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5681 = 7'he == total_offset_28[6:0] ? field_byte_28 : _GEN_5585; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5682 = 7'hf == total_offset_28[6:0] ? field_byte_28 : _GEN_5586; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5683 = 7'h10 == total_offset_28[6:0] ? field_byte_28 : _GEN_5587; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5684 = 7'h11 == total_offset_28[6:0] ? field_byte_28 : _GEN_5588; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5685 = 7'h12 == total_offset_28[6:0] ? field_byte_28 : _GEN_5589; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5686 = 7'h13 == total_offset_28[6:0] ? field_byte_28 : _GEN_5590; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5687 = 7'h14 == total_offset_28[6:0] ? field_byte_28 : _GEN_5591; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5688 = 7'h15 == total_offset_28[6:0] ? field_byte_28 : _GEN_5592; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5689 = 7'h16 == total_offset_28[6:0] ? field_byte_28 : _GEN_5593; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5690 = 7'h17 == total_offset_28[6:0] ? field_byte_28 : _GEN_5594; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5691 = 7'h18 == total_offset_28[6:0] ? field_byte_28 : _GEN_5595; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5692 = 7'h19 == total_offset_28[6:0] ? field_byte_28 : _GEN_5596; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5693 = 7'h1a == total_offset_28[6:0] ? field_byte_28 : _GEN_5597; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5694 = 7'h1b == total_offset_28[6:0] ? field_byte_28 : _GEN_5598; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5695 = 7'h1c == total_offset_28[6:0] ? field_byte_28 : _GEN_5599; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5696 = 7'h1d == total_offset_28[6:0] ? field_byte_28 : _GEN_5600; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5697 = 7'h1e == total_offset_28[6:0] ? field_byte_28 : _GEN_5601; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5698 = 7'h1f == total_offset_28[6:0] ? field_byte_28 : _GEN_5602; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5699 = 7'h20 == total_offset_28[6:0] ? field_byte_28 : _GEN_5603; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5700 = 7'h21 == total_offset_28[6:0] ? field_byte_28 : _GEN_5604; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5701 = 7'h22 == total_offset_28[6:0] ? field_byte_28 : _GEN_5605; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5702 = 7'h23 == total_offset_28[6:0] ? field_byte_28 : _GEN_5606; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5703 = 7'h24 == total_offset_28[6:0] ? field_byte_28 : _GEN_5607; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5704 = 7'h25 == total_offset_28[6:0] ? field_byte_28 : _GEN_5608; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5705 = 7'h26 == total_offset_28[6:0] ? field_byte_28 : _GEN_5609; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5706 = 7'h27 == total_offset_28[6:0] ? field_byte_28 : _GEN_5610; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5707 = 7'h28 == total_offset_28[6:0] ? field_byte_28 : _GEN_5611; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5708 = 7'h29 == total_offset_28[6:0] ? field_byte_28 : _GEN_5612; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5709 = 7'h2a == total_offset_28[6:0] ? field_byte_28 : _GEN_5613; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5710 = 7'h2b == total_offset_28[6:0] ? field_byte_28 : _GEN_5614; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5711 = 7'h2c == total_offset_28[6:0] ? field_byte_28 : _GEN_5615; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5712 = 7'h2d == total_offset_28[6:0] ? field_byte_28 : _GEN_5616; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5713 = 7'h2e == total_offset_28[6:0] ? field_byte_28 : _GEN_5617; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5714 = 7'h2f == total_offset_28[6:0] ? field_byte_28 : _GEN_5618; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5715 = 7'h30 == total_offset_28[6:0] ? field_byte_28 : _GEN_5619; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5716 = 7'h31 == total_offset_28[6:0] ? field_byte_28 : _GEN_5620; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5717 = 7'h32 == total_offset_28[6:0] ? field_byte_28 : _GEN_5621; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5718 = 7'h33 == total_offset_28[6:0] ? field_byte_28 : _GEN_5622; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5719 = 7'h34 == total_offset_28[6:0] ? field_byte_28 : _GEN_5623; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5720 = 7'h35 == total_offset_28[6:0] ? field_byte_28 : _GEN_5624; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5721 = 7'h36 == total_offset_28[6:0] ? field_byte_28 : _GEN_5625; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5722 = 7'h37 == total_offset_28[6:0] ? field_byte_28 : _GEN_5626; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5723 = 7'h38 == total_offset_28[6:0] ? field_byte_28 : _GEN_5627; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5724 = 7'h39 == total_offset_28[6:0] ? field_byte_28 : _GEN_5628; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5725 = 7'h3a == total_offset_28[6:0] ? field_byte_28 : _GEN_5629; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5726 = 7'h3b == total_offset_28[6:0] ? field_byte_28 : _GEN_5630; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5727 = 7'h3c == total_offset_28[6:0] ? field_byte_28 : _GEN_5631; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5728 = 7'h3d == total_offset_28[6:0] ? field_byte_28 : _GEN_5632; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5729 = 7'h3e == total_offset_28[6:0] ? field_byte_28 : _GEN_5633; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5730 = 7'h3f == total_offset_28[6:0] ? field_byte_28 : _GEN_5634; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5731 = 7'h40 == total_offset_28[6:0] ? field_byte_28 : _GEN_5635; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5732 = 7'h41 == total_offset_28[6:0] ? field_byte_28 : _GEN_5636; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5733 = 7'h42 == total_offset_28[6:0] ? field_byte_28 : _GEN_5637; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5734 = 7'h43 == total_offset_28[6:0] ? field_byte_28 : _GEN_5638; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5735 = 7'h44 == total_offset_28[6:0] ? field_byte_28 : _GEN_5639; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5736 = 7'h45 == total_offset_28[6:0] ? field_byte_28 : _GEN_5640; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5737 = 7'h46 == total_offset_28[6:0] ? field_byte_28 : _GEN_5641; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5738 = 7'h47 == total_offset_28[6:0] ? field_byte_28 : _GEN_5642; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5739 = 7'h48 == total_offset_28[6:0] ? field_byte_28 : _GEN_5643; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5740 = 7'h49 == total_offset_28[6:0] ? field_byte_28 : _GEN_5644; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5741 = 7'h4a == total_offset_28[6:0] ? field_byte_28 : _GEN_5645; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5742 = 7'h4b == total_offset_28[6:0] ? field_byte_28 : _GEN_5646; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5743 = 7'h4c == total_offset_28[6:0] ? field_byte_28 : _GEN_5647; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5744 = 7'h4d == total_offset_28[6:0] ? field_byte_28 : _GEN_5648; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5745 = 7'h4e == total_offset_28[6:0] ? field_byte_28 : _GEN_5649; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5746 = 7'h4f == total_offset_28[6:0] ? field_byte_28 : _GEN_5650; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5747 = 7'h50 == total_offset_28[6:0] ? field_byte_28 : _GEN_5651; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5748 = 7'h51 == total_offset_28[6:0] ? field_byte_28 : _GEN_5652; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5749 = 7'h52 == total_offset_28[6:0] ? field_byte_28 : _GEN_5653; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5750 = 7'h53 == total_offset_28[6:0] ? field_byte_28 : _GEN_5654; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5751 = 7'h54 == total_offset_28[6:0] ? field_byte_28 : _GEN_5655; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5752 = 7'h55 == total_offset_28[6:0] ? field_byte_28 : _GEN_5656; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5753 = 7'h56 == total_offset_28[6:0] ? field_byte_28 : _GEN_5657; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5754 = 7'h57 == total_offset_28[6:0] ? field_byte_28 : _GEN_5658; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5755 = 7'h58 == total_offset_28[6:0] ? field_byte_28 : _GEN_5659; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5756 = 7'h59 == total_offset_28[6:0] ? field_byte_28 : _GEN_5660; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5757 = 7'h5a == total_offset_28[6:0] ? field_byte_28 : _GEN_5661; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5758 = 7'h5b == total_offset_28[6:0] ? field_byte_28 : _GEN_5662; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5759 = 7'h5c == total_offset_28[6:0] ? field_byte_28 : _GEN_5663; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5760 = 7'h5d == total_offset_28[6:0] ? field_byte_28 : _GEN_5664; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5761 = 7'h5e == total_offset_28[6:0] ? field_byte_28 : _GEN_5665; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5762 = 7'h5f == total_offset_28[6:0] ? field_byte_28 : _GEN_5666; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5763 = 8'h4 < length_3 ? _GEN_5667 : _GEN_5571; // @[executor.scala 290:56]
  wire [7:0] _GEN_5764 = 8'h4 < length_3 ? _GEN_5668 : _GEN_5572; // @[executor.scala 290:56]
  wire [7:0] _GEN_5765 = 8'h4 < length_3 ? _GEN_5669 : _GEN_5573; // @[executor.scala 290:56]
  wire [7:0] _GEN_5766 = 8'h4 < length_3 ? _GEN_5670 : _GEN_5574; // @[executor.scala 290:56]
  wire [7:0] _GEN_5767 = 8'h4 < length_3 ? _GEN_5671 : _GEN_5575; // @[executor.scala 290:56]
  wire [7:0] _GEN_5768 = 8'h4 < length_3 ? _GEN_5672 : _GEN_5576; // @[executor.scala 290:56]
  wire [7:0] _GEN_5769 = 8'h4 < length_3 ? _GEN_5673 : _GEN_5577; // @[executor.scala 290:56]
  wire [7:0] _GEN_5770 = 8'h4 < length_3 ? _GEN_5674 : _GEN_5578; // @[executor.scala 290:56]
  wire [7:0] _GEN_5771 = 8'h4 < length_3 ? _GEN_5675 : _GEN_5579; // @[executor.scala 290:56]
  wire [7:0] _GEN_5772 = 8'h4 < length_3 ? _GEN_5676 : _GEN_5580; // @[executor.scala 290:56]
  wire [7:0] _GEN_5773 = 8'h4 < length_3 ? _GEN_5677 : _GEN_5581; // @[executor.scala 290:56]
  wire [7:0] _GEN_5774 = 8'h4 < length_3 ? _GEN_5678 : _GEN_5582; // @[executor.scala 290:56]
  wire [7:0] _GEN_5775 = 8'h4 < length_3 ? _GEN_5679 : _GEN_5583; // @[executor.scala 290:56]
  wire [7:0] _GEN_5776 = 8'h4 < length_3 ? _GEN_5680 : _GEN_5584; // @[executor.scala 290:56]
  wire [7:0] _GEN_5777 = 8'h4 < length_3 ? _GEN_5681 : _GEN_5585; // @[executor.scala 290:56]
  wire [7:0] _GEN_5778 = 8'h4 < length_3 ? _GEN_5682 : _GEN_5586; // @[executor.scala 290:56]
  wire [7:0] _GEN_5779 = 8'h4 < length_3 ? _GEN_5683 : _GEN_5587; // @[executor.scala 290:56]
  wire [7:0] _GEN_5780 = 8'h4 < length_3 ? _GEN_5684 : _GEN_5588; // @[executor.scala 290:56]
  wire [7:0] _GEN_5781 = 8'h4 < length_3 ? _GEN_5685 : _GEN_5589; // @[executor.scala 290:56]
  wire [7:0] _GEN_5782 = 8'h4 < length_3 ? _GEN_5686 : _GEN_5590; // @[executor.scala 290:56]
  wire [7:0] _GEN_5783 = 8'h4 < length_3 ? _GEN_5687 : _GEN_5591; // @[executor.scala 290:56]
  wire [7:0] _GEN_5784 = 8'h4 < length_3 ? _GEN_5688 : _GEN_5592; // @[executor.scala 290:56]
  wire [7:0] _GEN_5785 = 8'h4 < length_3 ? _GEN_5689 : _GEN_5593; // @[executor.scala 290:56]
  wire [7:0] _GEN_5786 = 8'h4 < length_3 ? _GEN_5690 : _GEN_5594; // @[executor.scala 290:56]
  wire [7:0] _GEN_5787 = 8'h4 < length_3 ? _GEN_5691 : _GEN_5595; // @[executor.scala 290:56]
  wire [7:0] _GEN_5788 = 8'h4 < length_3 ? _GEN_5692 : _GEN_5596; // @[executor.scala 290:56]
  wire [7:0] _GEN_5789 = 8'h4 < length_3 ? _GEN_5693 : _GEN_5597; // @[executor.scala 290:56]
  wire [7:0] _GEN_5790 = 8'h4 < length_3 ? _GEN_5694 : _GEN_5598; // @[executor.scala 290:56]
  wire [7:0] _GEN_5791 = 8'h4 < length_3 ? _GEN_5695 : _GEN_5599; // @[executor.scala 290:56]
  wire [7:0] _GEN_5792 = 8'h4 < length_3 ? _GEN_5696 : _GEN_5600; // @[executor.scala 290:56]
  wire [7:0] _GEN_5793 = 8'h4 < length_3 ? _GEN_5697 : _GEN_5601; // @[executor.scala 290:56]
  wire [7:0] _GEN_5794 = 8'h4 < length_3 ? _GEN_5698 : _GEN_5602; // @[executor.scala 290:56]
  wire [7:0] _GEN_5795 = 8'h4 < length_3 ? _GEN_5699 : _GEN_5603; // @[executor.scala 290:56]
  wire [7:0] _GEN_5796 = 8'h4 < length_3 ? _GEN_5700 : _GEN_5604; // @[executor.scala 290:56]
  wire [7:0] _GEN_5797 = 8'h4 < length_3 ? _GEN_5701 : _GEN_5605; // @[executor.scala 290:56]
  wire [7:0] _GEN_5798 = 8'h4 < length_3 ? _GEN_5702 : _GEN_5606; // @[executor.scala 290:56]
  wire [7:0] _GEN_5799 = 8'h4 < length_3 ? _GEN_5703 : _GEN_5607; // @[executor.scala 290:56]
  wire [7:0] _GEN_5800 = 8'h4 < length_3 ? _GEN_5704 : _GEN_5608; // @[executor.scala 290:56]
  wire [7:0] _GEN_5801 = 8'h4 < length_3 ? _GEN_5705 : _GEN_5609; // @[executor.scala 290:56]
  wire [7:0] _GEN_5802 = 8'h4 < length_3 ? _GEN_5706 : _GEN_5610; // @[executor.scala 290:56]
  wire [7:0] _GEN_5803 = 8'h4 < length_3 ? _GEN_5707 : _GEN_5611; // @[executor.scala 290:56]
  wire [7:0] _GEN_5804 = 8'h4 < length_3 ? _GEN_5708 : _GEN_5612; // @[executor.scala 290:56]
  wire [7:0] _GEN_5805 = 8'h4 < length_3 ? _GEN_5709 : _GEN_5613; // @[executor.scala 290:56]
  wire [7:0] _GEN_5806 = 8'h4 < length_3 ? _GEN_5710 : _GEN_5614; // @[executor.scala 290:56]
  wire [7:0] _GEN_5807 = 8'h4 < length_3 ? _GEN_5711 : _GEN_5615; // @[executor.scala 290:56]
  wire [7:0] _GEN_5808 = 8'h4 < length_3 ? _GEN_5712 : _GEN_5616; // @[executor.scala 290:56]
  wire [7:0] _GEN_5809 = 8'h4 < length_3 ? _GEN_5713 : _GEN_5617; // @[executor.scala 290:56]
  wire [7:0] _GEN_5810 = 8'h4 < length_3 ? _GEN_5714 : _GEN_5618; // @[executor.scala 290:56]
  wire [7:0] _GEN_5811 = 8'h4 < length_3 ? _GEN_5715 : _GEN_5619; // @[executor.scala 290:56]
  wire [7:0] _GEN_5812 = 8'h4 < length_3 ? _GEN_5716 : _GEN_5620; // @[executor.scala 290:56]
  wire [7:0] _GEN_5813 = 8'h4 < length_3 ? _GEN_5717 : _GEN_5621; // @[executor.scala 290:56]
  wire [7:0] _GEN_5814 = 8'h4 < length_3 ? _GEN_5718 : _GEN_5622; // @[executor.scala 290:56]
  wire [7:0] _GEN_5815 = 8'h4 < length_3 ? _GEN_5719 : _GEN_5623; // @[executor.scala 290:56]
  wire [7:0] _GEN_5816 = 8'h4 < length_3 ? _GEN_5720 : _GEN_5624; // @[executor.scala 290:56]
  wire [7:0] _GEN_5817 = 8'h4 < length_3 ? _GEN_5721 : _GEN_5625; // @[executor.scala 290:56]
  wire [7:0] _GEN_5818 = 8'h4 < length_3 ? _GEN_5722 : _GEN_5626; // @[executor.scala 290:56]
  wire [7:0] _GEN_5819 = 8'h4 < length_3 ? _GEN_5723 : _GEN_5627; // @[executor.scala 290:56]
  wire [7:0] _GEN_5820 = 8'h4 < length_3 ? _GEN_5724 : _GEN_5628; // @[executor.scala 290:56]
  wire [7:0] _GEN_5821 = 8'h4 < length_3 ? _GEN_5725 : _GEN_5629; // @[executor.scala 290:56]
  wire [7:0] _GEN_5822 = 8'h4 < length_3 ? _GEN_5726 : _GEN_5630; // @[executor.scala 290:56]
  wire [7:0] _GEN_5823 = 8'h4 < length_3 ? _GEN_5727 : _GEN_5631; // @[executor.scala 290:56]
  wire [7:0] _GEN_5824 = 8'h4 < length_3 ? _GEN_5728 : _GEN_5632; // @[executor.scala 290:56]
  wire [7:0] _GEN_5825 = 8'h4 < length_3 ? _GEN_5729 : _GEN_5633; // @[executor.scala 290:56]
  wire [7:0] _GEN_5826 = 8'h4 < length_3 ? _GEN_5730 : _GEN_5634; // @[executor.scala 290:56]
  wire [7:0] _GEN_5827 = 8'h4 < length_3 ? _GEN_5731 : _GEN_5635; // @[executor.scala 290:56]
  wire [7:0] _GEN_5828 = 8'h4 < length_3 ? _GEN_5732 : _GEN_5636; // @[executor.scala 290:56]
  wire [7:0] _GEN_5829 = 8'h4 < length_3 ? _GEN_5733 : _GEN_5637; // @[executor.scala 290:56]
  wire [7:0] _GEN_5830 = 8'h4 < length_3 ? _GEN_5734 : _GEN_5638; // @[executor.scala 290:56]
  wire [7:0] _GEN_5831 = 8'h4 < length_3 ? _GEN_5735 : _GEN_5639; // @[executor.scala 290:56]
  wire [7:0] _GEN_5832 = 8'h4 < length_3 ? _GEN_5736 : _GEN_5640; // @[executor.scala 290:56]
  wire [7:0] _GEN_5833 = 8'h4 < length_3 ? _GEN_5737 : _GEN_5641; // @[executor.scala 290:56]
  wire [7:0] _GEN_5834 = 8'h4 < length_3 ? _GEN_5738 : _GEN_5642; // @[executor.scala 290:56]
  wire [7:0] _GEN_5835 = 8'h4 < length_3 ? _GEN_5739 : _GEN_5643; // @[executor.scala 290:56]
  wire [7:0] _GEN_5836 = 8'h4 < length_3 ? _GEN_5740 : _GEN_5644; // @[executor.scala 290:56]
  wire [7:0] _GEN_5837 = 8'h4 < length_3 ? _GEN_5741 : _GEN_5645; // @[executor.scala 290:56]
  wire [7:0] _GEN_5838 = 8'h4 < length_3 ? _GEN_5742 : _GEN_5646; // @[executor.scala 290:56]
  wire [7:0] _GEN_5839 = 8'h4 < length_3 ? _GEN_5743 : _GEN_5647; // @[executor.scala 290:56]
  wire [7:0] _GEN_5840 = 8'h4 < length_3 ? _GEN_5744 : _GEN_5648; // @[executor.scala 290:56]
  wire [7:0] _GEN_5841 = 8'h4 < length_3 ? _GEN_5745 : _GEN_5649; // @[executor.scala 290:56]
  wire [7:0] _GEN_5842 = 8'h4 < length_3 ? _GEN_5746 : _GEN_5650; // @[executor.scala 290:56]
  wire [7:0] _GEN_5843 = 8'h4 < length_3 ? _GEN_5747 : _GEN_5651; // @[executor.scala 290:56]
  wire [7:0] _GEN_5844 = 8'h4 < length_3 ? _GEN_5748 : _GEN_5652; // @[executor.scala 290:56]
  wire [7:0] _GEN_5845 = 8'h4 < length_3 ? _GEN_5749 : _GEN_5653; // @[executor.scala 290:56]
  wire [7:0] _GEN_5846 = 8'h4 < length_3 ? _GEN_5750 : _GEN_5654; // @[executor.scala 290:56]
  wire [7:0] _GEN_5847 = 8'h4 < length_3 ? _GEN_5751 : _GEN_5655; // @[executor.scala 290:56]
  wire [7:0] _GEN_5848 = 8'h4 < length_3 ? _GEN_5752 : _GEN_5656; // @[executor.scala 290:56]
  wire [7:0] _GEN_5849 = 8'h4 < length_3 ? _GEN_5753 : _GEN_5657; // @[executor.scala 290:56]
  wire [7:0] _GEN_5850 = 8'h4 < length_3 ? _GEN_5754 : _GEN_5658; // @[executor.scala 290:56]
  wire [7:0] _GEN_5851 = 8'h4 < length_3 ? _GEN_5755 : _GEN_5659; // @[executor.scala 290:56]
  wire [7:0] _GEN_5852 = 8'h4 < length_3 ? _GEN_5756 : _GEN_5660; // @[executor.scala 290:56]
  wire [7:0] _GEN_5853 = 8'h4 < length_3 ? _GEN_5757 : _GEN_5661; // @[executor.scala 290:56]
  wire [7:0] _GEN_5854 = 8'h4 < length_3 ? _GEN_5758 : _GEN_5662; // @[executor.scala 290:56]
  wire [7:0] _GEN_5855 = 8'h4 < length_3 ? _GEN_5759 : _GEN_5663; // @[executor.scala 290:56]
  wire [7:0] _GEN_5856 = 8'h4 < length_3 ? _GEN_5760 : _GEN_5664; // @[executor.scala 290:56]
  wire [7:0] _GEN_5857 = 8'h4 < length_3 ? _GEN_5761 : _GEN_5665; // @[executor.scala 290:56]
  wire [7:0] _GEN_5858 = 8'h4 < length_3 ? _GEN_5762 : _GEN_5666; // @[executor.scala 290:56]
  wire [7:0] field_byte_29 = field_3[23:16]; // @[executor.scala 287:53]
  wire [7:0] total_offset_29 = offset_3 + 8'h5; // @[executor.scala 289:53]
  wire [7:0] _GEN_5859 = 7'h0 == total_offset_29[6:0] ? field_byte_29 : _GEN_5763; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5860 = 7'h1 == total_offset_29[6:0] ? field_byte_29 : _GEN_5764; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5861 = 7'h2 == total_offset_29[6:0] ? field_byte_29 : _GEN_5765; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5862 = 7'h3 == total_offset_29[6:0] ? field_byte_29 : _GEN_5766; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5863 = 7'h4 == total_offset_29[6:0] ? field_byte_29 : _GEN_5767; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5864 = 7'h5 == total_offset_29[6:0] ? field_byte_29 : _GEN_5768; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5865 = 7'h6 == total_offset_29[6:0] ? field_byte_29 : _GEN_5769; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5866 = 7'h7 == total_offset_29[6:0] ? field_byte_29 : _GEN_5770; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5867 = 7'h8 == total_offset_29[6:0] ? field_byte_29 : _GEN_5771; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5868 = 7'h9 == total_offset_29[6:0] ? field_byte_29 : _GEN_5772; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5869 = 7'ha == total_offset_29[6:0] ? field_byte_29 : _GEN_5773; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5870 = 7'hb == total_offset_29[6:0] ? field_byte_29 : _GEN_5774; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5871 = 7'hc == total_offset_29[6:0] ? field_byte_29 : _GEN_5775; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5872 = 7'hd == total_offset_29[6:0] ? field_byte_29 : _GEN_5776; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5873 = 7'he == total_offset_29[6:0] ? field_byte_29 : _GEN_5777; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5874 = 7'hf == total_offset_29[6:0] ? field_byte_29 : _GEN_5778; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5875 = 7'h10 == total_offset_29[6:0] ? field_byte_29 : _GEN_5779; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5876 = 7'h11 == total_offset_29[6:0] ? field_byte_29 : _GEN_5780; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5877 = 7'h12 == total_offset_29[6:0] ? field_byte_29 : _GEN_5781; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5878 = 7'h13 == total_offset_29[6:0] ? field_byte_29 : _GEN_5782; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5879 = 7'h14 == total_offset_29[6:0] ? field_byte_29 : _GEN_5783; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5880 = 7'h15 == total_offset_29[6:0] ? field_byte_29 : _GEN_5784; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5881 = 7'h16 == total_offset_29[6:0] ? field_byte_29 : _GEN_5785; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5882 = 7'h17 == total_offset_29[6:0] ? field_byte_29 : _GEN_5786; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5883 = 7'h18 == total_offset_29[6:0] ? field_byte_29 : _GEN_5787; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5884 = 7'h19 == total_offset_29[6:0] ? field_byte_29 : _GEN_5788; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5885 = 7'h1a == total_offset_29[6:0] ? field_byte_29 : _GEN_5789; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5886 = 7'h1b == total_offset_29[6:0] ? field_byte_29 : _GEN_5790; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5887 = 7'h1c == total_offset_29[6:0] ? field_byte_29 : _GEN_5791; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5888 = 7'h1d == total_offset_29[6:0] ? field_byte_29 : _GEN_5792; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5889 = 7'h1e == total_offset_29[6:0] ? field_byte_29 : _GEN_5793; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5890 = 7'h1f == total_offset_29[6:0] ? field_byte_29 : _GEN_5794; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5891 = 7'h20 == total_offset_29[6:0] ? field_byte_29 : _GEN_5795; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5892 = 7'h21 == total_offset_29[6:0] ? field_byte_29 : _GEN_5796; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5893 = 7'h22 == total_offset_29[6:0] ? field_byte_29 : _GEN_5797; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5894 = 7'h23 == total_offset_29[6:0] ? field_byte_29 : _GEN_5798; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5895 = 7'h24 == total_offset_29[6:0] ? field_byte_29 : _GEN_5799; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5896 = 7'h25 == total_offset_29[6:0] ? field_byte_29 : _GEN_5800; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5897 = 7'h26 == total_offset_29[6:0] ? field_byte_29 : _GEN_5801; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5898 = 7'h27 == total_offset_29[6:0] ? field_byte_29 : _GEN_5802; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5899 = 7'h28 == total_offset_29[6:0] ? field_byte_29 : _GEN_5803; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5900 = 7'h29 == total_offset_29[6:0] ? field_byte_29 : _GEN_5804; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5901 = 7'h2a == total_offset_29[6:0] ? field_byte_29 : _GEN_5805; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5902 = 7'h2b == total_offset_29[6:0] ? field_byte_29 : _GEN_5806; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5903 = 7'h2c == total_offset_29[6:0] ? field_byte_29 : _GEN_5807; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5904 = 7'h2d == total_offset_29[6:0] ? field_byte_29 : _GEN_5808; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5905 = 7'h2e == total_offset_29[6:0] ? field_byte_29 : _GEN_5809; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5906 = 7'h2f == total_offset_29[6:0] ? field_byte_29 : _GEN_5810; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5907 = 7'h30 == total_offset_29[6:0] ? field_byte_29 : _GEN_5811; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5908 = 7'h31 == total_offset_29[6:0] ? field_byte_29 : _GEN_5812; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5909 = 7'h32 == total_offset_29[6:0] ? field_byte_29 : _GEN_5813; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5910 = 7'h33 == total_offset_29[6:0] ? field_byte_29 : _GEN_5814; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5911 = 7'h34 == total_offset_29[6:0] ? field_byte_29 : _GEN_5815; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5912 = 7'h35 == total_offset_29[6:0] ? field_byte_29 : _GEN_5816; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5913 = 7'h36 == total_offset_29[6:0] ? field_byte_29 : _GEN_5817; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5914 = 7'h37 == total_offset_29[6:0] ? field_byte_29 : _GEN_5818; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5915 = 7'h38 == total_offset_29[6:0] ? field_byte_29 : _GEN_5819; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5916 = 7'h39 == total_offset_29[6:0] ? field_byte_29 : _GEN_5820; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5917 = 7'h3a == total_offset_29[6:0] ? field_byte_29 : _GEN_5821; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5918 = 7'h3b == total_offset_29[6:0] ? field_byte_29 : _GEN_5822; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5919 = 7'h3c == total_offset_29[6:0] ? field_byte_29 : _GEN_5823; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5920 = 7'h3d == total_offset_29[6:0] ? field_byte_29 : _GEN_5824; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5921 = 7'h3e == total_offset_29[6:0] ? field_byte_29 : _GEN_5825; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5922 = 7'h3f == total_offset_29[6:0] ? field_byte_29 : _GEN_5826; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5923 = 7'h40 == total_offset_29[6:0] ? field_byte_29 : _GEN_5827; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5924 = 7'h41 == total_offset_29[6:0] ? field_byte_29 : _GEN_5828; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5925 = 7'h42 == total_offset_29[6:0] ? field_byte_29 : _GEN_5829; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5926 = 7'h43 == total_offset_29[6:0] ? field_byte_29 : _GEN_5830; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5927 = 7'h44 == total_offset_29[6:0] ? field_byte_29 : _GEN_5831; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5928 = 7'h45 == total_offset_29[6:0] ? field_byte_29 : _GEN_5832; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5929 = 7'h46 == total_offset_29[6:0] ? field_byte_29 : _GEN_5833; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5930 = 7'h47 == total_offset_29[6:0] ? field_byte_29 : _GEN_5834; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5931 = 7'h48 == total_offset_29[6:0] ? field_byte_29 : _GEN_5835; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5932 = 7'h49 == total_offset_29[6:0] ? field_byte_29 : _GEN_5836; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5933 = 7'h4a == total_offset_29[6:0] ? field_byte_29 : _GEN_5837; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5934 = 7'h4b == total_offset_29[6:0] ? field_byte_29 : _GEN_5838; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5935 = 7'h4c == total_offset_29[6:0] ? field_byte_29 : _GEN_5839; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5936 = 7'h4d == total_offset_29[6:0] ? field_byte_29 : _GEN_5840; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5937 = 7'h4e == total_offset_29[6:0] ? field_byte_29 : _GEN_5841; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5938 = 7'h4f == total_offset_29[6:0] ? field_byte_29 : _GEN_5842; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5939 = 7'h50 == total_offset_29[6:0] ? field_byte_29 : _GEN_5843; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5940 = 7'h51 == total_offset_29[6:0] ? field_byte_29 : _GEN_5844; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5941 = 7'h52 == total_offset_29[6:0] ? field_byte_29 : _GEN_5845; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5942 = 7'h53 == total_offset_29[6:0] ? field_byte_29 : _GEN_5846; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5943 = 7'h54 == total_offset_29[6:0] ? field_byte_29 : _GEN_5847; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5944 = 7'h55 == total_offset_29[6:0] ? field_byte_29 : _GEN_5848; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5945 = 7'h56 == total_offset_29[6:0] ? field_byte_29 : _GEN_5849; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5946 = 7'h57 == total_offset_29[6:0] ? field_byte_29 : _GEN_5850; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5947 = 7'h58 == total_offset_29[6:0] ? field_byte_29 : _GEN_5851; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5948 = 7'h59 == total_offset_29[6:0] ? field_byte_29 : _GEN_5852; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5949 = 7'h5a == total_offset_29[6:0] ? field_byte_29 : _GEN_5853; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5950 = 7'h5b == total_offset_29[6:0] ? field_byte_29 : _GEN_5854; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5951 = 7'h5c == total_offset_29[6:0] ? field_byte_29 : _GEN_5855; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5952 = 7'h5d == total_offset_29[6:0] ? field_byte_29 : _GEN_5856; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5953 = 7'h5e == total_offset_29[6:0] ? field_byte_29 : _GEN_5857; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5954 = 7'h5f == total_offset_29[6:0] ? field_byte_29 : _GEN_5858; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_5955 = 8'h5 < length_3 ? _GEN_5859 : _GEN_5763; // @[executor.scala 290:56]
  wire [7:0] _GEN_5956 = 8'h5 < length_3 ? _GEN_5860 : _GEN_5764; // @[executor.scala 290:56]
  wire [7:0] _GEN_5957 = 8'h5 < length_3 ? _GEN_5861 : _GEN_5765; // @[executor.scala 290:56]
  wire [7:0] _GEN_5958 = 8'h5 < length_3 ? _GEN_5862 : _GEN_5766; // @[executor.scala 290:56]
  wire [7:0] _GEN_5959 = 8'h5 < length_3 ? _GEN_5863 : _GEN_5767; // @[executor.scala 290:56]
  wire [7:0] _GEN_5960 = 8'h5 < length_3 ? _GEN_5864 : _GEN_5768; // @[executor.scala 290:56]
  wire [7:0] _GEN_5961 = 8'h5 < length_3 ? _GEN_5865 : _GEN_5769; // @[executor.scala 290:56]
  wire [7:0] _GEN_5962 = 8'h5 < length_3 ? _GEN_5866 : _GEN_5770; // @[executor.scala 290:56]
  wire [7:0] _GEN_5963 = 8'h5 < length_3 ? _GEN_5867 : _GEN_5771; // @[executor.scala 290:56]
  wire [7:0] _GEN_5964 = 8'h5 < length_3 ? _GEN_5868 : _GEN_5772; // @[executor.scala 290:56]
  wire [7:0] _GEN_5965 = 8'h5 < length_3 ? _GEN_5869 : _GEN_5773; // @[executor.scala 290:56]
  wire [7:0] _GEN_5966 = 8'h5 < length_3 ? _GEN_5870 : _GEN_5774; // @[executor.scala 290:56]
  wire [7:0] _GEN_5967 = 8'h5 < length_3 ? _GEN_5871 : _GEN_5775; // @[executor.scala 290:56]
  wire [7:0] _GEN_5968 = 8'h5 < length_3 ? _GEN_5872 : _GEN_5776; // @[executor.scala 290:56]
  wire [7:0] _GEN_5969 = 8'h5 < length_3 ? _GEN_5873 : _GEN_5777; // @[executor.scala 290:56]
  wire [7:0] _GEN_5970 = 8'h5 < length_3 ? _GEN_5874 : _GEN_5778; // @[executor.scala 290:56]
  wire [7:0] _GEN_5971 = 8'h5 < length_3 ? _GEN_5875 : _GEN_5779; // @[executor.scala 290:56]
  wire [7:0] _GEN_5972 = 8'h5 < length_3 ? _GEN_5876 : _GEN_5780; // @[executor.scala 290:56]
  wire [7:0] _GEN_5973 = 8'h5 < length_3 ? _GEN_5877 : _GEN_5781; // @[executor.scala 290:56]
  wire [7:0] _GEN_5974 = 8'h5 < length_3 ? _GEN_5878 : _GEN_5782; // @[executor.scala 290:56]
  wire [7:0] _GEN_5975 = 8'h5 < length_3 ? _GEN_5879 : _GEN_5783; // @[executor.scala 290:56]
  wire [7:0] _GEN_5976 = 8'h5 < length_3 ? _GEN_5880 : _GEN_5784; // @[executor.scala 290:56]
  wire [7:0] _GEN_5977 = 8'h5 < length_3 ? _GEN_5881 : _GEN_5785; // @[executor.scala 290:56]
  wire [7:0] _GEN_5978 = 8'h5 < length_3 ? _GEN_5882 : _GEN_5786; // @[executor.scala 290:56]
  wire [7:0] _GEN_5979 = 8'h5 < length_3 ? _GEN_5883 : _GEN_5787; // @[executor.scala 290:56]
  wire [7:0] _GEN_5980 = 8'h5 < length_3 ? _GEN_5884 : _GEN_5788; // @[executor.scala 290:56]
  wire [7:0] _GEN_5981 = 8'h5 < length_3 ? _GEN_5885 : _GEN_5789; // @[executor.scala 290:56]
  wire [7:0] _GEN_5982 = 8'h5 < length_3 ? _GEN_5886 : _GEN_5790; // @[executor.scala 290:56]
  wire [7:0] _GEN_5983 = 8'h5 < length_3 ? _GEN_5887 : _GEN_5791; // @[executor.scala 290:56]
  wire [7:0] _GEN_5984 = 8'h5 < length_3 ? _GEN_5888 : _GEN_5792; // @[executor.scala 290:56]
  wire [7:0] _GEN_5985 = 8'h5 < length_3 ? _GEN_5889 : _GEN_5793; // @[executor.scala 290:56]
  wire [7:0] _GEN_5986 = 8'h5 < length_3 ? _GEN_5890 : _GEN_5794; // @[executor.scala 290:56]
  wire [7:0] _GEN_5987 = 8'h5 < length_3 ? _GEN_5891 : _GEN_5795; // @[executor.scala 290:56]
  wire [7:0] _GEN_5988 = 8'h5 < length_3 ? _GEN_5892 : _GEN_5796; // @[executor.scala 290:56]
  wire [7:0] _GEN_5989 = 8'h5 < length_3 ? _GEN_5893 : _GEN_5797; // @[executor.scala 290:56]
  wire [7:0] _GEN_5990 = 8'h5 < length_3 ? _GEN_5894 : _GEN_5798; // @[executor.scala 290:56]
  wire [7:0] _GEN_5991 = 8'h5 < length_3 ? _GEN_5895 : _GEN_5799; // @[executor.scala 290:56]
  wire [7:0] _GEN_5992 = 8'h5 < length_3 ? _GEN_5896 : _GEN_5800; // @[executor.scala 290:56]
  wire [7:0] _GEN_5993 = 8'h5 < length_3 ? _GEN_5897 : _GEN_5801; // @[executor.scala 290:56]
  wire [7:0] _GEN_5994 = 8'h5 < length_3 ? _GEN_5898 : _GEN_5802; // @[executor.scala 290:56]
  wire [7:0] _GEN_5995 = 8'h5 < length_3 ? _GEN_5899 : _GEN_5803; // @[executor.scala 290:56]
  wire [7:0] _GEN_5996 = 8'h5 < length_3 ? _GEN_5900 : _GEN_5804; // @[executor.scala 290:56]
  wire [7:0] _GEN_5997 = 8'h5 < length_3 ? _GEN_5901 : _GEN_5805; // @[executor.scala 290:56]
  wire [7:0] _GEN_5998 = 8'h5 < length_3 ? _GEN_5902 : _GEN_5806; // @[executor.scala 290:56]
  wire [7:0] _GEN_5999 = 8'h5 < length_3 ? _GEN_5903 : _GEN_5807; // @[executor.scala 290:56]
  wire [7:0] _GEN_6000 = 8'h5 < length_3 ? _GEN_5904 : _GEN_5808; // @[executor.scala 290:56]
  wire [7:0] _GEN_6001 = 8'h5 < length_3 ? _GEN_5905 : _GEN_5809; // @[executor.scala 290:56]
  wire [7:0] _GEN_6002 = 8'h5 < length_3 ? _GEN_5906 : _GEN_5810; // @[executor.scala 290:56]
  wire [7:0] _GEN_6003 = 8'h5 < length_3 ? _GEN_5907 : _GEN_5811; // @[executor.scala 290:56]
  wire [7:0] _GEN_6004 = 8'h5 < length_3 ? _GEN_5908 : _GEN_5812; // @[executor.scala 290:56]
  wire [7:0] _GEN_6005 = 8'h5 < length_3 ? _GEN_5909 : _GEN_5813; // @[executor.scala 290:56]
  wire [7:0] _GEN_6006 = 8'h5 < length_3 ? _GEN_5910 : _GEN_5814; // @[executor.scala 290:56]
  wire [7:0] _GEN_6007 = 8'h5 < length_3 ? _GEN_5911 : _GEN_5815; // @[executor.scala 290:56]
  wire [7:0] _GEN_6008 = 8'h5 < length_3 ? _GEN_5912 : _GEN_5816; // @[executor.scala 290:56]
  wire [7:0] _GEN_6009 = 8'h5 < length_3 ? _GEN_5913 : _GEN_5817; // @[executor.scala 290:56]
  wire [7:0] _GEN_6010 = 8'h5 < length_3 ? _GEN_5914 : _GEN_5818; // @[executor.scala 290:56]
  wire [7:0] _GEN_6011 = 8'h5 < length_3 ? _GEN_5915 : _GEN_5819; // @[executor.scala 290:56]
  wire [7:0] _GEN_6012 = 8'h5 < length_3 ? _GEN_5916 : _GEN_5820; // @[executor.scala 290:56]
  wire [7:0] _GEN_6013 = 8'h5 < length_3 ? _GEN_5917 : _GEN_5821; // @[executor.scala 290:56]
  wire [7:0] _GEN_6014 = 8'h5 < length_3 ? _GEN_5918 : _GEN_5822; // @[executor.scala 290:56]
  wire [7:0] _GEN_6015 = 8'h5 < length_3 ? _GEN_5919 : _GEN_5823; // @[executor.scala 290:56]
  wire [7:0] _GEN_6016 = 8'h5 < length_3 ? _GEN_5920 : _GEN_5824; // @[executor.scala 290:56]
  wire [7:0] _GEN_6017 = 8'h5 < length_3 ? _GEN_5921 : _GEN_5825; // @[executor.scala 290:56]
  wire [7:0] _GEN_6018 = 8'h5 < length_3 ? _GEN_5922 : _GEN_5826; // @[executor.scala 290:56]
  wire [7:0] _GEN_6019 = 8'h5 < length_3 ? _GEN_5923 : _GEN_5827; // @[executor.scala 290:56]
  wire [7:0] _GEN_6020 = 8'h5 < length_3 ? _GEN_5924 : _GEN_5828; // @[executor.scala 290:56]
  wire [7:0] _GEN_6021 = 8'h5 < length_3 ? _GEN_5925 : _GEN_5829; // @[executor.scala 290:56]
  wire [7:0] _GEN_6022 = 8'h5 < length_3 ? _GEN_5926 : _GEN_5830; // @[executor.scala 290:56]
  wire [7:0] _GEN_6023 = 8'h5 < length_3 ? _GEN_5927 : _GEN_5831; // @[executor.scala 290:56]
  wire [7:0] _GEN_6024 = 8'h5 < length_3 ? _GEN_5928 : _GEN_5832; // @[executor.scala 290:56]
  wire [7:0] _GEN_6025 = 8'h5 < length_3 ? _GEN_5929 : _GEN_5833; // @[executor.scala 290:56]
  wire [7:0] _GEN_6026 = 8'h5 < length_3 ? _GEN_5930 : _GEN_5834; // @[executor.scala 290:56]
  wire [7:0] _GEN_6027 = 8'h5 < length_3 ? _GEN_5931 : _GEN_5835; // @[executor.scala 290:56]
  wire [7:0] _GEN_6028 = 8'h5 < length_3 ? _GEN_5932 : _GEN_5836; // @[executor.scala 290:56]
  wire [7:0] _GEN_6029 = 8'h5 < length_3 ? _GEN_5933 : _GEN_5837; // @[executor.scala 290:56]
  wire [7:0] _GEN_6030 = 8'h5 < length_3 ? _GEN_5934 : _GEN_5838; // @[executor.scala 290:56]
  wire [7:0] _GEN_6031 = 8'h5 < length_3 ? _GEN_5935 : _GEN_5839; // @[executor.scala 290:56]
  wire [7:0] _GEN_6032 = 8'h5 < length_3 ? _GEN_5936 : _GEN_5840; // @[executor.scala 290:56]
  wire [7:0] _GEN_6033 = 8'h5 < length_3 ? _GEN_5937 : _GEN_5841; // @[executor.scala 290:56]
  wire [7:0] _GEN_6034 = 8'h5 < length_3 ? _GEN_5938 : _GEN_5842; // @[executor.scala 290:56]
  wire [7:0] _GEN_6035 = 8'h5 < length_3 ? _GEN_5939 : _GEN_5843; // @[executor.scala 290:56]
  wire [7:0] _GEN_6036 = 8'h5 < length_3 ? _GEN_5940 : _GEN_5844; // @[executor.scala 290:56]
  wire [7:0] _GEN_6037 = 8'h5 < length_3 ? _GEN_5941 : _GEN_5845; // @[executor.scala 290:56]
  wire [7:0] _GEN_6038 = 8'h5 < length_3 ? _GEN_5942 : _GEN_5846; // @[executor.scala 290:56]
  wire [7:0] _GEN_6039 = 8'h5 < length_3 ? _GEN_5943 : _GEN_5847; // @[executor.scala 290:56]
  wire [7:0] _GEN_6040 = 8'h5 < length_3 ? _GEN_5944 : _GEN_5848; // @[executor.scala 290:56]
  wire [7:0] _GEN_6041 = 8'h5 < length_3 ? _GEN_5945 : _GEN_5849; // @[executor.scala 290:56]
  wire [7:0] _GEN_6042 = 8'h5 < length_3 ? _GEN_5946 : _GEN_5850; // @[executor.scala 290:56]
  wire [7:0] _GEN_6043 = 8'h5 < length_3 ? _GEN_5947 : _GEN_5851; // @[executor.scala 290:56]
  wire [7:0] _GEN_6044 = 8'h5 < length_3 ? _GEN_5948 : _GEN_5852; // @[executor.scala 290:56]
  wire [7:0] _GEN_6045 = 8'h5 < length_3 ? _GEN_5949 : _GEN_5853; // @[executor.scala 290:56]
  wire [7:0] _GEN_6046 = 8'h5 < length_3 ? _GEN_5950 : _GEN_5854; // @[executor.scala 290:56]
  wire [7:0] _GEN_6047 = 8'h5 < length_3 ? _GEN_5951 : _GEN_5855; // @[executor.scala 290:56]
  wire [7:0] _GEN_6048 = 8'h5 < length_3 ? _GEN_5952 : _GEN_5856; // @[executor.scala 290:56]
  wire [7:0] _GEN_6049 = 8'h5 < length_3 ? _GEN_5953 : _GEN_5857; // @[executor.scala 290:56]
  wire [7:0] _GEN_6050 = 8'h5 < length_3 ? _GEN_5954 : _GEN_5858; // @[executor.scala 290:56]
  wire [7:0] field_byte_30 = field_3[15:8]; // @[executor.scala 287:53]
  wire [7:0] total_offset_30 = offset_3 + 8'h6; // @[executor.scala 289:53]
  wire [7:0] _GEN_6051 = 7'h0 == total_offset_30[6:0] ? field_byte_30 : _GEN_5955; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6052 = 7'h1 == total_offset_30[6:0] ? field_byte_30 : _GEN_5956; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6053 = 7'h2 == total_offset_30[6:0] ? field_byte_30 : _GEN_5957; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6054 = 7'h3 == total_offset_30[6:0] ? field_byte_30 : _GEN_5958; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6055 = 7'h4 == total_offset_30[6:0] ? field_byte_30 : _GEN_5959; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6056 = 7'h5 == total_offset_30[6:0] ? field_byte_30 : _GEN_5960; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6057 = 7'h6 == total_offset_30[6:0] ? field_byte_30 : _GEN_5961; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6058 = 7'h7 == total_offset_30[6:0] ? field_byte_30 : _GEN_5962; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6059 = 7'h8 == total_offset_30[6:0] ? field_byte_30 : _GEN_5963; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6060 = 7'h9 == total_offset_30[6:0] ? field_byte_30 : _GEN_5964; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6061 = 7'ha == total_offset_30[6:0] ? field_byte_30 : _GEN_5965; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6062 = 7'hb == total_offset_30[6:0] ? field_byte_30 : _GEN_5966; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6063 = 7'hc == total_offset_30[6:0] ? field_byte_30 : _GEN_5967; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6064 = 7'hd == total_offset_30[6:0] ? field_byte_30 : _GEN_5968; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6065 = 7'he == total_offset_30[6:0] ? field_byte_30 : _GEN_5969; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6066 = 7'hf == total_offset_30[6:0] ? field_byte_30 : _GEN_5970; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6067 = 7'h10 == total_offset_30[6:0] ? field_byte_30 : _GEN_5971; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6068 = 7'h11 == total_offset_30[6:0] ? field_byte_30 : _GEN_5972; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6069 = 7'h12 == total_offset_30[6:0] ? field_byte_30 : _GEN_5973; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6070 = 7'h13 == total_offset_30[6:0] ? field_byte_30 : _GEN_5974; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6071 = 7'h14 == total_offset_30[6:0] ? field_byte_30 : _GEN_5975; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6072 = 7'h15 == total_offset_30[6:0] ? field_byte_30 : _GEN_5976; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6073 = 7'h16 == total_offset_30[6:0] ? field_byte_30 : _GEN_5977; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6074 = 7'h17 == total_offset_30[6:0] ? field_byte_30 : _GEN_5978; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6075 = 7'h18 == total_offset_30[6:0] ? field_byte_30 : _GEN_5979; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6076 = 7'h19 == total_offset_30[6:0] ? field_byte_30 : _GEN_5980; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6077 = 7'h1a == total_offset_30[6:0] ? field_byte_30 : _GEN_5981; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6078 = 7'h1b == total_offset_30[6:0] ? field_byte_30 : _GEN_5982; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6079 = 7'h1c == total_offset_30[6:0] ? field_byte_30 : _GEN_5983; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6080 = 7'h1d == total_offset_30[6:0] ? field_byte_30 : _GEN_5984; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6081 = 7'h1e == total_offset_30[6:0] ? field_byte_30 : _GEN_5985; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6082 = 7'h1f == total_offset_30[6:0] ? field_byte_30 : _GEN_5986; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6083 = 7'h20 == total_offset_30[6:0] ? field_byte_30 : _GEN_5987; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6084 = 7'h21 == total_offset_30[6:0] ? field_byte_30 : _GEN_5988; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6085 = 7'h22 == total_offset_30[6:0] ? field_byte_30 : _GEN_5989; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6086 = 7'h23 == total_offset_30[6:0] ? field_byte_30 : _GEN_5990; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6087 = 7'h24 == total_offset_30[6:0] ? field_byte_30 : _GEN_5991; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6088 = 7'h25 == total_offset_30[6:0] ? field_byte_30 : _GEN_5992; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6089 = 7'h26 == total_offset_30[6:0] ? field_byte_30 : _GEN_5993; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6090 = 7'h27 == total_offset_30[6:0] ? field_byte_30 : _GEN_5994; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6091 = 7'h28 == total_offset_30[6:0] ? field_byte_30 : _GEN_5995; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6092 = 7'h29 == total_offset_30[6:0] ? field_byte_30 : _GEN_5996; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6093 = 7'h2a == total_offset_30[6:0] ? field_byte_30 : _GEN_5997; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6094 = 7'h2b == total_offset_30[6:0] ? field_byte_30 : _GEN_5998; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6095 = 7'h2c == total_offset_30[6:0] ? field_byte_30 : _GEN_5999; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6096 = 7'h2d == total_offset_30[6:0] ? field_byte_30 : _GEN_6000; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6097 = 7'h2e == total_offset_30[6:0] ? field_byte_30 : _GEN_6001; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6098 = 7'h2f == total_offset_30[6:0] ? field_byte_30 : _GEN_6002; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6099 = 7'h30 == total_offset_30[6:0] ? field_byte_30 : _GEN_6003; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6100 = 7'h31 == total_offset_30[6:0] ? field_byte_30 : _GEN_6004; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6101 = 7'h32 == total_offset_30[6:0] ? field_byte_30 : _GEN_6005; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6102 = 7'h33 == total_offset_30[6:0] ? field_byte_30 : _GEN_6006; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6103 = 7'h34 == total_offset_30[6:0] ? field_byte_30 : _GEN_6007; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6104 = 7'h35 == total_offset_30[6:0] ? field_byte_30 : _GEN_6008; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6105 = 7'h36 == total_offset_30[6:0] ? field_byte_30 : _GEN_6009; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6106 = 7'h37 == total_offset_30[6:0] ? field_byte_30 : _GEN_6010; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6107 = 7'h38 == total_offset_30[6:0] ? field_byte_30 : _GEN_6011; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6108 = 7'h39 == total_offset_30[6:0] ? field_byte_30 : _GEN_6012; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6109 = 7'h3a == total_offset_30[6:0] ? field_byte_30 : _GEN_6013; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6110 = 7'h3b == total_offset_30[6:0] ? field_byte_30 : _GEN_6014; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6111 = 7'h3c == total_offset_30[6:0] ? field_byte_30 : _GEN_6015; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6112 = 7'h3d == total_offset_30[6:0] ? field_byte_30 : _GEN_6016; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6113 = 7'h3e == total_offset_30[6:0] ? field_byte_30 : _GEN_6017; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6114 = 7'h3f == total_offset_30[6:0] ? field_byte_30 : _GEN_6018; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6115 = 7'h40 == total_offset_30[6:0] ? field_byte_30 : _GEN_6019; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6116 = 7'h41 == total_offset_30[6:0] ? field_byte_30 : _GEN_6020; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6117 = 7'h42 == total_offset_30[6:0] ? field_byte_30 : _GEN_6021; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6118 = 7'h43 == total_offset_30[6:0] ? field_byte_30 : _GEN_6022; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6119 = 7'h44 == total_offset_30[6:0] ? field_byte_30 : _GEN_6023; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6120 = 7'h45 == total_offset_30[6:0] ? field_byte_30 : _GEN_6024; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6121 = 7'h46 == total_offset_30[6:0] ? field_byte_30 : _GEN_6025; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6122 = 7'h47 == total_offset_30[6:0] ? field_byte_30 : _GEN_6026; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6123 = 7'h48 == total_offset_30[6:0] ? field_byte_30 : _GEN_6027; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6124 = 7'h49 == total_offset_30[6:0] ? field_byte_30 : _GEN_6028; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6125 = 7'h4a == total_offset_30[6:0] ? field_byte_30 : _GEN_6029; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6126 = 7'h4b == total_offset_30[6:0] ? field_byte_30 : _GEN_6030; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6127 = 7'h4c == total_offset_30[6:0] ? field_byte_30 : _GEN_6031; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6128 = 7'h4d == total_offset_30[6:0] ? field_byte_30 : _GEN_6032; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6129 = 7'h4e == total_offset_30[6:0] ? field_byte_30 : _GEN_6033; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6130 = 7'h4f == total_offset_30[6:0] ? field_byte_30 : _GEN_6034; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6131 = 7'h50 == total_offset_30[6:0] ? field_byte_30 : _GEN_6035; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6132 = 7'h51 == total_offset_30[6:0] ? field_byte_30 : _GEN_6036; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6133 = 7'h52 == total_offset_30[6:0] ? field_byte_30 : _GEN_6037; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6134 = 7'h53 == total_offset_30[6:0] ? field_byte_30 : _GEN_6038; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6135 = 7'h54 == total_offset_30[6:0] ? field_byte_30 : _GEN_6039; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6136 = 7'h55 == total_offset_30[6:0] ? field_byte_30 : _GEN_6040; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6137 = 7'h56 == total_offset_30[6:0] ? field_byte_30 : _GEN_6041; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6138 = 7'h57 == total_offset_30[6:0] ? field_byte_30 : _GEN_6042; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6139 = 7'h58 == total_offset_30[6:0] ? field_byte_30 : _GEN_6043; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6140 = 7'h59 == total_offset_30[6:0] ? field_byte_30 : _GEN_6044; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6141 = 7'h5a == total_offset_30[6:0] ? field_byte_30 : _GEN_6045; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6142 = 7'h5b == total_offset_30[6:0] ? field_byte_30 : _GEN_6046; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6143 = 7'h5c == total_offset_30[6:0] ? field_byte_30 : _GEN_6047; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6144 = 7'h5d == total_offset_30[6:0] ? field_byte_30 : _GEN_6048; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6145 = 7'h5e == total_offset_30[6:0] ? field_byte_30 : _GEN_6049; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6146 = 7'h5f == total_offset_30[6:0] ? field_byte_30 : _GEN_6050; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6147 = 8'h6 < length_3 ? _GEN_6051 : _GEN_5955; // @[executor.scala 290:56]
  wire [7:0] _GEN_6148 = 8'h6 < length_3 ? _GEN_6052 : _GEN_5956; // @[executor.scala 290:56]
  wire [7:0] _GEN_6149 = 8'h6 < length_3 ? _GEN_6053 : _GEN_5957; // @[executor.scala 290:56]
  wire [7:0] _GEN_6150 = 8'h6 < length_3 ? _GEN_6054 : _GEN_5958; // @[executor.scala 290:56]
  wire [7:0] _GEN_6151 = 8'h6 < length_3 ? _GEN_6055 : _GEN_5959; // @[executor.scala 290:56]
  wire [7:0] _GEN_6152 = 8'h6 < length_3 ? _GEN_6056 : _GEN_5960; // @[executor.scala 290:56]
  wire [7:0] _GEN_6153 = 8'h6 < length_3 ? _GEN_6057 : _GEN_5961; // @[executor.scala 290:56]
  wire [7:0] _GEN_6154 = 8'h6 < length_3 ? _GEN_6058 : _GEN_5962; // @[executor.scala 290:56]
  wire [7:0] _GEN_6155 = 8'h6 < length_3 ? _GEN_6059 : _GEN_5963; // @[executor.scala 290:56]
  wire [7:0] _GEN_6156 = 8'h6 < length_3 ? _GEN_6060 : _GEN_5964; // @[executor.scala 290:56]
  wire [7:0] _GEN_6157 = 8'h6 < length_3 ? _GEN_6061 : _GEN_5965; // @[executor.scala 290:56]
  wire [7:0] _GEN_6158 = 8'h6 < length_3 ? _GEN_6062 : _GEN_5966; // @[executor.scala 290:56]
  wire [7:0] _GEN_6159 = 8'h6 < length_3 ? _GEN_6063 : _GEN_5967; // @[executor.scala 290:56]
  wire [7:0] _GEN_6160 = 8'h6 < length_3 ? _GEN_6064 : _GEN_5968; // @[executor.scala 290:56]
  wire [7:0] _GEN_6161 = 8'h6 < length_3 ? _GEN_6065 : _GEN_5969; // @[executor.scala 290:56]
  wire [7:0] _GEN_6162 = 8'h6 < length_3 ? _GEN_6066 : _GEN_5970; // @[executor.scala 290:56]
  wire [7:0] _GEN_6163 = 8'h6 < length_3 ? _GEN_6067 : _GEN_5971; // @[executor.scala 290:56]
  wire [7:0] _GEN_6164 = 8'h6 < length_3 ? _GEN_6068 : _GEN_5972; // @[executor.scala 290:56]
  wire [7:0] _GEN_6165 = 8'h6 < length_3 ? _GEN_6069 : _GEN_5973; // @[executor.scala 290:56]
  wire [7:0] _GEN_6166 = 8'h6 < length_3 ? _GEN_6070 : _GEN_5974; // @[executor.scala 290:56]
  wire [7:0] _GEN_6167 = 8'h6 < length_3 ? _GEN_6071 : _GEN_5975; // @[executor.scala 290:56]
  wire [7:0] _GEN_6168 = 8'h6 < length_3 ? _GEN_6072 : _GEN_5976; // @[executor.scala 290:56]
  wire [7:0] _GEN_6169 = 8'h6 < length_3 ? _GEN_6073 : _GEN_5977; // @[executor.scala 290:56]
  wire [7:0] _GEN_6170 = 8'h6 < length_3 ? _GEN_6074 : _GEN_5978; // @[executor.scala 290:56]
  wire [7:0] _GEN_6171 = 8'h6 < length_3 ? _GEN_6075 : _GEN_5979; // @[executor.scala 290:56]
  wire [7:0] _GEN_6172 = 8'h6 < length_3 ? _GEN_6076 : _GEN_5980; // @[executor.scala 290:56]
  wire [7:0] _GEN_6173 = 8'h6 < length_3 ? _GEN_6077 : _GEN_5981; // @[executor.scala 290:56]
  wire [7:0] _GEN_6174 = 8'h6 < length_3 ? _GEN_6078 : _GEN_5982; // @[executor.scala 290:56]
  wire [7:0] _GEN_6175 = 8'h6 < length_3 ? _GEN_6079 : _GEN_5983; // @[executor.scala 290:56]
  wire [7:0] _GEN_6176 = 8'h6 < length_3 ? _GEN_6080 : _GEN_5984; // @[executor.scala 290:56]
  wire [7:0] _GEN_6177 = 8'h6 < length_3 ? _GEN_6081 : _GEN_5985; // @[executor.scala 290:56]
  wire [7:0] _GEN_6178 = 8'h6 < length_3 ? _GEN_6082 : _GEN_5986; // @[executor.scala 290:56]
  wire [7:0] _GEN_6179 = 8'h6 < length_3 ? _GEN_6083 : _GEN_5987; // @[executor.scala 290:56]
  wire [7:0] _GEN_6180 = 8'h6 < length_3 ? _GEN_6084 : _GEN_5988; // @[executor.scala 290:56]
  wire [7:0] _GEN_6181 = 8'h6 < length_3 ? _GEN_6085 : _GEN_5989; // @[executor.scala 290:56]
  wire [7:0] _GEN_6182 = 8'h6 < length_3 ? _GEN_6086 : _GEN_5990; // @[executor.scala 290:56]
  wire [7:0] _GEN_6183 = 8'h6 < length_3 ? _GEN_6087 : _GEN_5991; // @[executor.scala 290:56]
  wire [7:0] _GEN_6184 = 8'h6 < length_3 ? _GEN_6088 : _GEN_5992; // @[executor.scala 290:56]
  wire [7:0] _GEN_6185 = 8'h6 < length_3 ? _GEN_6089 : _GEN_5993; // @[executor.scala 290:56]
  wire [7:0] _GEN_6186 = 8'h6 < length_3 ? _GEN_6090 : _GEN_5994; // @[executor.scala 290:56]
  wire [7:0] _GEN_6187 = 8'h6 < length_3 ? _GEN_6091 : _GEN_5995; // @[executor.scala 290:56]
  wire [7:0] _GEN_6188 = 8'h6 < length_3 ? _GEN_6092 : _GEN_5996; // @[executor.scala 290:56]
  wire [7:0] _GEN_6189 = 8'h6 < length_3 ? _GEN_6093 : _GEN_5997; // @[executor.scala 290:56]
  wire [7:0] _GEN_6190 = 8'h6 < length_3 ? _GEN_6094 : _GEN_5998; // @[executor.scala 290:56]
  wire [7:0] _GEN_6191 = 8'h6 < length_3 ? _GEN_6095 : _GEN_5999; // @[executor.scala 290:56]
  wire [7:0] _GEN_6192 = 8'h6 < length_3 ? _GEN_6096 : _GEN_6000; // @[executor.scala 290:56]
  wire [7:0] _GEN_6193 = 8'h6 < length_3 ? _GEN_6097 : _GEN_6001; // @[executor.scala 290:56]
  wire [7:0] _GEN_6194 = 8'h6 < length_3 ? _GEN_6098 : _GEN_6002; // @[executor.scala 290:56]
  wire [7:0] _GEN_6195 = 8'h6 < length_3 ? _GEN_6099 : _GEN_6003; // @[executor.scala 290:56]
  wire [7:0] _GEN_6196 = 8'h6 < length_3 ? _GEN_6100 : _GEN_6004; // @[executor.scala 290:56]
  wire [7:0] _GEN_6197 = 8'h6 < length_3 ? _GEN_6101 : _GEN_6005; // @[executor.scala 290:56]
  wire [7:0] _GEN_6198 = 8'h6 < length_3 ? _GEN_6102 : _GEN_6006; // @[executor.scala 290:56]
  wire [7:0] _GEN_6199 = 8'h6 < length_3 ? _GEN_6103 : _GEN_6007; // @[executor.scala 290:56]
  wire [7:0] _GEN_6200 = 8'h6 < length_3 ? _GEN_6104 : _GEN_6008; // @[executor.scala 290:56]
  wire [7:0] _GEN_6201 = 8'h6 < length_3 ? _GEN_6105 : _GEN_6009; // @[executor.scala 290:56]
  wire [7:0] _GEN_6202 = 8'h6 < length_3 ? _GEN_6106 : _GEN_6010; // @[executor.scala 290:56]
  wire [7:0] _GEN_6203 = 8'h6 < length_3 ? _GEN_6107 : _GEN_6011; // @[executor.scala 290:56]
  wire [7:0] _GEN_6204 = 8'h6 < length_3 ? _GEN_6108 : _GEN_6012; // @[executor.scala 290:56]
  wire [7:0] _GEN_6205 = 8'h6 < length_3 ? _GEN_6109 : _GEN_6013; // @[executor.scala 290:56]
  wire [7:0] _GEN_6206 = 8'h6 < length_3 ? _GEN_6110 : _GEN_6014; // @[executor.scala 290:56]
  wire [7:0] _GEN_6207 = 8'h6 < length_3 ? _GEN_6111 : _GEN_6015; // @[executor.scala 290:56]
  wire [7:0] _GEN_6208 = 8'h6 < length_3 ? _GEN_6112 : _GEN_6016; // @[executor.scala 290:56]
  wire [7:0] _GEN_6209 = 8'h6 < length_3 ? _GEN_6113 : _GEN_6017; // @[executor.scala 290:56]
  wire [7:0] _GEN_6210 = 8'h6 < length_3 ? _GEN_6114 : _GEN_6018; // @[executor.scala 290:56]
  wire [7:0] _GEN_6211 = 8'h6 < length_3 ? _GEN_6115 : _GEN_6019; // @[executor.scala 290:56]
  wire [7:0] _GEN_6212 = 8'h6 < length_3 ? _GEN_6116 : _GEN_6020; // @[executor.scala 290:56]
  wire [7:0] _GEN_6213 = 8'h6 < length_3 ? _GEN_6117 : _GEN_6021; // @[executor.scala 290:56]
  wire [7:0] _GEN_6214 = 8'h6 < length_3 ? _GEN_6118 : _GEN_6022; // @[executor.scala 290:56]
  wire [7:0] _GEN_6215 = 8'h6 < length_3 ? _GEN_6119 : _GEN_6023; // @[executor.scala 290:56]
  wire [7:0] _GEN_6216 = 8'h6 < length_3 ? _GEN_6120 : _GEN_6024; // @[executor.scala 290:56]
  wire [7:0] _GEN_6217 = 8'h6 < length_3 ? _GEN_6121 : _GEN_6025; // @[executor.scala 290:56]
  wire [7:0] _GEN_6218 = 8'h6 < length_3 ? _GEN_6122 : _GEN_6026; // @[executor.scala 290:56]
  wire [7:0] _GEN_6219 = 8'h6 < length_3 ? _GEN_6123 : _GEN_6027; // @[executor.scala 290:56]
  wire [7:0] _GEN_6220 = 8'h6 < length_3 ? _GEN_6124 : _GEN_6028; // @[executor.scala 290:56]
  wire [7:0] _GEN_6221 = 8'h6 < length_3 ? _GEN_6125 : _GEN_6029; // @[executor.scala 290:56]
  wire [7:0] _GEN_6222 = 8'h6 < length_3 ? _GEN_6126 : _GEN_6030; // @[executor.scala 290:56]
  wire [7:0] _GEN_6223 = 8'h6 < length_3 ? _GEN_6127 : _GEN_6031; // @[executor.scala 290:56]
  wire [7:0] _GEN_6224 = 8'h6 < length_3 ? _GEN_6128 : _GEN_6032; // @[executor.scala 290:56]
  wire [7:0] _GEN_6225 = 8'h6 < length_3 ? _GEN_6129 : _GEN_6033; // @[executor.scala 290:56]
  wire [7:0] _GEN_6226 = 8'h6 < length_3 ? _GEN_6130 : _GEN_6034; // @[executor.scala 290:56]
  wire [7:0] _GEN_6227 = 8'h6 < length_3 ? _GEN_6131 : _GEN_6035; // @[executor.scala 290:56]
  wire [7:0] _GEN_6228 = 8'h6 < length_3 ? _GEN_6132 : _GEN_6036; // @[executor.scala 290:56]
  wire [7:0] _GEN_6229 = 8'h6 < length_3 ? _GEN_6133 : _GEN_6037; // @[executor.scala 290:56]
  wire [7:0] _GEN_6230 = 8'h6 < length_3 ? _GEN_6134 : _GEN_6038; // @[executor.scala 290:56]
  wire [7:0] _GEN_6231 = 8'h6 < length_3 ? _GEN_6135 : _GEN_6039; // @[executor.scala 290:56]
  wire [7:0] _GEN_6232 = 8'h6 < length_3 ? _GEN_6136 : _GEN_6040; // @[executor.scala 290:56]
  wire [7:0] _GEN_6233 = 8'h6 < length_3 ? _GEN_6137 : _GEN_6041; // @[executor.scala 290:56]
  wire [7:0] _GEN_6234 = 8'h6 < length_3 ? _GEN_6138 : _GEN_6042; // @[executor.scala 290:56]
  wire [7:0] _GEN_6235 = 8'h6 < length_3 ? _GEN_6139 : _GEN_6043; // @[executor.scala 290:56]
  wire [7:0] _GEN_6236 = 8'h6 < length_3 ? _GEN_6140 : _GEN_6044; // @[executor.scala 290:56]
  wire [7:0] _GEN_6237 = 8'h6 < length_3 ? _GEN_6141 : _GEN_6045; // @[executor.scala 290:56]
  wire [7:0] _GEN_6238 = 8'h6 < length_3 ? _GEN_6142 : _GEN_6046; // @[executor.scala 290:56]
  wire [7:0] _GEN_6239 = 8'h6 < length_3 ? _GEN_6143 : _GEN_6047; // @[executor.scala 290:56]
  wire [7:0] _GEN_6240 = 8'h6 < length_3 ? _GEN_6144 : _GEN_6048; // @[executor.scala 290:56]
  wire [7:0] _GEN_6241 = 8'h6 < length_3 ? _GEN_6145 : _GEN_6049; // @[executor.scala 290:56]
  wire [7:0] _GEN_6242 = 8'h6 < length_3 ? _GEN_6146 : _GEN_6050; // @[executor.scala 290:56]
  wire [7:0] field_byte_31 = field_3[7:0]; // @[executor.scala 287:53]
  wire [7:0] total_offset_31 = offset_3 + 8'h7; // @[executor.scala 289:53]
  wire [7:0] _GEN_6243 = 7'h0 == total_offset_31[6:0] ? field_byte_31 : _GEN_6147; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6244 = 7'h1 == total_offset_31[6:0] ? field_byte_31 : _GEN_6148; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6245 = 7'h2 == total_offset_31[6:0] ? field_byte_31 : _GEN_6149; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6246 = 7'h3 == total_offset_31[6:0] ? field_byte_31 : _GEN_6150; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6247 = 7'h4 == total_offset_31[6:0] ? field_byte_31 : _GEN_6151; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6248 = 7'h5 == total_offset_31[6:0] ? field_byte_31 : _GEN_6152; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6249 = 7'h6 == total_offset_31[6:0] ? field_byte_31 : _GEN_6153; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6250 = 7'h7 == total_offset_31[6:0] ? field_byte_31 : _GEN_6154; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6251 = 7'h8 == total_offset_31[6:0] ? field_byte_31 : _GEN_6155; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6252 = 7'h9 == total_offset_31[6:0] ? field_byte_31 : _GEN_6156; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6253 = 7'ha == total_offset_31[6:0] ? field_byte_31 : _GEN_6157; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6254 = 7'hb == total_offset_31[6:0] ? field_byte_31 : _GEN_6158; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6255 = 7'hc == total_offset_31[6:0] ? field_byte_31 : _GEN_6159; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6256 = 7'hd == total_offset_31[6:0] ? field_byte_31 : _GEN_6160; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6257 = 7'he == total_offset_31[6:0] ? field_byte_31 : _GEN_6161; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6258 = 7'hf == total_offset_31[6:0] ? field_byte_31 : _GEN_6162; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6259 = 7'h10 == total_offset_31[6:0] ? field_byte_31 : _GEN_6163; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6260 = 7'h11 == total_offset_31[6:0] ? field_byte_31 : _GEN_6164; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6261 = 7'h12 == total_offset_31[6:0] ? field_byte_31 : _GEN_6165; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6262 = 7'h13 == total_offset_31[6:0] ? field_byte_31 : _GEN_6166; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6263 = 7'h14 == total_offset_31[6:0] ? field_byte_31 : _GEN_6167; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6264 = 7'h15 == total_offset_31[6:0] ? field_byte_31 : _GEN_6168; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6265 = 7'h16 == total_offset_31[6:0] ? field_byte_31 : _GEN_6169; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6266 = 7'h17 == total_offset_31[6:0] ? field_byte_31 : _GEN_6170; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6267 = 7'h18 == total_offset_31[6:0] ? field_byte_31 : _GEN_6171; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6268 = 7'h19 == total_offset_31[6:0] ? field_byte_31 : _GEN_6172; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6269 = 7'h1a == total_offset_31[6:0] ? field_byte_31 : _GEN_6173; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6270 = 7'h1b == total_offset_31[6:0] ? field_byte_31 : _GEN_6174; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6271 = 7'h1c == total_offset_31[6:0] ? field_byte_31 : _GEN_6175; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6272 = 7'h1d == total_offset_31[6:0] ? field_byte_31 : _GEN_6176; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6273 = 7'h1e == total_offset_31[6:0] ? field_byte_31 : _GEN_6177; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6274 = 7'h1f == total_offset_31[6:0] ? field_byte_31 : _GEN_6178; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6275 = 7'h20 == total_offset_31[6:0] ? field_byte_31 : _GEN_6179; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6276 = 7'h21 == total_offset_31[6:0] ? field_byte_31 : _GEN_6180; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6277 = 7'h22 == total_offset_31[6:0] ? field_byte_31 : _GEN_6181; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6278 = 7'h23 == total_offset_31[6:0] ? field_byte_31 : _GEN_6182; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6279 = 7'h24 == total_offset_31[6:0] ? field_byte_31 : _GEN_6183; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6280 = 7'h25 == total_offset_31[6:0] ? field_byte_31 : _GEN_6184; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6281 = 7'h26 == total_offset_31[6:0] ? field_byte_31 : _GEN_6185; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6282 = 7'h27 == total_offset_31[6:0] ? field_byte_31 : _GEN_6186; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6283 = 7'h28 == total_offset_31[6:0] ? field_byte_31 : _GEN_6187; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6284 = 7'h29 == total_offset_31[6:0] ? field_byte_31 : _GEN_6188; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6285 = 7'h2a == total_offset_31[6:0] ? field_byte_31 : _GEN_6189; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6286 = 7'h2b == total_offset_31[6:0] ? field_byte_31 : _GEN_6190; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6287 = 7'h2c == total_offset_31[6:0] ? field_byte_31 : _GEN_6191; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6288 = 7'h2d == total_offset_31[6:0] ? field_byte_31 : _GEN_6192; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6289 = 7'h2e == total_offset_31[6:0] ? field_byte_31 : _GEN_6193; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6290 = 7'h2f == total_offset_31[6:0] ? field_byte_31 : _GEN_6194; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6291 = 7'h30 == total_offset_31[6:0] ? field_byte_31 : _GEN_6195; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6292 = 7'h31 == total_offset_31[6:0] ? field_byte_31 : _GEN_6196; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6293 = 7'h32 == total_offset_31[6:0] ? field_byte_31 : _GEN_6197; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6294 = 7'h33 == total_offset_31[6:0] ? field_byte_31 : _GEN_6198; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6295 = 7'h34 == total_offset_31[6:0] ? field_byte_31 : _GEN_6199; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6296 = 7'h35 == total_offset_31[6:0] ? field_byte_31 : _GEN_6200; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6297 = 7'h36 == total_offset_31[6:0] ? field_byte_31 : _GEN_6201; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6298 = 7'h37 == total_offset_31[6:0] ? field_byte_31 : _GEN_6202; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6299 = 7'h38 == total_offset_31[6:0] ? field_byte_31 : _GEN_6203; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6300 = 7'h39 == total_offset_31[6:0] ? field_byte_31 : _GEN_6204; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6301 = 7'h3a == total_offset_31[6:0] ? field_byte_31 : _GEN_6205; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6302 = 7'h3b == total_offset_31[6:0] ? field_byte_31 : _GEN_6206; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6303 = 7'h3c == total_offset_31[6:0] ? field_byte_31 : _GEN_6207; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6304 = 7'h3d == total_offset_31[6:0] ? field_byte_31 : _GEN_6208; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6305 = 7'h3e == total_offset_31[6:0] ? field_byte_31 : _GEN_6209; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6306 = 7'h3f == total_offset_31[6:0] ? field_byte_31 : _GEN_6210; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6307 = 7'h40 == total_offset_31[6:0] ? field_byte_31 : _GEN_6211; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6308 = 7'h41 == total_offset_31[6:0] ? field_byte_31 : _GEN_6212; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6309 = 7'h42 == total_offset_31[6:0] ? field_byte_31 : _GEN_6213; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6310 = 7'h43 == total_offset_31[6:0] ? field_byte_31 : _GEN_6214; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6311 = 7'h44 == total_offset_31[6:0] ? field_byte_31 : _GEN_6215; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6312 = 7'h45 == total_offset_31[6:0] ? field_byte_31 : _GEN_6216; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6313 = 7'h46 == total_offset_31[6:0] ? field_byte_31 : _GEN_6217; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6314 = 7'h47 == total_offset_31[6:0] ? field_byte_31 : _GEN_6218; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6315 = 7'h48 == total_offset_31[6:0] ? field_byte_31 : _GEN_6219; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6316 = 7'h49 == total_offset_31[6:0] ? field_byte_31 : _GEN_6220; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6317 = 7'h4a == total_offset_31[6:0] ? field_byte_31 : _GEN_6221; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6318 = 7'h4b == total_offset_31[6:0] ? field_byte_31 : _GEN_6222; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6319 = 7'h4c == total_offset_31[6:0] ? field_byte_31 : _GEN_6223; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6320 = 7'h4d == total_offset_31[6:0] ? field_byte_31 : _GEN_6224; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6321 = 7'h4e == total_offset_31[6:0] ? field_byte_31 : _GEN_6225; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6322 = 7'h4f == total_offset_31[6:0] ? field_byte_31 : _GEN_6226; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6323 = 7'h50 == total_offset_31[6:0] ? field_byte_31 : _GEN_6227; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6324 = 7'h51 == total_offset_31[6:0] ? field_byte_31 : _GEN_6228; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6325 = 7'h52 == total_offset_31[6:0] ? field_byte_31 : _GEN_6229; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6326 = 7'h53 == total_offset_31[6:0] ? field_byte_31 : _GEN_6230; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6327 = 7'h54 == total_offset_31[6:0] ? field_byte_31 : _GEN_6231; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6328 = 7'h55 == total_offset_31[6:0] ? field_byte_31 : _GEN_6232; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6329 = 7'h56 == total_offset_31[6:0] ? field_byte_31 : _GEN_6233; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6330 = 7'h57 == total_offset_31[6:0] ? field_byte_31 : _GEN_6234; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6331 = 7'h58 == total_offset_31[6:0] ? field_byte_31 : _GEN_6235; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6332 = 7'h59 == total_offset_31[6:0] ? field_byte_31 : _GEN_6236; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6333 = 7'h5a == total_offset_31[6:0] ? field_byte_31 : _GEN_6237; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6334 = 7'h5b == total_offset_31[6:0] ? field_byte_31 : _GEN_6238; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6335 = 7'h5c == total_offset_31[6:0] ? field_byte_31 : _GEN_6239; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6336 = 7'h5d == total_offset_31[6:0] ? field_byte_31 : _GEN_6240; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6337 = 7'h5e == total_offset_31[6:0] ? field_byte_31 : _GEN_6241; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6338 = 7'h5f == total_offset_31[6:0] ? field_byte_31 : _GEN_6242; // @[executor.scala 291:60 executor.scala 291:60]
  wire [7:0] _GEN_6339 = 8'h7 < length_3 ? _GEN_6243 : _GEN_6147; // @[executor.scala 290:56]
  wire [7:0] _GEN_6340 = 8'h7 < length_3 ? _GEN_6244 : _GEN_6148; // @[executor.scala 290:56]
  wire [7:0] _GEN_6341 = 8'h7 < length_3 ? _GEN_6245 : _GEN_6149; // @[executor.scala 290:56]
  wire [7:0] _GEN_6342 = 8'h7 < length_3 ? _GEN_6246 : _GEN_6150; // @[executor.scala 290:56]
  wire [7:0] _GEN_6343 = 8'h7 < length_3 ? _GEN_6247 : _GEN_6151; // @[executor.scala 290:56]
  wire [7:0] _GEN_6344 = 8'h7 < length_3 ? _GEN_6248 : _GEN_6152; // @[executor.scala 290:56]
  wire [7:0] _GEN_6345 = 8'h7 < length_3 ? _GEN_6249 : _GEN_6153; // @[executor.scala 290:56]
  wire [7:0] _GEN_6346 = 8'h7 < length_3 ? _GEN_6250 : _GEN_6154; // @[executor.scala 290:56]
  wire [7:0] _GEN_6347 = 8'h7 < length_3 ? _GEN_6251 : _GEN_6155; // @[executor.scala 290:56]
  wire [7:0] _GEN_6348 = 8'h7 < length_3 ? _GEN_6252 : _GEN_6156; // @[executor.scala 290:56]
  wire [7:0] _GEN_6349 = 8'h7 < length_3 ? _GEN_6253 : _GEN_6157; // @[executor.scala 290:56]
  wire [7:0] _GEN_6350 = 8'h7 < length_3 ? _GEN_6254 : _GEN_6158; // @[executor.scala 290:56]
  wire [7:0] _GEN_6351 = 8'h7 < length_3 ? _GEN_6255 : _GEN_6159; // @[executor.scala 290:56]
  wire [7:0] _GEN_6352 = 8'h7 < length_3 ? _GEN_6256 : _GEN_6160; // @[executor.scala 290:56]
  wire [7:0] _GEN_6353 = 8'h7 < length_3 ? _GEN_6257 : _GEN_6161; // @[executor.scala 290:56]
  wire [7:0] _GEN_6354 = 8'h7 < length_3 ? _GEN_6258 : _GEN_6162; // @[executor.scala 290:56]
  wire [7:0] _GEN_6355 = 8'h7 < length_3 ? _GEN_6259 : _GEN_6163; // @[executor.scala 290:56]
  wire [7:0] _GEN_6356 = 8'h7 < length_3 ? _GEN_6260 : _GEN_6164; // @[executor.scala 290:56]
  wire [7:0] _GEN_6357 = 8'h7 < length_3 ? _GEN_6261 : _GEN_6165; // @[executor.scala 290:56]
  wire [7:0] _GEN_6358 = 8'h7 < length_3 ? _GEN_6262 : _GEN_6166; // @[executor.scala 290:56]
  wire [7:0] _GEN_6359 = 8'h7 < length_3 ? _GEN_6263 : _GEN_6167; // @[executor.scala 290:56]
  wire [7:0] _GEN_6360 = 8'h7 < length_3 ? _GEN_6264 : _GEN_6168; // @[executor.scala 290:56]
  wire [7:0] _GEN_6361 = 8'h7 < length_3 ? _GEN_6265 : _GEN_6169; // @[executor.scala 290:56]
  wire [7:0] _GEN_6362 = 8'h7 < length_3 ? _GEN_6266 : _GEN_6170; // @[executor.scala 290:56]
  wire [7:0] _GEN_6363 = 8'h7 < length_3 ? _GEN_6267 : _GEN_6171; // @[executor.scala 290:56]
  wire [7:0] _GEN_6364 = 8'h7 < length_3 ? _GEN_6268 : _GEN_6172; // @[executor.scala 290:56]
  wire [7:0] _GEN_6365 = 8'h7 < length_3 ? _GEN_6269 : _GEN_6173; // @[executor.scala 290:56]
  wire [7:0] _GEN_6366 = 8'h7 < length_3 ? _GEN_6270 : _GEN_6174; // @[executor.scala 290:56]
  wire [7:0] _GEN_6367 = 8'h7 < length_3 ? _GEN_6271 : _GEN_6175; // @[executor.scala 290:56]
  wire [7:0] _GEN_6368 = 8'h7 < length_3 ? _GEN_6272 : _GEN_6176; // @[executor.scala 290:56]
  wire [7:0] _GEN_6369 = 8'h7 < length_3 ? _GEN_6273 : _GEN_6177; // @[executor.scala 290:56]
  wire [7:0] _GEN_6370 = 8'h7 < length_3 ? _GEN_6274 : _GEN_6178; // @[executor.scala 290:56]
  wire [7:0] _GEN_6371 = 8'h7 < length_3 ? _GEN_6275 : _GEN_6179; // @[executor.scala 290:56]
  wire [7:0] _GEN_6372 = 8'h7 < length_3 ? _GEN_6276 : _GEN_6180; // @[executor.scala 290:56]
  wire [7:0] _GEN_6373 = 8'h7 < length_3 ? _GEN_6277 : _GEN_6181; // @[executor.scala 290:56]
  wire [7:0] _GEN_6374 = 8'h7 < length_3 ? _GEN_6278 : _GEN_6182; // @[executor.scala 290:56]
  wire [7:0] _GEN_6375 = 8'h7 < length_3 ? _GEN_6279 : _GEN_6183; // @[executor.scala 290:56]
  wire [7:0] _GEN_6376 = 8'h7 < length_3 ? _GEN_6280 : _GEN_6184; // @[executor.scala 290:56]
  wire [7:0] _GEN_6377 = 8'h7 < length_3 ? _GEN_6281 : _GEN_6185; // @[executor.scala 290:56]
  wire [7:0] _GEN_6378 = 8'h7 < length_3 ? _GEN_6282 : _GEN_6186; // @[executor.scala 290:56]
  wire [7:0] _GEN_6379 = 8'h7 < length_3 ? _GEN_6283 : _GEN_6187; // @[executor.scala 290:56]
  wire [7:0] _GEN_6380 = 8'h7 < length_3 ? _GEN_6284 : _GEN_6188; // @[executor.scala 290:56]
  wire [7:0] _GEN_6381 = 8'h7 < length_3 ? _GEN_6285 : _GEN_6189; // @[executor.scala 290:56]
  wire [7:0] _GEN_6382 = 8'h7 < length_3 ? _GEN_6286 : _GEN_6190; // @[executor.scala 290:56]
  wire [7:0] _GEN_6383 = 8'h7 < length_3 ? _GEN_6287 : _GEN_6191; // @[executor.scala 290:56]
  wire [7:0] _GEN_6384 = 8'h7 < length_3 ? _GEN_6288 : _GEN_6192; // @[executor.scala 290:56]
  wire [7:0] _GEN_6385 = 8'h7 < length_3 ? _GEN_6289 : _GEN_6193; // @[executor.scala 290:56]
  wire [7:0] _GEN_6386 = 8'h7 < length_3 ? _GEN_6290 : _GEN_6194; // @[executor.scala 290:56]
  wire [7:0] _GEN_6387 = 8'h7 < length_3 ? _GEN_6291 : _GEN_6195; // @[executor.scala 290:56]
  wire [7:0] _GEN_6388 = 8'h7 < length_3 ? _GEN_6292 : _GEN_6196; // @[executor.scala 290:56]
  wire [7:0] _GEN_6389 = 8'h7 < length_3 ? _GEN_6293 : _GEN_6197; // @[executor.scala 290:56]
  wire [7:0] _GEN_6390 = 8'h7 < length_3 ? _GEN_6294 : _GEN_6198; // @[executor.scala 290:56]
  wire [7:0] _GEN_6391 = 8'h7 < length_3 ? _GEN_6295 : _GEN_6199; // @[executor.scala 290:56]
  wire [7:0] _GEN_6392 = 8'h7 < length_3 ? _GEN_6296 : _GEN_6200; // @[executor.scala 290:56]
  wire [7:0] _GEN_6393 = 8'h7 < length_3 ? _GEN_6297 : _GEN_6201; // @[executor.scala 290:56]
  wire [7:0] _GEN_6394 = 8'h7 < length_3 ? _GEN_6298 : _GEN_6202; // @[executor.scala 290:56]
  wire [7:0] _GEN_6395 = 8'h7 < length_3 ? _GEN_6299 : _GEN_6203; // @[executor.scala 290:56]
  wire [7:0] _GEN_6396 = 8'h7 < length_3 ? _GEN_6300 : _GEN_6204; // @[executor.scala 290:56]
  wire [7:0] _GEN_6397 = 8'h7 < length_3 ? _GEN_6301 : _GEN_6205; // @[executor.scala 290:56]
  wire [7:0] _GEN_6398 = 8'h7 < length_3 ? _GEN_6302 : _GEN_6206; // @[executor.scala 290:56]
  wire [7:0] _GEN_6399 = 8'h7 < length_3 ? _GEN_6303 : _GEN_6207; // @[executor.scala 290:56]
  wire [7:0] _GEN_6400 = 8'h7 < length_3 ? _GEN_6304 : _GEN_6208; // @[executor.scala 290:56]
  wire [7:0] _GEN_6401 = 8'h7 < length_3 ? _GEN_6305 : _GEN_6209; // @[executor.scala 290:56]
  wire [7:0] _GEN_6402 = 8'h7 < length_3 ? _GEN_6306 : _GEN_6210; // @[executor.scala 290:56]
  wire [7:0] _GEN_6403 = 8'h7 < length_3 ? _GEN_6307 : _GEN_6211; // @[executor.scala 290:56]
  wire [7:0] _GEN_6404 = 8'h7 < length_3 ? _GEN_6308 : _GEN_6212; // @[executor.scala 290:56]
  wire [7:0] _GEN_6405 = 8'h7 < length_3 ? _GEN_6309 : _GEN_6213; // @[executor.scala 290:56]
  wire [7:0] _GEN_6406 = 8'h7 < length_3 ? _GEN_6310 : _GEN_6214; // @[executor.scala 290:56]
  wire [7:0] _GEN_6407 = 8'h7 < length_3 ? _GEN_6311 : _GEN_6215; // @[executor.scala 290:56]
  wire [7:0] _GEN_6408 = 8'h7 < length_3 ? _GEN_6312 : _GEN_6216; // @[executor.scala 290:56]
  wire [7:0] _GEN_6409 = 8'h7 < length_3 ? _GEN_6313 : _GEN_6217; // @[executor.scala 290:56]
  wire [7:0] _GEN_6410 = 8'h7 < length_3 ? _GEN_6314 : _GEN_6218; // @[executor.scala 290:56]
  wire [7:0] _GEN_6411 = 8'h7 < length_3 ? _GEN_6315 : _GEN_6219; // @[executor.scala 290:56]
  wire [7:0] _GEN_6412 = 8'h7 < length_3 ? _GEN_6316 : _GEN_6220; // @[executor.scala 290:56]
  wire [7:0] _GEN_6413 = 8'h7 < length_3 ? _GEN_6317 : _GEN_6221; // @[executor.scala 290:56]
  wire [7:0] _GEN_6414 = 8'h7 < length_3 ? _GEN_6318 : _GEN_6222; // @[executor.scala 290:56]
  wire [7:0] _GEN_6415 = 8'h7 < length_3 ? _GEN_6319 : _GEN_6223; // @[executor.scala 290:56]
  wire [7:0] _GEN_6416 = 8'h7 < length_3 ? _GEN_6320 : _GEN_6224; // @[executor.scala 290:56]
  wire [7:0] _GEN_6417 = 8'h7 < length_3 ? _GEN_6321 : _GEN_6225; // @[executor.scala 290:56]
  wire [7:0] _GEN_6418 = 8'h7 < length_3 ? _GEN_6322 : _GEN_6226; // @[executor.scala 290:56]
  wire [7:0] _GEN_6419 = 8'h7 < length_3 ? _GEN_6323 : _GEN_6227; // @[executor.scala 290:56]
  wire [7:0] _GEN_6420 = 8'h7 < length_3 ? _GEN_6324 : _GEN_6228; // @[executor.scala 290:56]
  wire [7:0] _GEN_6421 = 8'h7 < length_3 ? _GEN_6325 : _GEN_6229; // @[executor.scala 290:56]
  wire [7:0] _GEN_6422 = 8'h7 < length_3 ? _GEN_6326 : _GEN_6230; // @[executor.scala 290:56]
  wire [7:0] _GEN_6423 = 8'h7 < length_3 ? _GEN_6327 : _GEN_6231; // @[executor.scala 290:56]
  wire [7:0] _GEN_6424 = 8'h7 < length_3 ? _GEN_6328 : _GEN_6232; // @[executor.scala 290:56]
  wire [7:0] _GEN_6425 = 8'h7 < length_3 ? _GEN_6329 : _GEN_6233; // @[executor.scala 290:56]
  wire [7:0] _GEN_6426 = 8'h7 < length_3 ? _GEN_6330 : _GEN_6234; // @[executor.scala 290:56]
  wire [7:0] _GEN_6427 = 8'h7 < length_3 ? _GEN_6331 : _GEN_6235; // @[executor.scala 290:56]
  wire [7:0] _GEN_6428 = 8'h7 < length_3 ? _GEN_6332 : _GEN_6236; // @[executor.scala 290:56]
  wire [7:0] _GEN_6429 = 8'h7 < length_3 ? _GEN_6333 : _GEN_6237; // @[executor.scala 290:56]
  wire [7:0] _GEN_6430 = 8'h7 < length_3 ? _GEN_6334 : _GEN_6238; // @[executor.scala 290:56]
  wire [7:0] _GEN_6431 = 8'h7 < length_3 ? _GEN_6335 : _GEN_6239; // @[executor.scala 290:56]
  wire [7:0] _GEN_6432 = 8'h7 < length_3 ? _GEN_6336 : _GEN_6240; // @[executor.scala 290:56]
  wire [7:0] _GEN_6433 = 8'h7 < length_3 ? _GEN_6337 : _GEN_6241; // @[executor.scala 290:56]
  wire [7:0] _GEN_6434 = 8'h7 < length_3 ? _GEN_6338 : _GEN_6242; // @[executor.scala 290:56]
  wire [63:0] _GEN_6435 = length_3 == 8'h0 ? field_3 : _GEN_4802; // @[executor.scala 283:67 executor.scala 284:51]
  assign io_pipe_phv_out_data_0 = length_3 == 8'h0 ? _GEN_4803 : _GEN_6339; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_1 = length_3 == 8'h0 ? _GEN_4804 : _GEN_6340; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_2 = length_3 == 8'h0 ? _GEN_4805 : _GEN_6341; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_3 = length_3 == 8'h0 ? _GEN_4806 : _GEN_6342; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_4 = length_3 == 8'h0 ? _GEN_4807 : _GEN_6343; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_5 = length_3 == 8'h0 ? _GEN_4808 : _GEN_6344; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_6 = length_3 == 8'h0 ? _GEN_4809 : _GEN_6345; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_7 = length_3 == 8'h0 ? _GEN_4810 : _GEN_6346; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_8 = length_3 == 8'h0 ? _GEN_4811 : _GEN_6347; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_9 = length_3 == 8'h0 ? _GEN_4812 : _GEN_6348; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_10 = length_3 == 8'h0 ? _GEN_4813 : _GEN_6349; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_11 = length_3 == 8'h0 ? _GEN_4814 : _GEN_6350; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_12 = length_3 == 8'h0 ? _GEN_4815 : _GEN_6351; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_13 = length_3 == 8'h0 ? _GEN_4816 : _GEN_6352; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_14 = length_3 == 8'h0 ? _GEN_4817 : _GEN_6353; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_15 = length_3 == 8'h0 ? _GEN_4818 : _GEN_6354; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_16 = length_3 == 8'h0 ? _GEN_4819 : _GEN_6355; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_17 = length_3 == 8'h0 ? _GEN_4820 : _GEN_6356; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_18 = length_3 == 8'h0 ? _GEN_4821 : _GEN_6357; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_19 = length_3 == 8'h0 ? _GEN_4822 : _GEN_6358; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_20 = length_3 == 8'h0 ? _GEN_4823 : _GEN_6359; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_21 = length_3 == 8'h0 ? _GEN_4824 : _GEN_6360; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_22 = length_3 == 8'h0 ? _GEN_4825 : _GEN_6361; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_23 = length_3 == 8'h0 ? _GEN_4826 : _GEN_6362; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_24 = length_3 == 8'h0 ? _GEN_4827 : _GEN_6363; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_25 = length_3 == 8'h0 ? _GEN_4828 : _GEN_6364; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_26 = length_3 == 8'h0 ? _GEN_4829 : _GEN_6365; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_27 = length_3 == 8'h0 ? _GEN_4830 : _GEN_6366; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_28 = length_3 == 8'h0 ? _GEN_4831 : _GEN_6367; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_29 = length_3 == 8'h0 ? _GEN_4832 : _GEN_6368; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_30 = length_3 == 8'h0 ? _GEN_4833 : _GEN_6369; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_31 = length_3 == 8'h0 ? _GEN_4834 : _GEN_6370; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_32 = length_3 == 8'h0 ? _GEN_4835 : _GEN_6371; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_33 = length_3 == 8'h0 ? _GEN_4836 : _GEN_6372; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_34 = length_3 == 8'h0 ? _GEN_4837 : _GEN_6373; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_35 = length_3 == 8'h0 ? _GEN_4838 : _GEN_6374; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_36 = length_3 == 8'h0 ? _GEN_4839 : _GEN_6375; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_37 = length_3 == 8'h0 ? _GEN_4840 : _GEN_6376; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_38 = length_3 == 8'h0 ? _GEN_4841 : _GEN_6377; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_39 = length_3 == 8'h0 ? _GEN_4842 : _GEN_6378; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_40 = length_3 == 8'h0 ? _GEN_4843 : _GEN_6379; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_41 = length_3 == 8'h0 ? _GEN_4844 : _GEN_6380; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_42 = length_3 == 8'h0 ? _GEN_4845 : _GEN_6381; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_43 = length_3 == 8'h0 ? _GEN_4846 : _GEN_6382; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_44 = length_3 == 8'h0 ? _GEN_4847 : _GEN_6383; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_45 = length_3 == 8'h0 ? _GEN_4848 : _GEN_6384; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_46 = length_3 == 8'h0 ? _GEN_4849 : _GEN_6385; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_47 = length_3 == 8'h0 ? _GEN_4850 : _GEN_6386; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_48 = length_3 == 8'h0 ? _GEN_4851 : _GEN_6387; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_49 = length_3 == 8'h0 ? _GEN_4852 : _GEN_6388; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_50 = length_3 == 8'h0 ? _GEN_4853 : _GEN_6389; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_51 = length_3 == 8'h0 ? _GEN_4854 : _GEN_6390; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_52 = length_3 == 8'h0 ? _GEN_4855 : _GEN_6391; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_53 = length_3 == 8'h0 ? _GEN_4856 : _GEN_6392; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_54 = length_3 == 8'h0 ? _GEN_4857 : _GEN_6393; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_55 = length_3 == 8'h0 ? _GEN_4858 : _GEN_6394; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_56 = length_3 == 8'h0 ? _GEN_4859 : _GEN_6395; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_57 = length_3 == 8'h0 ? _GEN_4860 : _GEN_6396; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_58 = length_3 == 8'h0 ? _GEN_4861 : _GEN_6397; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_59 = length_3 == 8'h0 ? _GEN_4862 : _GEN_6398; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_60 = length_3 == 8'h0 ? _GEN_4863 : _GEN_6399; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_61 = length_3 == 8'h0 ? _GEN_4864 : _GEN_6400; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_62 = length_3 == 8'h0 ? _GEN_4865 : _GEN_6401; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_63 = length_3 == 8'h0 ? _GEN_4866 : _GEN_6402; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_64 = length_3 == 8'h0 ? _GEN_4867 : _GEN_6403; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_65 = length_3 == 8'h0 ? _GEN_4868 : _GEN_6404; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_66 = length_3 == 8'h0 ? _GEN_4869 : _GEN_6405; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_67 = length_3 == 8'h0 ? _GEN_4870 : _GEN_6406; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_68 = length_3 == 8'h0 ? _GEN_4871 : _GEN_6407; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_69 = length_3 == 8'h0 ? _GEN_4872 : _GEN_6408; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_70 = length_3 == 8'h0 ? _GEN_4873 : _GEN_6409; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_71 = length_3 == 8'h0 ? _GEN_4874 : _GEN_6410; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_72 = length_3 == 8'h0 ? _GEN_4875 : _GEN_6411; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_73 = length_3 == 8'h0 ? _GEN_4876 : _GEN_6412; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_74 = length_3 == 8'h0 ? _GEN_4877 : _GEN_6413; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_75 = length_3 == 8'h0 ? _GEN_4878 : _GEN_6414; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_76 = length_3 == 8'h0 ? _GEN_4879 : _GEN_6415; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_77 = length_3 == 8'h0 ? _GEN_4880 : _GEN_6416; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_78 = length_3 == 8'h0 ? _GEN_4881 : _GEN_6417; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_79 = length_3 == 8'h0 ? _GEN_4882 : _GEN_6418; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_80 = length_3 == 8'h0 ? _GEN_4883 : _GEN_6419; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_81 = length_3 == 8'h0 ? _GEN_4884 : _GEN_6420; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_82 = length_3 == 8'h0 ? _GEN_4885 : _GEN_6421; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_83 = length_3 == 8'h0 ? _GEN_4886 : _GEN_6422; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_84 = length_3 == 8'h0 ? _GEN_4887 : _GEN_6423; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_85 = length_3 == 8'h0 ? _GEN_4888 : _GEN_6424; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_86 = length_3 == 8'h0 ? _GEN_4889 : _GEN_6425; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_87 = length_3 == 8'h0 ? _GEN_4890 : _GEN_6426; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_88 = length_3 == 8'h0 ? _GEN_4891 : _GEN_6427; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_89 = length_3 == 8'h0 ? _GEN_4892 : _GEN_6428; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_90 = length_3 == 8'h0 ? _GEN_4893 : _GEN_6429; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_91 = length_3 == 8'h0 ? _GEN_4894 : _GEN_6430; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_92 = length_3 == 8'h0 ? _GEN_4895 : _GEN_6431; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_93 = length_3 == 8'h0 ? _GEN_4896 : _GEN_6432; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_94 = length_3 == 8'h0 ? _GEN_4897 : _GEN_6433; // @[executor.scala 283:67]
  assign io_pipe_phv_out_data_95 = length_3 == 8'h0 ? _GEN_4898 : _GEN_6434; // @[executor.scala 283:67]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 270:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 270:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 270:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 270:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 270:25]
  assign io_pipe_phv_out_next_processor_id = _GEN_6435[1:0];
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 269:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 269:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 269:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 269:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 269:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 269:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 269:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 269:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 269:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 269:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 269:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 269:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 269:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 269:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 269:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 269:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 269:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 269:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 269:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 269:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 269:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 269:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 269:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 269:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 269:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 269:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 269:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 269:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 269:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 269:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 269:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 269:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 269:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 269:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 269:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 269:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 269:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 269:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 269:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 269:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 269:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 269:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 269:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 269:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 269:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 269:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 269:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 269:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 269:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 269:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 269:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 269:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 269:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 269:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 269:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 269:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 269:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 269:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 269:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 269:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 269:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 269:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 269:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 269:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 269:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 269:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 269:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 269:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 269:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 269:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 269:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 269:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 269:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 269:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 269:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 269:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 269:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 269:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 269:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 269:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 269:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 269:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 269:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 269:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 269:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 269:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 269:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 269:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 269:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 269:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 269:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 269:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 269:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 269:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 269:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 269:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 269:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 269:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 269:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 269:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 269:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 269:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 269:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 269:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 269:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 269:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 269:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 269:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 269:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 269:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 269:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 269:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 269:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 269:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 269:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 269:13]
    offset_0 <= io_offset_in_0; // @[executor.scala 275:16]
    offset_1 <= io_offset_in_1; // @[executor.scala 275:16]
    offset_2 <= io_offset_in_2; // @[executor.scala 275:16]
    offset_3 <= io_offset_in_3; // @[executor.scala 275:16]
    length_0 <= io_length_in_0; // @[executor.scala 276:16]
    length_1 <= io_length_in_1; // @[executor.scala 276:16]
    length_2 <= io_length_in_2; // @[executor.scala 276:16]
    length_3 <= io_length_in_3; // @[executor.scala 276:16]
    field_0 <= io_field_in_0; // @[executor.scala 277:16]
    field_1 <= io_field_in_1; // @[executor.scala 277:16]
    field_2 <= io_field_in_2; // @[executor.scala 277:16]
    field_3 <= io_field_in_3; // @[executor.scala 277:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_header_0 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  phv_header_1 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  phv_header_2 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  phv_header_3 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  phv_header_4 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  phv_header_5 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  phv_header_6 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  phv_header_7 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  phv_header_8 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  phv_header_9 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  phv_header_10 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  phv_header_11 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  phv_header_12 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  phv_header_13 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  phv_header_14 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  phv_header_15 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  offset_0 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  offset_1 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  offset_2 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  offset_3 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  length_0 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  length_1 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  length_2 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  length_3 = _RAND_123[7:0];
  _RAND_124 = {2{`RANDOM}};
  field_0 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  field_1 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  field_2 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  field_3 = _RAND_127[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Executor(
  input         clock,
  input         reset,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  input         io_hit,
  input  [63:0] io_match_value,
  input         io_action_mod_en,
  input  [7:0]  io_action_mod_addr,
  input  [63:0] io_action_mod_data_0,
  input  [63:0] io_action_mod_data_1
);
  wire  pipe1_clock; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[executor.scala 299:23]
  wire [1:0] pipe1_io_pipe_phv_in_next_processor_id; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 299:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 299:23]
  wire [1:0] pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 299:23]
  wire  pipe1_io_hit; // @[executor.scala 299:23]
  wire [63:0] pipe1_io_match_value; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_args_out_0; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_args_out_1; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_args_out_2; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_args_out_3; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_args_out_4; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_args_out_5; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_args_out_6; // @[executor.scala 299:23]
  wire [31:0] pipe1_io_vliw_out_0; // @[executor.scala 299:23]
  wire [31:0] pipe1_io_vliw_out_1; // @[executor.scala 299:23]
  wire [31:0] pipe1_io_vliw_out_2; // @[executor.scala 299:23]
  wire [31:0] pipe1_io_vliw_out_3; // @[executor.scala 299:23]
  wire  pipe1_io_action_mod_en; // @[executor.scala 299:23]
  wire [7:0] pipe1_io_action_mod_addr; // @[executor.scala 299:23]
  wire [63:0] pipe1_io_action_mod_data_0; // @[executor.scala 299:23]
  wire [63:0] pipe1_io_action_mod_data_1; // @[executor.scala 299:23]
  wire  pipe2_clock; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[executor.scala 300:23]
  wire [1:0] pipe2_io_pipe_phv_in_next_processor_id; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 300:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 300:23]
  wire [1:0] pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_in_0; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_in_1; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_in_2; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_in_3; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_in_4; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_in_5; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_in_6; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_in_0; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_in_1; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_in_2; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_in_3; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_out_0; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_out_1; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_out_2; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_out_3; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_out_4; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_out_5; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_args_out_6; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_out_0; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_out_1; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_out_2; // @[executor.scala 300:23]
  wire [31:0] pipe2_io_vliw_out_3; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_offset_out_0; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_offset_out_1; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_offset_out_2; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_offset_out_3; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_length_out_0; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_length_out_1; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_length_out_2; // @[executor.scala 300:23]
  wire [7:0] pipe2_io_length_out_3; // @[executor.scala 300:23]
  wire  pipe3_clock; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[executor.scala 301:23]
  wire [1:0] pipe3_io_pipe_phv_in_next_processor_id; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 301:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 301:23]
  wire [1:0] pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_args_in_0; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_args_in_1; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_args_in_2; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_args_in_3; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_args_in_4; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_args_in_5; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_args_in_6; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_in_0; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_in_1; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_in_2; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_in_3; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_offset_in_0; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_offset_in_1; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_offset_in_2; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_offset_in_3; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_length_in_0; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_length_in_1; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_length_in_2; // @[executor.scala 301:23]
  wire [7:0] pipe3_io_length_in_3; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_out_0; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_out_1; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_out_2; // @[executor.scala 301:23]
  wire [31:0] pipe3_io_vliw_out_3; // @[executor.scala 301:23]
  wire [63:0] pipe3_io_field_out_0; // @[executor.scala 301:23]
  wire [63:0] pipe3_io_field_out_1; // @[executor.scala 301:23]
  wire [63:0] pipe3_io_field_out_2; // @[executor.scala 301:23]
  wire [63:0] pipe3_io_field_out_3; // @[executor.scala 301:23]
  wire  pipe4_clock; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[executor.scala 302:23]
  wire [1:0] pipe4_io_pipe_phv_in_next_processor_id; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 302:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 302:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 302:23]
  wire [1:0] pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_in_0; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_in_1; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_in_2; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_in_3; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_in_0; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_in_1; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_in_2; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_in_3; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_out_0; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_out_1; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_out_2; // @[executor.scala 302:23]
  wire [31:0] pipe4_io_vliw_out_3; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_out_0; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_out_1; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_out_2; // @[executor.scala 302:23]
  wire [63:0] pipe4_io_field_out_3; // @[executor.scala 302:23]
  wire  pipe5_clock; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[executor.scala 303:23]
  wire [1:0] pipe5_io_pipe_phv_in_next_processor_id; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 303:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 303:23]
  wire [1:0] pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 303:23]
  wire [31:0] pipe5_io_vliw_in_0; // @[executor.scala 303:23]
  wire [31:0] pipe5_io_vliw_in_1; // @[executor.scala 303:23]
  wire [31:0] pipe5_io_vliw_in_2; // @[executor.scala 303:23]
  wire [31:0] pipe5_io_vliw_in_3; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_in_0; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_in_1; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_in_2; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_in_3; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_offset_out_0; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_offset_out_1; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_offset_out_2; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_offset_out_3; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_length_out_0; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_length_out_1; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_length_out_2; // @[executor.scala 303:23]
  wire [7:0] pipe5_io_length_out_3; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_out_0; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_out_1; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_out_2; // @[executor.scala 303:23]
  wire [63:0] pipe5_io_field_out_3; // @[executor.scala 303:23]
  wire  pipe6_clock; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[executor.scala 304:23]
  wire [1:0] pipe6_io_pipe_phv_in_next_processor_id; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 304:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 304:23]
  wire [1:0] pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_offset_in_0; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_offset_in_1; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_offset_in_2; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_offset_in_3; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_length_in_0; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_length_in_1; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_length_in_2; // @[executor.scala 304:23]
  wire [7:0] pipe6_io_length_in_3; // @[executor.scala 304:23]
  wire [63:0] pipe6_io_field_in_0; // @[executor.scala 304:23]
  wire [63:0] pipe6_io_field_in_1; // @[executor.scala 304:23]
  wire [63:0] pipe6_io_field_in_2; // @[executor.scala 304:23]
  wire [63:0] pipe6_io_field_in_3; // @[executor.scala 304:23]
  ActionReader pipe1 ( // @[executor.scala 299:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_hit(pipe1_io_hit),
    .io_match_value(pipe1_io_match_value),
    .io_args_out_0(pipe1_io_args_out_0),
    .io_args_out_1(pipe1_io_args_out_1),
    .io_args_out_2(pipe1_io_args_out_2),
    .io_args_out_3(pipe1_io_args_out_3),
    .io_args_out_4(pipe1_io_args_out_4),
    .io_args_out_5(pipe1_io_args_out_5),
    .io_args_out_6(pipe1_io_args_out_6),
    .io_vliw_out_0(pipe1_io_vliw_out_0),
    .io_vliw_out_1(pipe1_io_vliw_out_1),
    .io_vliw_out_2(pipe1_io_vliw_out_2),
    .io_vliw_out_3(pipe1_io_vliw_out_3),
    .io_action_mod_en(pipe1_io_action_mod_en),
    .io_action_mod_addr(pipe1_io_action_mod_addr),
    .io_action_mod_data_0(pipe1_io_action_mod_data_0),
    .io_action_mod_data_1(pipe1_io_action_mod_data_1)
  );
  PrimitiveGetOffset pipe2 ( // @[executor.scala 300:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_args_in_0(pipe2_io_args_in_0),
    .io_args_in_1(pipe2_io_args_in_1),
    .io_args_in_2(pipe2_io_args_in_2),
    .io_args_in_3(pipe2_io_args_in_3),
    .io_args_in_4(pipe2_io_args_in_4),
    .io_args_in_5(pipe2_io_args_in_5),
    .io_args_in_6(pipe2_io_args_in_6),
    .io_vliw_in_0(pipe2_io_vliw_in_0),
    .io_vliw_in_1(pipe2_io_vliw_in_1),
    .io_vliw_in_2(pipe2_io_vliw_in_2),
    .io_vliw_in_3(pipe2_io_vliw_in_3),
    .io_args_out_0(pipe2_io_args_out_0),
    .io_args_out_1(pipe2_io_args_out_1),
    .io_args_out_2(pipe2_io_args_out_2),
    .io_args_out_3(pipe2_io_args_out_3),
    .io_args_out_4(pipe2_io_args_out_4),
    .io_args_out_5(pipe2_io_args_out_5),
    .io_args_out_6(pipe2_io_args_out_6),
    .io_vliw_out_0(pipe2_io_vliw_out_0),
    .io_vliw_out_1(pipe2_io_vliw_out_1),
    .io_vliw_out_2(pipe2_io_vliw_out_2),
    .io_vliw_out_3(pipe2_io_vliw_out_3),
    .io_offset_out_0(pipe2_io_offset_out_0),
    .io_offset_out_1(pipe2_io_offset_out_1),
    .io_offset_out_2(pipe2_io_offset_out_2),
    .io_offset_out_3(pipe2_io_offset_out_3),
    .io_length_out_0(pipe2_io_length_out_0),
    .io_length_out_1(pipe2_io_length_out_1),
    .io_length_out_2(pipe2_io_length_out_2),
    .io_length_out_3(pipe2_io_length_out_3)
  );
  PrimitiveGetSource pipe3 ( // @[executor.scala 301:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_args_in_0(pipe3_io_args_in_0),
    .io_args_in_1(pipe3_io_args_in_1),
    .io_args_in_2(pipe3_io_args_in_2),
    .io_args_in_3(pipe3_io_args_in_3),
    .io_args_in_4(pipe3_io_args_in_4),
    .io_args_in_5(pipe3_io_args_in_5),
    .io_args_in_6(pipe3_io_args_in_6),
    .io_vliw_in_0(pipe3_io_vliw_in_0),
    .io_vliw_in_1(pipe3_io_vliw_in_1),
    .io_vliw_in_2(pipe3_io_vliw_in_2),
    .io_vliw_in_3(pipe3_io_vliw_in_3),
    .io_offset_in_0(pipe3_io_offset_in_0),
    .io_offset_in_1(pipe3_io_offset_in_1),
    .io_offset_in_2(pipe3_io_offset_in_2),
    .io_offset_in_3(pipe3_io_offset_in_3),
    .io_length_in_0(pipe3_io_length_in_0),
    .io_length_in_1(pipe3_io_length_in_1),
    .io_length_in_2(pipe3_io_length_in_2),
    .io_length_in_3(pipe3_io_length_in_3),
    .io_vliw_out_0(pipe3_io_vliw_out_0),
    .io_vliw_out_1(pipe3_io_vliw_out_1),
    .io_vliw_out_2(pipe3_io_vliw_out_2),
    .io_vliw_out_3(pipe3_io_vliw_out_3),
    .io_field_out_0(pipe3_io_field_out_0),
    .io_field_out_1(pipe3_io_field_out_1),
    .io_field_out_2(pipe3_io_field_out_2),
    .io_field_out_3(pipe3_io_field_out_3)
  );
  PrimitiveALU pipe4 ( // @[executor.scala 302:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_vliw_in_0(pipe4_io_vliw_in_0),
    .io_vliw_in_1(pipe4_io_vliw_in_1),
    .io_vliw_in_2(pipe4_io_vliw_in_2),
    .io_vliw_in_3(pipe4_io_vliw_in_3),
    .io_field_in_0(pipe4_io_field_in_0),
    .io_field_in_1(pipe4_io_field_in_1),
    .io_field_in_2(pipe4_io_field_in_2),
    .io_field_in_3(pipe4_io_field_in_3),
    .io_vliw_out_0(pipe4_io_vliw_out_0),
    .io_vliw_out_1(pipe4_io_vliw_out_1),
    .io_vliw_out_2(pipe4_io_vliw_out_2),
    .io_vliw_out_3(pipe4_io_vliw_out_3),
    .io_field_out_0(pipe4_io_field_out_0),
    .io_field_out_1(pipe4_io_field_out_1),
    .io_field_out_2(pipe4_io_field_out_2),
    .io_field_out_3(pipe4_io_field_out_3)
  );
  PrimitiveGetWriteBackOffset pipe5 ( // @[executor.scala 303:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_vliw_in_0(pipe5_io_vliw_in_0),
    .io_vliw_in_1(pipe5_io_vliw_in_1),
    .io_vliw_in_2(pipe5_io_vliw_in_2),
    .io_vliw_in_3(pipe5_io_vliw_in_3),
    .io_field_in_0(pipe5_io_field_in_0),
    .io_field_in_1(pipe5_io_field_in_1),
    .io_field_in_2(pipe5_io_field_in_2),
    .io_field_in_3(pipe5_io_field_in_3),
    .io_offset_out_0(pipe5_io_offset_out_0),
    .io_offset_out_1(pipe5_io_offset_out_1),
    .io_offset_out_2(pipe5_io_offset_out_2),
    .io_offset_out_3(pipe5_io_offset_out_3),
    .io_length_out_0(pipe5_io_length_out_0),
    .io_length_out_1(pipe5_io_length_out_1),
    .io_length_out_2(pipe5_io_length_out_2),
    .io_length_out_3(pipe5_io_length_out_3),
    .io_field_out_0(pipe5_io_field_out_0),
    .io_field_out_1(pipe5_io_field_out_1),
    .io_field_out_2(pipe5_io_field_out_2),
    .io_field_out_3(pipe5_io_field_out_3)
  );
  PrimitiveWriteBack pipe6 ( // @[executor.scala 304:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_offset_in_0(pipe6_io_offset_in_0),
    .io_offset_in_1(pipe6_io_offset_in_1),
    .io_offset_in_2(pipe6_io_offset_in_2),
    .io_offset_in_3(pipe6_io_offset_in_3),
    .io_length_in_0(pipe6_io_length_in_0),
    .io_length_in_1(pipe6_io_length_in_1),
    .io_length_in_2(pipe6_io_length_in_2),
    .io_length_in_3(pipe6_io_length_in_3),
    .io_field_in_0(pipe6_io_field_in_0),
    .io_field_in_1(pipe6_io_field_in_1),
    .io_field_in_2(pipe6_io_field_in_2),
    .io_field_in_3(pipe6_io_field_in_3)
  );
  assign io_pipe_phv_out_data_0 = pipe6_io_pipe_phv_out_data_0; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_1 = pipe6_io_pipe_phv_out_data_1; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_2 = pipe6_io_pipe_phv_out_data_2; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_3 = pipe6_io_pipe_phv_out_data_3; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_4 = pipe6_io_pipe_phv_out_data_4; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_5 = pipe6_io_pipe_phv_out_data_5; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_6 = pipe6_io_pipe_phv_out_data_6; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_7 = pipe6_io_pipe_phv_out_data_7; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_8 = pipe6_io_pipe_phv_out_data_8; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_9 = pipe6_io_pipe_phv_out_data_9; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_10 = pipe6_io_pipe_phv_out_data_10; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_11 = pipe6_io_pipe_phv_out_data_11; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_12 = pipe6_io_pipe_phv_out_data_12; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_13 = pipe6_io_pipe_phv_out_data_13; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_14 = pipe6_io_pipe_phv_out_data_14; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_15 = pipe6_io_pipe_phv_out_data_15; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_16 = pipe6_io_pipe_phv_out_data_16; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_17 = pipe6_io_pipe_phv_out_data_17; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_18 = pipe6_io_pipe_phv_out_data_18; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_19 = pipe6_io_pipe_phv_out_data_19; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_20 = pipe6_io_pipe_phv_out_data_20; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_21 = pipe6_io_pipe_phv_out_data_21; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_22 = pipe6_io_pipe_phv_out_data_22; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_23 = pipe6_io_pipe_phv_out_data_23; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_24 = pipe6_io_pipe_phv_out_data_24; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_25 = pipe6_io_pipe_phv_out_data_25; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_26 = pipe6_io_pipe_phv_out_data_26; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_27 = pipe6_io_pipe_phv_out_data_27; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_28 = pipe6_io_pipe_phv_out_data_28; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_29 = pipe6_io_pipe_phv_out_data_29; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_30 = pipe6_io_pipe_phv_out_data_30; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_31 = pipe6_io_pipe_phv_out_data_31; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_32 = pipe6_io_pipe_phv_out_data_32; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_33 = pipe6_io_pipe_phv_out_data_33; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_34 = pipe6_io_pipe_phv_out_data_34; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_35 = pipe6_io_pipe_phv_out_data_35; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_36 = pipe6_io_pipe_phv_out_data_36; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_37 = pipe6_io_pipe_phv_out_data_37; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_38 = pipe6_io_pipe_phv_out_data_38; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_39 = pipe6_io_pipe_phv_out_data_39; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_40 = pipe6_io_pipe_phv_out_data_40; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_41 = pipe6_io_pipe_phv_out_data_41; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_42 = pipe6_io_pipe_phv_out_data_42; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_43 = pipe6_io_pipe_phv_out_data_43; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_44 = pipe6_io_pipe_phv_out_data_44; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_45 = pipe6_io_pipe_phv_out_data_45; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_46 = pipe6_io_pipe_phv_out_data_46; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_47 = pipe6_io_pipe_phv_out_data_47; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_48 = pipe6_io_pipe_phv_out_data_48; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_49 = pipe6_io_pipe_phv_out_data_49; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_50 = pipe6_io_pipe_phv_out_data_50; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_51 = pipe6_io_pipe_phv_out_data_51; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_52 = pipe6_io_pipe_phv_out_data_52; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_53 = pipe6_io_pipe_phv_out_data_53; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_54 = pipe6_io_pipe_phv_out_data_54; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_55 = pipe6_io_pipe_phv_out_data_55; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_56 = pipe6_io_pipe_phv_out_data_56; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_57 = pipe6_io_pipe_phv_out_data_57; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_58 = pipe6_io_pipe_phv_out_data_58; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_59 = pipe6_io_pipe_phv_out_data_59; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_60 = pipe6_io_pipe_phv_out_data_60; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_61 = pipe6_io_pipe_phv_out_data_61; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_62 = pipe6_io_pipe_phv_out_data_62; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_63 = pipe6_io_pipe_phv_out_data_63; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_64 = pipe6_io_pipe_phv_out_data_64; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_65 = pipe6_io_pipe_phv_out_data_65; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_66 = pipe6_io_pipe_phv_out_data_66; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_67 = pipe6_io_pipe_phv_out_data_67; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_68 = pipe6_io_pipe_phv_out_data_68; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_69 = pipe6_io_pipe_phv_out_data_69; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_70 = pipe6_io_pipe_phv_out_data_70; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_71 = pipe6_io_pipe_phv_out_data_71; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_72 = pipe6_io_pipe_phv_out_data_72; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_73 = pipe6_io_pipe_phv_out_data_73; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_74 = pipe6_io_pipe_phv_out_data_74; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_75 = pipe6_io_pipe_phv_out_data_75; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_76 = pipe6_io_pipe_phv_out_data_76; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_77 = pipe6_io_pipe_phv_out_data_77; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_78 = pipe6_io_pipe_phv_out_data_78; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_79 = pipe6_io_pipe_phv_out_data_79; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_80 = pipe6_io_pipe_phv_out_data_80; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_81 = pipe6_io_pipe_phv_out_data_81; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_82 = pipe6_io_pipe_phv_out_data_82; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_83 = pipe6_io_pipe_phv_out_data_83; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_84 = pipe6_io_pipe_phv_out_data_84; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_85 = pipe6_io_pipe_phv_out_data_85; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_86 = pipe6_io_pipe_phv_out_data_86; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_87 = pipe6_io_pipe_phv_out_data_87; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_88 = pipe6_io_pipe_phv_out_data_88; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_89 = pipe6_io_pipe_phv_out_data_89; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_90 = pipe6_io_pipe_phv_out_data_90; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_91 = pipe6_io_pipe_phv_out_data_91; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_92 = pipe6_io_pipe_phv_out_data_92; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_93 = pipe6_io_pipe_phv_out_data_93; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_94 = pipe6_io_pipe_phv_out_data_94; // @[executor.scala 334:27]
  assign io_pipe_phv_out_data_95 = pipe6_io_pipe_phv_out_data_95; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_0 = pipe6_io_pipe_phv_out_header_0; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_1 = pipe6_io_pipe_phv_out_header_1; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_2 = pipe6_io_pipe_phv_out_header_2; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_3 = pipe6_io_pipe_phv_out_header_3; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_4 = pipe6_io_pipe_phv_out_header_4; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_5 = pipe6_io_pipe_phv_out_header_5; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_6 = pipe6_io_pipe_phv_out_header_6; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_7 = pipe6_io_pipe_phv_out_header_7; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_8 = pipe6_io_pipe_phv_out_header_8; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_9 = pipe6_io_pipe_phv_out_header_9; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_10 = pipe6_io_pipe_phv_out_header_10; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_11 = pipe6_io_pipe_phv_out_header_11; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_12 = pipe6_io_pipe_phv_out_header_12; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_13 = pipe6_io_pipe_phv_out_header_13; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_14 = pipe6_io_pipe_phv_out_header_14; // @[executor.scala 334:27]
  assign io_pipe_phv_out_header_15 = pipe6_io_pipe_phv_out_header_15; // @[executor.scala 334:27]
  assign io_pipe_phv_out_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 334:27]
  assign io_pipe_phv_out_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 334:27]
  assign io_pipe_phv_out_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 334:27]
  assign io_pipe_phv_out_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 334:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[executor.scala 306:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[executor.scala 306:26]
  assign pipe1_io_hit = io_hit; // @[executor.scala 307:26]
  assign pipe1_io_match_value = io_match_value; // @[executor.scala 308:26]
  assign pipe1_io_action_mod_en = io_action_mod_en; // @[executor.scala 309:26]
  assign pipe1_io_action_mod_addr = io_action_mod_addr; // @[executor.scala 309:26]
  assign pipe1_io_action_mod_data_0 = io_action_mod_data_0; // @[executor.scala 309:26]
  assign pipe1_io_action_mod_data_1 = io_action_mod_data_1; // @[executor.scala 309:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 311:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 311:26]
  assign pipe2_io_args_in_0 = pipe1_io_args_out_0; // @[executor.scala 312:26]
  assign pipe2_io_args_in_1 = pipe1_io_args_out_1; // @[executor.scala 312:26]
  assign pipe2_io_args_in_2 = pipe1_io_args_out_2; // @[executor.scala 312:26]
  assign pipe2_io_args_in_3 = pipe1_io_args_out_3; // @[executor.scala 312:26]
  assign pipe2_io_args_in_4 = pipe1_io_args_out_4; // @[executor.scala 312:26]
  assign pipe2_io_args_in_5 = pipe1_io_args_out_5; // @[executor.scala 312:26]
  assign pipe2_io_args_in_6 = pipe1_io_args_out_6; // @[executor.scala 312:26]
  assign pipe2_io_vliw_in_0 = pipe1_io_vliw_out_0; // @[executor.scala 313:26]
  assign pipe2_io_vliw_in_1 = pipe1_io_vliw_out_1; // @[executor.scala 313:26]
  assign pipe2_io_vliw_in_2 = pipe1_io_vliw_out_2; // @[executor.scala 313:26]
  assign pipe2_io_vliw_in_3 = pipe1_io_vliw_out_3; // @[executor.scala 313:26]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 315:26]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 315:26]
  assign pipe3_io_args_in_0 = pipe2_io_args_out_0; // @[executor.scala 316:26]
  assign pipe3_io_args_in_1 = pipe2_io_args_out_1; // @[executor.scala 316:26]
  assign pipe3_io_args_in_2 = pipe2_io_args_out_2; // @[executor.scala 316:26]
  assign pipe3_io_args_in_3 = pipe2_io_args_out_3; // @[executor.scala 316:26]
  assign pipe3_io_args_in_4 = pipe2_io_args_out_4; // @[executor.scala 316:26]
  assign pipe3_io_args_in_5 = pipe2_io_args_out_5; // @[executor.scala 316:26]
  assign pipe3_io_args_in_6 = pipe2_io_args_out_6; // @[executor.scala 316:26]
  assign pipe3_io_vliw_in_0 = pipe2_io_vliw_out_0; // @[executor.scala 317:26]
  assign pipe3_io_vliw_in_1 = pipe2_io_vliw_out_1; // @[executor.scala 317:26]
  assign pipe3_io_vliw_in_2 = pipe2_io_vliw_out_2; // @[executor.scala 317:26]
  assign pipe3_io_vliw_in_3 = pipe2_io_vliw_out_3; // @[executor.scala 317:26]
  assign pipe3_io_offset_in_0 = pipe2_io_offset_out_0; // @[executor.scala 318:26]
  assign pipe3_io_offset_in_1 = pipe2_io_offset_out_1; // @[executor.scala 318:26]
  assign pipe3_io_offset_in_2 = pipe2_io_offset_out_2; // @[executor.scala 318:26]
  assign pipe3_io_offset_in_3 = pipe2_io_offset_out_3; // @[executor.scala 318:26]
  assign pipe3_io_length_in_0 = pipe2_io_length_out_0; // @[executor.scala 319:26]
  assign pipe3_io_length_in_1 = pipe2_io_length_out_1; // @[executor.scala 319:26]
  assign pipe3_io_length_in_2 = pipe2_io_length_out_2; // @[executor.scala 319:26]
  assign pipe3_io_length_in_3 = pipe2_io_length_out_3; // @[executor.scala 319:26]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 321:26]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 321:26]
  assign pipe4_io_vliw_in_0 = pipe3_io_vliw_out_0; // @[executor.scala 322:26]
  assign pipe4_io_vliw_in_1 = pipe3_io_vliw_out_1; // @[executor.scala 322:26]
  assign pipe4_io_vliw_in_2 = pipe3_io_vliw_out_2; // @[executor.scala 322:26]
  assign pipe4_io_vliw_in_3 = pipe3_io_vliw_out_3; // @[executor.scala 322:26]
  assign pipe4_io_field_in_0 = pipe3_io_field_out_0; // @[executor.scala 323:26]
  assign pipe4_io_field_in_1 = pipe3_io_field_out_1; // @[executor.scala 323:26]
  assign pipe4_io_field_in_2 = pipe3_io_field_out_2; // @[executor.scala 323:26]
  assign pipe4_io_field_in_3 = pipe3_io_field_out_3; // @[executor.scala 323:26]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 325:26]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 325:26]
  assign pipe5_io_vliw_in_0 = pipe4_io_vliw_out_0; // @[executor.scala 326:26]
  assign pipe5_io_vliw_in_1 = pipe4_io_vliw_out_1; // @[executor.scala 326:26]
  assign pipe5_io_vliw_in_2 = pipe4_io_vliw_out_2; // @[executor.scala 326:26]
  assign pipe5_io_vliw_in_3 = pipe4_io_vliw_out_3; // @[executor.scala 326:26]
  assign pipe5_io_field_in_0 = pipe4_io_field_out_0; // @[executor.scala 327:26]
  assign pipe5_io_field_in_1 = pipe4_io_field_out_1; // @[executor.scala 327:26]
  assign pipe5_io_field_in_2 = pipe4_io_field_out_2; // @[executor.scala 327:26]
  assign pipe5_io_field_in_3 = pipe4_io_field_out_3; // @[executor.scala 327:26]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 329:26]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 329:26]
  assign pipe6_io_offset_in_0 = pipe5_io_offset_out_0; // @[executor.scala 331:26]
  assign pipe6_io_offset_in_1 = pipe5_io_offset_out_1; // @[executor.scala 331:26]
  assign pipe6_io_offset_in_2 = pipe5_io_offset_out_2; // @[executor.scala 331:26]
  assign pipe6_io_offset_in_3 = pipe5_io_offset_out_3; // @[executor.scala 331:26]
  assign pipe6_io_length_in_0 = pipe5_io_length_out_0; // @[executor.scala 332:26]
  assign pipe6_io_length_in_1 = pipe5_io_length_out_1; // @[executor.scala 332:26]
  assign pipe6_io_length_in_2 = pipe5_io_length_out_2; // @[executor.scala 332:26]
  assign pipe6_io_length_in_3 = pipe5_io_length_out_3; // @[executor.scala 332:26]
  assign pipe6_io_field_in_0 = pipe5_io_field_out_0; // @[executor.scala 330:26]
  assign pipe6_io_field_in_1 = pipe5_io_field_out_1; // @[executor.scala 330:26]
  assign pipe6_io_field_in_2 = pipe5_io_field_out_2; // @[executor.scala 330:26]
  assign pipe6_io_field_in_3 = pipe5_io_field_out_3; // @[executor.scala 330:26]
endmodule
