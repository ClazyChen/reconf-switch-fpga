module PrimitiveWriteBack(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [31:0] io_field_in_0,
  input  [31:0] io_field_in_1,
  input  [31:0] io_field_in_2,
  input  [31:0] io_field_in_3,
  input  [3:0]  io_mask_in_0,
  input  [3:0]  io_mask_in_1,
  input  [3:0]  io_mask_in_2,
  input  [3:0]  io_mask_in_3,
  input  [5:0]  io_dst_offset_in_0,
  input  [5:0]  io_dst_offset_in_1,
  input  [5:0]  io_dst_offset_in_2,
  input  [5:0]  io_dst_offset_in_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 448:22]
  reg [7:0] phv_data_1; // @[executor.scala 448:22]
  reg [7:0] phv_data_2; // @[executor.scala 448:22]
  reg [7:0] phv_data_3; // @[executor.scala 448:22]
  reg [7:0] phv_data_4; // @[executor.scala 448:22]
  reg [7:0] phv_data_5; // @[executor.scala 448:22]
  reg [7:0] phv_data_6; // @[executor.scala 448:22]
  reg [7:0] phv_data_7; // @[executor.scala 448:22]
  reg [7:0] phv_data_8; // @[executor.scala 448:22]
  reg [7:0] phv_data_9; // @[executor.scala 448:22]
  reg [7:0] phv_data_10; // @[executor.scala 448:22]
  reg [7:0] phv_data_11; // @[executor.scala 448:22]
  reg [7:0] phv_data_12; // @[executor.scala 448:22]
  reg [7:0] phv_data_13; // @[executor.scala 448:22]
  reg [7:0] phv_data_14; // @[executor.scala 448:22]
  reg [7:0] phv_data_15; // @[executor.scala 448:22]
  reg [7:0] phv_data_16; // @[executor.scala 448:22]
  reg [7:0] phv_data_17; // @[executor.scala 448:22]
  reg [7:0] phv_data_18; // @[executor.scala 448:22]
  reg [7:0] phv_data_19; // @[executor.scala 448:22]
  reg [7:0] phv_data_20; // @[executor.scala 448:22]
  reg [7:0] phv_data_21; // @[executor.scala 448:22]
  reg [7:0] phv_data_22; // @[executor.scala 448:22]
  reg [7:0] phv_data_23; // @[executor.scala 448:22]
  reg [7:0] phv_data_24; // @[executor.scala 448:22]
  reg [7:0] phv_data_25; // @[executor.scala 448:22]
  reg [7:0] phv_data_26; // @[executor.scala 448:22]
  reg [7:0] phv_data_27; // @[executor.scala 448:22]
  reg [7:0] phv_data_28; // @[executor.scala 448:22]
  reg [7:0] phv_data_29; // @[executor.scala 448:22]
  reg [7:0] phv_data_30; // @[executor.scala 448:22]
  reg [7:0] phv_data_31; // @[executor.scala 448:22]
  reg [7:0] phv_data_32; // @[executor.scala 448:22]
  reg [7:0] phv_data_33; // @[executor.scala 448:22]
  reg [7:0] phv_data_34; // @[executor.scala 448:22]
  reg [7:0] phv_data_35; // @[executor.scala 448:22]
  reg [7:0] phv_data_36; // @[executor.scala 448:22]
  reg [7:0] phv_data_37; // @[executor.scala 448:22]
  reg [7:0] phv_data_38; // @[executor.scala 448:22]
  reg [7:0] phv_data_39; // @[executor.scala 448:22]
  reg [7:0] phv_data_40; // @[executor.scala 448:22]
  reg [7:0] phv_data_41; // @[executor.scala 448:22]
  reg [7:0] phv_data_42; // @[executor.scala 448:22]
  reg [7:0] phv_data_43; // @[executor.scala 448:22]
  reg [7:0] phv_data_44; // @[executor.scala 448:22]
  reg [7:0] phv_data_45; // @[executor.scala 448:22]
  reg [7:0] phv_data_46; // @[executor.scala 448:22]
  reg [7:0] phv_data_47; // @[executor.scala 448:22]
  reg [7:0] phv_data_48; // @[executor.scala 448:22]
  reg [7:0] phv_data_49; // @[executor.scala 448:22]
  reg [7:0] phv_data_50; // @[executor.scala 448:22]
  reg [7:0] phv_data_51; // @[executor.scala 448:22]
  reg [7:0] phv_data_52; // @[executor.scala 448:22]
  reg [7:0] phv_data_53; // @[executor.scala 448:22]
  reg [7:0] phv_data_54; // @[executor.scala 448:22]
  reg [7:0] phv_data_55; // @[executor.scala 448:22]
  reg [7:0] phv_data_56; // @[executor.scala 448:22]
  reg [7:0] phv_data_57; // @[executor.scala 448:22]
  reg [7:0] phv_data_58; // @[executor.scala 448:22]
  reg [7:0] phv_data_59; // @[executor.scala 448:22]
  reg [7:0] phv_data_60; // @[executor.scala 448:22]
  reg [7:0] phv_data_61; // @[executor.scala 448:22]
  reg [7:0] phv_data_62; // @[executor.scala 448:22]
  reg [7:0] phv_data_63; // @[executor.scala 448:22]
  reg [7:0] phv_data_64; // @[executor.scala 448:22]
  reg [7:0] phv_data_65; // @[executor.scala 448:22]
  reg [7:0] phv_data_66; // @[executor.scala 448:22]
  reg [7:0] phv_data_67; // @[executor.scala 448:22]
  reg [7:0] phv_data_68; // @[executor.scala 448:22]
  reg [7:0] phv_data_69; // @[executor.scala 448:22]
  reg [7:0] phv_data_70; // @[executor.scala 448:22]
  reg [7:0] phv_data_71; // @[executor.scala 448:22]
  reg [7:0] phv_data_72; // @[executor.scala 448:22]
  reg [7:0] phv_data_73; // @[executor.scala 448:22]
  reg [7:0] phv_data_74; // @[executor.scala 448:22]
  reg [7:0] phv_data_75; // @[executor.scala 448:22]
  reg [7:0] phv_data_76; // @[executor.scala 448:22]
  reg [7:0] phv_data_77; // @[executor.scala 448:22]
  reg [7:0] phv_data_78; // @[executor.scala 448:22]
  reg [7:0] phv_data_79; // @[executor.scala 448:22]
  reg [7:0] phv_data_80; // @[executor.scala 448:22]
  reg [7:0] phv_data_81; // @[executor.scala 448:22]
  reg [7:0] phv_data_82; // @[executor.scala 448:22]
  reg [7:0] phv_data_83; // @[executor.scala 448:22]
  reg [7:0] phv_data_84; // @[executor.scala 448:22]
  reg [7:0] phv_data_85; // @[executor.scala 448:22]
  reg [7:0] phv_data_86; // @[executor.scala 448:22]
  reg [7:0] phv_data_87; // @[executor.scala 448:22]
  reg [7:0] phv_data_88; // @[executor.scala 448:22]
  reg [7:0] phv_data_89; // @[executor.scala 448:22]
  reg [7:0] phv_data_90; // @[executor.scala 448:22]
  reg [7:0] phv_data_91; // @[executor.scala 448:22]
  reg [7:0] phv_data_92; // @[executor.scala 448:22]
  reg [7:0] phv_data_93; // @[executor.scala 448:22]
  reg [7:0] phv_data_94; // @[executor.scala 448:22]
  reg [7:0] phv_data_95; // @[executor.scala 448:22]
  reg [7:0] phv_data_96; // @[executor.scala 448:22]
  reg [7:0] phv_data_97; // @[executor.scala 448:22]
  reg [7:0] phv_data_98; // @[executor.scala 448:22]
  reg [7:0] phv_data_99; // @[executor.scala 448:22]
  reg [7:0] phv_data_100; // @[executor.scala 448:22]
  reg [7:0] phv_data_101; // @[executor.scala 448:22]
  reg [7:0] phv_data_102; // @[executor.scala 448:22]
  reg [7:0] phv_data_103; // @[executor.scala 448:22]
  reg [7:0] phv_data_104; // @[executor.scala 448:22]
  reg [7:0] phv_data_105; // @[executor.scala 448:22]
  reg [7:0] phv_data_106; // @[executor.scala 448:22]
  reg [7:0] phv_data_107; // @[executor.scala 448:22]
  reg [7:0] phv_data_108; // @[executor.scala 448:22]
  reg [7:0] phv_data_109; // @[executor.scala 448:22]
  reg [7:0] phv_data_110; // @[executor.scala 448:22]
  reg [7:0] phv_data_111; // @[executor.scala 448:22]
  reg [7:0] phv_data_112; // @[executor.scala 448:22]
  reg [7:0] phv_data_113; // @[executor.scala 448:22]
  reg [7:0] phv_data_114; // @[executor.scala 448:22]
  reg [7:0] phv_data_115; // @[executor.scala 448:22]
  reg [7:0] phv_data_116; // @[executor.scala 448:22]
  reg [7:0] phv_data_117; // @[executor.scala 448:22]
  reg [7:0] phv_data_118; // @[executor.scala 448:22]
  reg [7:0] phv_data_119; // @[executor.scala 448:22]
  reg [7:0] phv_data_120; // @[executor.scala 448:22]
  reg [7:0] phv_data_121; // @[executor.scala 448:22]
  reg [7:0] phv_data_122; // @[executor.scala 448:22]
  reg [7:0] phv_data_123; // @[executor.scala 448:22]
  reg [7:0] phv_data_124; // @[executor.scala 448:22]
  reg [7:0] phv_data_125; // @[executor.scala 448:22]
  reg [7:0] phv_data_126; // @[executor.scala 448:22]
  reg [7:0] phv_data_127; // @[executor.scala 448:22]
  reg [7:0] phv_data_128; // @[executor.scala 448:22]
  reg [7:0] phv_data_129; // @[executor.scala 448:22]
  reg [7:0] phv_data_130; // @[executor.scala 448:22]
  reg [7:0] phv_data_131; // @[executor.scala 448:22]
  reg [7:0] phv_data_132; // @[executor.scala 448:22]
  reg [7:0] phv_data_133; // @[executor.scala 448:22]
  reg [7:0] phv_data_134; // @[executor.scala 448:22]
  reg [7:0] phv_data_135; // @[executor.scala 448:22]
  reg [7:0] phv_data_136; // @[executor.scala 448:22]
  reg [7:0] phv_data_137; // @[executor.scala 448:22]
  reg [7:0] phv_data_138; // @[executor.scala 448:22]
  reg [7:0] phv_data_139; // @[executor.scala 448:22]
  reg [7:0] phv_data_140; // @[executor.scala 448:22]
  reg [7:0] phv_data_141; // @[executor.scala 448:22]
  reg [7:0] phv_data_142; // @[executor.scala 448:22]
  reg [7:0] phv_data_143; // @[executor.scala 448:22]
  reg [7:0] phv_data_144; // @[executor.scala 448:22]
  reg [7:0] phv_data_145; // @[executor.scala 448:22]
  reg [7:0] phv_data_146; // @[executor.scala 448:22]
  reg [7:0] phv_data_147; // @[executor.scala 448:22]
  reg [7:0] phv_data_148; // @[executor.scala 448:22]
  reg [7:0] phv_data_149; // @[executor.scala 448:22]
  reg [7:0] phv_data_150; // @[executor.scala 448:22]
  reg [7:0] phv_data_151; // @[executor.scala 448:22]
  reg [7:0] phv_data_152; // @[executor.scala 448:22]
  reg [7:0] phv_data_153; // @[executor.scala 448:22]
  reg [7:0] phv_data_154; // @[executor.scala 448:22]
  reg [7:0] phv_data_155; // @[executor.scala 448:22]
  reg [7:0] phv_data_156; // @[executor.scala 448:22]
  reg [7:0] phv_data_157; // @[executor.scala 448:22]
  reg [7:0] phv_data_158; // @[executor.scala 448:22]
  reg [7:0] phv_data_159; // @[executor.scala 448:22]
  reg [7:0] phv_data_160; // @[executor.scala 448:22]
  reg [7:0] phv_data_161; // @[executor.scala 448:22]
  reg [7:0] phv_data_162; // @[executor.scala 448:22]
  reg [7:0] phv_data_163; // @[executor.scala 448:22]
  reg [7:0] phv_data_164; // @[executor.scala 448:22]
  reg [7:0] phv_data_165; // @[executor.scala 448:22]
  reg [7:0] phv_data_166; // @[executor.scala 448:22]
  reg [7:0] phv_data_167; // @[executor.scala 448:22]
  reg [7:0] phv_data_168; // @[executor.scala 448:22]
  reg [7:0] phv_data_169; // @[executor.scala 448:22]
  reg [7:0] phv_data_170; // @[executor.scala 448:22]
  reg [7:0] phv_data_171; // @[executor.scala 448:22]
  reg [7:0] phv_data_172; // @[executor.scala 448:22]
  reg [7:0] phv_data_173; // @[executor.scala 448:22]
  reg [7:0] phv_data_174; // @[executor.scala 448:22]
  reg [7:0] phv_data_175; // @[executor.scala 448:22]
  reg [7:0] phv_data_176; // @[executor.scala 448:22]
  reg [7:0] phv_data_177; // @[executor.scala 448:22]
  reg [7:0] phv_data_178; // @[executor.scala 448:22]
  reg [7:0] phv_data_179; // @[executor.scala 448:22]
  reg [7:0] phv_data_180; // @[executor.scala 448:22]
  reg [7:0] phv_data_181; // @[executor.scala 448:22]
  reg [7:0] phv_data_182; // @[executor.scala 448:22]
  reg [7:0] phv_data_183; // @[executor.scala 448:22]
  reg [7:0] phv_data_184; // @[executor.scala 448:22]
  reg [7:0] phv_data_185; // @[executor.scala 448:22]
  reg [7:0] phv_data_186; // @[executor.scala 448:22]
  reg [7:0] phv_data_187; // @[executor.scala 448:22]
  reg [7:0] phv_data_188; // @[executor.scala 448:22]
  reg [7:0] phv_data_189; // @[executor.scala 448:22]
  reg [7:0] phv_data_190; // @[executor.scala 448:22]
  reg [7:0] phv_data_191; // @[executor.scala 448:22]
  reg [7:0] phv_data_192; // @[executor.scala 448:22]
  reg [7:0] phv_data_193; // @[executor.scala 448:22]
  reg [7:0] phv_data_194; // @[executor.scala 448:22]
  reg [7:0] phv_data_195; // @[executor.scala 448:22]
  reg [7:0] phv_data_196; // @[executor.scala 448:22]
  reg [7:0] phv_data_197; // @[executor.scala 448:22]
  reg [7:0] phv_data_198; // @[executor.scala 448:22]
  reg [7:0] phv_data_199; // @[executor.scala 448:22]
  reg [7:0] phv_data_200; // @[executor.scala 448:22]
  reg [7:0] phv_data_201; // @[executor.scala 448:22]
  reg [7:0] phv_data_202; // @[executor.scala 448:22]
  reg [7:0] phv_data_203; // @[executor.scala 448:22]
  reg [7:0] phv_data_204; // @[executor.scala 448:22]
  reg [7:0] phv_data_205; // @[executor.scala 448:22]
  reg [7:0] phv_data_206; // @[executor.scala 448:22]
  reg [7:0] phv_data_207; // @[executor.scala 448:22]
  reg [7:0] phv_data_208; // @[executor.scala 448:22]
  reg [7:0] phv_data_209; // @[executor.scala 448:22]
  reg [7:0] phv_data_210; // @[executor.scala 448:22]
  reg [7:0] phv_data_211; // @[executor.scala 448:22]
  reg [7:0] phv_data_212; // @[executor.scala 448:22]
  reg [7:0] phv_data_213; // @[executor.scala 448:22]
  reg [7:0] phv_data_214; // @[executor.scala 448:22]
  reg [7:0] phv_data_215; // @[executor.scala 448:22]
  reg [7:0] phv_data_216; // @[executor.scala 448:22]
  reg [7:0] phv_data_217; // @[executor.scala 448:22]
  reg [7:0] phv_data_218; // @[executor.scala 448:22]
  reg [7:0] phv_data_219; // @[executor.scala 448:22]
  reg [7:0] phv_data_220; // @[executor.scala 448:22]
  reg [7:0] phv_data_221; // @[executor.scala 448:22]
  reg [7:0] phv_data_222; // @[executor.scala 448:22]
  reg [7:0] phv_data_223; // @[executor.scala 448:22]
  reg [7:0] phv_data_224; // @[executor.scala 448:22]
  reg [7:0] phv_data_225; // @[executor.scala 448:22]
  reg [7:0] phv_data_226; // @[executor.scala 448:22]
  reg [7:0] phv_data_227; // @[executor.scala 448:22]
  reg [7:0] phv_data_228; // @[executor.scala 448:22]
  reg [7:0] phv_data_229; // @[executor.scala 448:22]
  reg [7:0] phv_data_230; // @[executor.scala 448:22]
  reg [7:0] phv_data_231; // @[executor.scala 448:22]
  reg [7:0] phv_data_232; // @[executor.scala 448:22]
  reg [7:0] phv_data_233; // @[executor.scala 448:22]
  reg [7:0] phv_data_234; // @[executor.scala 448:22]
  reg [7:0] phv_data_235; // @[executor.scala 448:22]
  reg [7:0] phv_data_236; // @[executor.scala 448:22]
  reg [7:0] phv_data_237; // @[executor.scala 448:22]
  reg [7:0] phv_data_238; // @[executor.scala 448:22]
  reg [7:0] phv_data_239; // @[executor.scala 448:22]
  reg [7:0] phv_data_240; // @[executor.scala 448:22]
  reg [7:0] phv_data_241; // @[executor.scala 448:22]
  reg [7:0] phv_data_242; // @[executor.scala 448:22]
  reg [7:0] phv_data_243; // @[executor.scala 448:22]
  reg [7:0] phv_data_244; // @[executor.scala 448:22]
  reg [7:0] phv_data_245; // @[executor.scala 448:22]
  reg [7:0] phv_data_246; // @[executor.scala 448:22]
  reg [7:0] phv_data_247; // @[executor.scala 448:22]
  reg [7:0] phv_data_248; // @[executor.scala 448:22]
  reg [7:0] phv_data_249; // @[executor.scala 448:22]
  reg [7:0] phv_data_250; // @[executor.scala 448:22]
  reg [7:0] phv_data_251; // @[executor.scala 448:22]
  reg [7:0] phv_data_252; // @[executor.scala 448:22]
  reg [7:0] phv_data_253; // @[executor.scala 448:22]
  reg [7:0] phv_data_254; // @[executor.scala 448:22]
  reg [7:0] phv_data_255; // @[executor.scala 448:22]
  reg [7:0] phv_data_256; // @[executor.scala 448:22]
  reg [7:0] phv_data_257; // @[executor.scala 448:22]
  reg [7:0] phv_data_258; // @[executor.scala 448:22]
  reg [7:0] phv_data_259; // @[executor.scala 448:22]
  reg [7:0] phv_data_260; // @[executor.scala 448:22]
  reg [7:0] phv_data_261; // @[executor.scala 448:22]
  reg [7:0] phv_data_262; // @[executor.scala 448:22]
  reg [7:0] phv_data_263; // @[executor.scala 448:22]
  reg [7:0] phv_data_264; // @[executor.scala 448:22]
  reg [7:0] phv_data_265; // @[executor.scala 448:22]
  reg [7:0] phv_data_266; // @[executor.scala 448:22]
  reg [7:0] phv_data_267; // @[executor.scala 448:22]
  reg [7:0] phv_data_268; // @[executor.scala 448:22]
  reg [7:0] phv_data_269; // @[executor.scala 448:22]
  reg [7:0] phv_data_270; // @[executor.scala 448:22]
  reg [7:0] phv_data_271; // @[executor.scala 448:22]
  reg [7:0] phv_data_272; // @[executor.scala 448:22]
  reg [7:0] phv_data_273; // @[executor.scala 448:22]
  reg [7:0] phv_data_274; // @[executor.scala 448:22]
  reg [7:0] phv_data_275; // @[executor.scala 448:22]
  reg [7:0] phv_data_276; // @[executor.scala 448:22]
  reg [7:0] phv_data_277; // @[executor.scala 448:22]
  reg [7:0] phv_data_278; // @[executor.scala 448:22]
  reg [7:0] phv_data_279; // @[executor.scala 448:22]
  reg [7:0] phv_data_280; // @[executor.scala 448:22]
  reg [7:0] phv_data_281; // @[executor.scala 448:22]
  reg [7:0] phv_data_282; // @[executor.scala 448:22]
  reg [7:0] phv_data_283; // @[executor.scala 448:22]
  reg [7:0] phv_data_284; // @[executor.scala 448:22]
  reg [7:0] phv_data_285; // @[executor.scala 448:22]
  reg [7:0] phv_data_286; // @[executor.scala 448:22]
  reg [7:0] phv_data_287; // @[executor.scala 448:22]
  reg [7:0] phv_data_288; // @[executor.scala 448:22]
  reg [7:0] phv_data_289; // @[executor.scala 448:22]
  reg [7:0] phv_data_290; // @[executor.scala 448:22]
  reg [7:0] phv_data_291; // @[executor.scala 448:22]
  reg [7:0] phv_data_292; // @[executor.scala 448:22]
  reg [7:0] phv_data_293; // @[executor.scala 448:22]
  reg [7:0] phv_data_294; // @[executor.scala 448:22]
  reg [7:0] phv_data_295; // @[executor.scala 448:22]
  reg [7:0] phv_data_296; // @[executor.scala 448:22]
  reg [7:0] phv_data_297; // @[executor.scala 448:22]
  reg [7:0] phv_data_298; // @[executor.scala 448:22]
  reg [7:0] phv_data_299; // @[executor.scala 448:22]
  reg [7:0] phv_data_300; // @[executor.scala 448:22]
  reg [7:0] phv_data_301; // @[executor.scala 448:22]
  reg [7:0] phv_data_302; // @[executor.scala 448:22]
  reg [7:0] phv_data_303; // @[executor.scala 448:22]
  reg [7:0] phv_data_304; // @[executor.scala 448:22]
  reg [7:0] phv_data_305; // @[executor.scala 448:22]
  reg [7:0] phv_data_306; // @[executor.scala 448:22]
  reg [7:0] phv_data_307; // @[executor.scala 448:22]
  reg [7:0] phv_data_308; // @[executor.scala 448:22]
  reg [7:0] phv_data_309; // @[executor.scala 448:22]
  reg [7:0] phv_data_310; // @[executor.scala 448:22]
  reg [7:0] phv_data_311; // @[executor.scala 448:22]
  reg [7:0] phv_data_312; // @[executor.scala 448:22]
  reg [7:0] phv_data_313; // @[executor.scala 448:22]
  reg [7:0] phv_data_314; // @[executor.scala 448:22]
  reg [7:0] phv_data_315; // @[executor.scala 448:22]
  reg [7:0] phv_data_316; // @[executor.scala 448:22]
  reg [7:0] phv_data_317; // @[executor.scala 448:22]
  reg [7:0] phv_data_318; // @[executor.scala 448:22]
  reg [7:0] phv_data_319; // @[executor.scala 448:22]
  reg [7:0] phv_data_320; // @[executor.scala 448:22]
  reg [7:0] phv_data_321; // @[executor.scala 448:22]
  reg [7:0] phv_data_322; // @[executor.scala 448:22]
  reg [7:0] phv_data_323; // @[executor.scala 448:22]
  reg [7:0] phv_data_324; // @[executor.scala 448:22]
  reg [7:0] phv_data_325; // @[executor.scala 448:22]
  reg [7:0] phv_data_326; // @[executor.scala 448:22]
  reg [7:0] phv_data_327; // @[executor.scala 448:22]
  reg [7:0] phv_data_328; // @[executor.scala 448:22]
  reg [7:0] phv_data_329; // @[executor.scala 448:22]
  reg [7:0] phv_data_330; // @[executor.scala 448:22]
  reg [7:0] phv_data_331; // @[executor.scala 448:22]
  reg [7:0] phv_data_332; // @[executor.scala 448:22]
  reg [7:0] phv_data_333; // @[executor.scala 448:22]
  reg [7:0] phv_data_334; // @[executor.scala 448:22]
  reg [7:0] phv_data_335; // @[executor.scala 448:22]
  reg [7:0] phv_data_336; // @[executor.scala 448:22]
  reg [7:0] phv_data_337; // @[executor.scala 448:22]
  reg [7:0] phv_data_338; // @[executor.scala 448:22]
  reg [7:0] phv_data_339; // @[executor.scala 448:22]
  reg [7:0] phv_data_340; // @[executor.scala 448:22]
  reg [7:0] phv_data_341; // @[executor.scala 448:22]
  reg [7:0] phv_data_342; // @[executor.scala 448:22]
  reg [7:0] phv_data_343; // @[executor.scala 448:22]
  reg [7:0] phv_data_344; // @[executor.scala 448:22]
  reg [7:0] phv_data_345; // @[executor.scala 448:22]
  reg [7:0] phv_data_346; // @[executor.scala 448:22]
  reg [7:0] phv_data_347; // @[executor.scala 448:22]
  reg [7:0] phv_data_348; // @[executor.scala 448:22]
  reg [7:0] phv_data_349; // @[executor.scala 448:22]
  reg [7:0] phv_data_350; // @[executor.scala 448:22]
  reg [7:0] phv_data_351; // @[executor.scala 448:22]
  reg [7:0] phv_data_352; // @[executor.scala 448:22]
  reg [7:0] phv_data_353; // @[executor.scala 448:22]
  reg [7:0] phv_data_354; // @[executor.scala 448:22]
  reg [7:0] phv_data_355; // @[executor.scala 448:22]
  reg [7:0] phv_data_356; // @[executor.scala 448:22]
  reg [7:0] phv_data_357; // @[executor.scala 448:22]
  reg [7:0] phv_data_358; // @[executor.scala 448:22]
  reg [7:0] phv_data_359; // @[executor.scala 448:22]
  reg [7:0] phv_data_360; // @[executor.scala 448:22]
  reg [7:0] phv_data_361; // @[executor.scala 448:22]
  reg [7:0] phv_data_362; // @[executor.scala 448:22]
  reg [7:0] phv_data_363; // @[executor.scala 448:22]
  reg [7:0] phv_data_364; // @[executor.scala 448:22]
  reg [7:0] phv_data_365; // @[executor.scala 448:22]
  reg [7:0] phv_data_366; // @[executor.scala 448:22]
  reg [7:0] phv_data_367; // @[executor.scala 448:22]
  reg [7:0] phv_data_368; // @[executor.scala 448:22]
  reg [7:0] phv_data_369; // @[executor.scala 448:22]
  reg [7:0] phv_data_370; // @[executor.scala 448:22]
  reg [7:0] phv_data_371; // @[executor.scala 448:22]
  reg [7:0] phv_data_372; // @[executor.scala 448:22]
  reg [7:0] phv_data_373; // @[executor.scala 448:22]
  reg [7:0] phv_data_374; // @[executor.scala 448:22]
  reg [7:0] phv_data_375; // @[executor.scala 448:22]
  reg [7:0] phv_data_376; // @[executor.scala 448:22]
  reg [7:0] phv_data_377; // @[executor.scala 448:22]
  reg [7:0] phv_data_378; // @[executor.scala 448:22]
  reg [7:0] phv_data_379; // @[executor.scala 448:22]
  reg [7:0] phv_data_380; // @[executor.scala 448:22]
  reg [7:0] phv_data_381; // @[executor.scala 448:22]
  reg [7:0] phv_data_382; // @[executor.scala 448:22]
  reg [7:0] phv_data_383; // @[executor.scala 448:22]
  reg [7:0] phv_data_384; // @[executor.scala 448:22]
  reg [7:0] phv_data_385; // @[executor.scala 448:22]
  reg [7:0] phv_data_386; // @[executor.scala 448:22]
  reg [7:0] phv_data_387; // @[executor.scala 448:22]
  reg [7:0] phv_data_388; // @[executor.scala 448:22]
  reg [7:0] phv_data_389; // @[executor.scala 448:22]
  reg [7:0] phv_data_390; // @[executor.scala 448:22]
  reg [7:0] phv_data_391; // @[executor.scala 448:22]
  reg [7:0] phv_data_392; // @[executor.scala 448:22]
  reg [7:0] phv_data_393; // @[executor.scala 448:22]
  reg [7:0] phv_data_394; // @[executor.scala 448:22]
  reg [7:0] phv_data_395; // @[executor.scala 448:22]
  reg [7:0] phv_data_396; // @[executor.scala 448:22]
  reg [7:0] phv_data_397; // @[executor.scala 448:22]
  reg [7:0] phv_data_398; // @[executor.scala 448:22]
  reg [7:0] phv_data_399; // @[executor.scala 448:22]
  reg [7:0] phv_data_400; // @[executor.scala 448:22]
  reg [7:0] phv_data_401; // @[executor.scala 448:22]
  reg [7:0] phv_data_402; // @[executor.scala 448:22]
  reg [7:0] phv_data_403; // @[executor.scala 448:22]
  reg [7:0] phv_data_404; // @[executor.scala 448:22]
  reg [7:0] phv_data_405; // @[executor.scala 448:22]
  reg [7:0] phv_data_406; // @[executor.scala 448:22]
  reg [7:0] phv_data_407; // @[executor.scala 448:22]
  reg [7:0] phv_data_408; // @[executor.scala 448:22]
  reg [7:0] phv_data_409; // @[executor.scala 448:22]
  reg [7:0] phv_data_410; // @[executor.scala 448:22]
  reg [7:0] phv_data_411; // @[executor.scala 448:22]
  reg [7:0] phv_data_412; // @[executor.scala 448:22]
  reg [7:0] phv_data_413; // @[executor.scala 448:22]
  reg [7:0] phv_data_414; // @[executor.scala 448:22]
  reg [7:0] phv_data_415; // @[executor.scala 448:22]
  reg [7:0] phv_data_416; // @[executor.scala 448:22]
  reg [7:0] phv_data_417; // @[executor.scala 448:22]
  reg [7:0] phv_data_418; // @[executor.scala 448:22]
  reg [7:0] phv_data_419; // @[executor.scala 448:22]
  reg [7:0] phv_data_420; // @[executor.scala 448:22]
  reg [7:0] phv_data_421; // @[executor.scala 448:22]
  reg [7:0] phv_data_422; // @[executor.scala 448:22]
  reg [7:0] phv_data_423; // @[executor.scala 448:22]
  reg [7:0] phv_data_424; // @[executor.scala 448:22]
  reg [7:0] phv_data_425; // @[executor.scala 448:22]
  reg [7:0] phv_data_426; // @[executor.scala 448:22]
  reg [7:0] phv_data_427; // @[executor.scala 448:22]
  reg [7:0] phv_data_428; // @[executor.scala 448:22]
  reg [7:0] phv_data_429; // @[executor.scala 448:22]
  reg [7:0] phv_data_430; // @[executor.scala 448:22]
  reg [7:0] phv_data_431; // @[executor.scala 448:22]
  reg [7:0] phv_data_432; // @[executor.scala 448:22]
  reg [7:0] phv_data_433; // @[executor.scala 448:22]
  reg [7:0] phv_data_434; // @[executor.scala 448:22]
  reg [7:0] phv_data_435; // @[executor.scala 448:22]
  reg [7:0] phv_data_436; // @[executor.scala 448:22]
  reg [7:0] phv_data_437; // @[executor.scala 448:22]
  reg [7:0] phv_data_438; // @[executor.scala 448:22]
  reg [7:0] phv_data_439; // @[executor.scala 448:22]
  reg [7:0] phv_data_440; // @[executor.scala 448:22]
  reg [7:0] phv_data_441; // @[executor.scala 448:22]
  reg [7:0] phv_data_442; // @[executor.scala 448:22]
  reg [7:0] phv_data_443; // @[executor.scala 448:22]
  reg [7:0] phv_data_444; // @[executor.scala 448:22]
  reg [7:0] phv_data_445; // @[executor.scala 448:22]
  reg [7:0] phv_data_446; // @[executor.scala 448:22]
  reg [7:0] phv_data_447; // @[executor.scala 448:22]
  reg [7:0] phv_data_448; // @[executor.scala 448:22]
  reg [7:0] phv_data_449; // @[executor.scala 448:22]
  reg [7:0] phv_data_450; // @[executor.scala 448:22]
  reg [7:0] phv_data_451; // @[executor.scala 448:22]
  reg [7:0] phv_data_452; // @[executor.scala 448:22]
  reg [7:0] phv_data_453; // @[executor.scala 448:22]
  reg [7:0] phv_data_454; // @[executor.scala 448:22]
  reg [7:0] phv_data_455; // @[executor.scala 448:22]
  reg [7:0] phv_data_456; // @[executor.scala 448:22]
  reg [7:0] phv_data_457; // @[executor.scala 448:22]
  reg [7:0] phv_data_458; // @[executor.scala 448:22]
  reg [7:0] phv_data_459; // @[executor.scala 448:22]
  reg [7:0] phv_data_460; // @[executor.scala 448:22]
  reg [7:0] phv_data_461; // @[executor.scala 448:22]
  reg [7:0] phv_data_462; // @[executor.scala 448:22]
  reg [7:0] phv_data_463; // @[executor.scala 448:22]
  reg [7:0] phv_data_464; // @[executor.scala 448:22]
  reg [7:0] phv_data_465; // @[executor.scala 448:22]
  reg [7:0] phv_data_466; // @[executor.scala 448:22]
  reg [7:0] phv_data_467; // @[executor.scala 448:22]
  reg [7:0] phv_data_468; // @[executor.scala 448:22]
  reg [7:0] phv_data_469; // @[executor.scala 448:22]
  reg [7:0] phv_data_470; // @[executor.scala 448:22]
  reg [7:0] phv_data_471; // @[executor.scala 448:22]
  reg [7:0] phv_data_472; // @[executor.scala 448:22]
  reg [7:0] phv_data_473; // @[executor.scala 448:22]
  reg [7:0] phv_data_474; // @[executor.scala 448:22]
  reg [7:0] phv_data_475; // @[executor.scala 448:22]
  reg [7:0] phv_data_476; // @[executor.scala 448:22]
  reg [7:0] phv_data_477; // @[executor.scala 448:22]
  reg [7:0] phv_data_478; // @[executor.scala 448:22]
  reg [7:0] phv_data_479; // @[executor.scala 448:22]
  reg [7:0] phv_data_480; // @[executor.scala 448:22]
  reg [7:0] phv_data_481; // @[executor.scala 448:22]
  reg [7:0] phv_data_482; // @[executor.scala 448:22]
  reg [7:0] phv_data_483; // @[executor.scala 448:22]
  reg [7:0] phv_data_484; // @[executor.scala 448:22]
  reg [7:0] phv_data_485; // @[executor.scala 448:22]
  reg [7:0] phv_data_486; // @[executor.scala 448:22]
  reg [7:0] phv_data_487; // @[executor.scala 448:22]
  reg [7:0] phv_data_488; // @[executor.scala 448:22]
  reg [7:0] phv_data_489; // @[executor.scala 448:22]
  reg [7:0] phv_data_490; // @[executor.scala 448:22]
  reg [7:0] phv_data_491; // @[executor.scala 448:22]
  reg [7:0] phv_data_492; // @[executor.scala 448:22]
  reg [7:0] phv_data_493; // @[executor.scala 448:22]
  reg [7:0] phv_data_494; // @[executor.scala 448:22]
  reg [7:0] phv_data_495; // @[executor.scala 448:22]
  reg [7:0] phv_data_496; // @[executor.scala 448:22]
  reg [7:0] phv_data_497; // @[executor.scala 448:22]
  reg [7:0] phv_data_498; // @[executor.scala 448:22]
  reg [7:0] phv_data_499; // @[executor.scala 448:22]
  reg [7:0] phv_data_500; // @[executor.scala 448:22]
  reg [7:0] phv_data_501; // @[executor.scala 448:22]
  reg [7:0] phv_data_502; // @[executor.scala 448:22]
  reg [7:0] phv_data_503; // @[executor.scala 448:22]
  reg [7:0] phv_data_504; // @[executor.scala 448:22]
  reg [7:0] phv_data_505; // @[executor.scala 448:22]
  reg [7:0] phv_data_506; // @[executor.scala 448:22]
  reg [7:0] phv_data_507; // @[executor.scala 448:22]
  reg [7:0] phv_data_508; // @[executor.scala 448:22]
  reg [7:0] phv_data_509; // @[executor.scala 448:22]
  reg [7:0] phv_data_510; // @[executor.scala 448:22]
  reg [7:0] phv_data_511; // @[executor.scala 448:22]
  reg [15:0] phv_header_0; // @[executor.scala 448:22]
  reg [15:0] phv_header_1; // @[executor.scala 448:22]
  reg [15:0] phv_header_2; // @[executor.scala 448:22]
  reg [15:0] phv_header_3; // @[executor.scala 448:22]
  reg [15:0] phv_header_4; // @[executor.scala 448:22]
  reg [15:0] phv_header_5; // @[executor.scala 448:22]
  reg [15:0] phv_header_6; // @[executor.scala 448:22]
  reg [15:0] phv_header_7; // @[executor.scala 448:22]
  reg [15:0] phv_header_8; // @[executor.scala 448:22]
  reg [15:0] phv_header_9; // @[executor.scala 448:22]
  reg [15:0] phv_header_10; // @[executor.scala 448:22]
  reg [15:0] phv_header_11; // @[executor.scala 448:22]
  reg [15:0] phv_header_12; // @[executor.scala 448:22]
  reg [15:0] phv_header_13; // @[executor.scala 448:22]
  reg [15:0] phv_header_14; // @[executor.scala 448:22]
  reg [15:0] phv_header_15; // @[executor.scala 448:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 448:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 448:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 448:22]
  reg [3:0] phv_next_processor_id; // @[executor.scala 448:22]
  reg  phv_next_config_id; // @[executor.scala 448:22]
  reg  phv_is_valid_processor; // @[executor.scala 448:22]
  reg [31:0] vliw_0; // @[executor.scala 452:23]
  reg [31:0] vliw_1; // @[executor.scala 452:23]
  reg [31:0] vliw_2; // @[executor.scala 452:23]
  reg [31:0] vliw_3; // @[executor.scala 452:23]
  reg [31:0] field_0; // @[executor.scala 454:24]
  reg [31:0] field_1; // @[executor.scala 454:24]
  reg [31:0] field_2; // @[executor.scala 454:24]
  reg [31:0] field_3; // @[executor.scala 454:24]
  reg [3:0] mask_0; // @[executor.scala 456:23]
  reg [3:0] mask_1; // @[executor.scala 456:23]
  reg [3:0] mask_2; // @[executor.scala 456:23]
  reg [3:0] mask_3; // @[executor.scala 456:23]
  reg [5:0] dst_offset_0; // @[executor.scala 458:29]
  reg [5:0] dst_offset_1; // @[executor.scala 458:29]
  reg [5:0] dst_offset_2; // @[executor.scala 458:29]
  reg [5:0] dst_offset_3; // @[executor.scala 458:29]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2 = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8714 = {{2'd0}, dst_offset_0}; // @[executor.scala 473:49]
  wire [7:0] byte_ = field_0[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_0 = mask_0[0] ? byte_ : phv_data_3; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_1 = field_0[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_1 = mask_0[1] ? byte_1 : phv_data_2; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_2 = field_0[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2 = mask_0[2] ? byte_2 : phv_data_1; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] byte_3 = field_0[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_3 = mask_0[3] ? byte_3 : phv_data_0; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_4 = _GEN_8714 == 8'h0 ? _GEN_0 : phv_data_3; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_5 = _GEN_8714 == 8'h0 ? _GEN_1 : phv_data_2; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_6 = _GEN_8714 == 8'h0 ? _GEN_2 : phv_data_1; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_7 = _GEN_8714 == 8'h0 ? _GEN_3 : phv_data_0; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_8 = mask_0[0] ? byte_ : phv_data_7; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_9 = mask_0[1] ? byte_1 : phv_data_6; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_10 = mask_0[2] ? byte_2 : phv_data_5; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_11 = mask_0[3] ? byte_3 : phv_data_4; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_12 = _GEN_8714 == 8'h1 ? _GEN_8 : phv_data_7; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_13 = _GEN_8714 == 8'h1 ? _GEN_9 : phv_data_6; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_14 = _GEN_8714 == 8'h1 ? _GEN_10 : phv_data_5; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_15 = _GEN_8714 == 8'h1 ? _GEN_11 : phv_data_4; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_16 = mask_0[0] ? byte_ : phv_data_11; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_17 = mask_0[1] ? byte_1 : phv_data_10; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_18 = mask_0[2] ? byte_2 : phv_data_9; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_19 = mask_0[3] ? byte_3 : phv_data_8; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_20 = _GEN_8714 == 8'h2 ? _GEN_16 : phv_data_11; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_21 = _GEN_8714 == 8'h2 ? _GEN_17 : phv_data_10; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_22 = _GEN_8714 == 8'h2 ? _GEN_18 : phv_data_9; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_23 = _GEN_8714 == 8'h2 ? _GEN_19 : phv_data_8; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_24 = mask_0[0] ? byte_ : phv_data_15; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_25 = mask_0[1] ? byte_1 : phv_data_14; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_26 = mask_0[2] ? byte_2 : phv_data_13; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_27 = mask_0[3] ? byte_3 : phv_data_12; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_28 = _GEN_8714 == 8'h3 ? _GEN_24 : phv_data_15; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_29 = _GEN_8714 == 8'h3 ? _GEN_25 : phv_data_14; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_30 = _GEN_8714 == 8'h3 ? _GEN_26 : phv_data_13; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_31 = _GEN_8714 == 8'h3 ? _GEN_27 : phv_data_12; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_32 = mask_0[0] ? byte_ : phv_data_19; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_33 = mask_0[1] ? byte_1 : phv_data_18; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_34 = mask_0[2] ? byte_2 : phv_data_17; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_35 = mask_0[3] ? byte_3 : phv_data_16; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_36 = _GEN_8714 == 8'h4 ? _GEN_32 : phv_data_19; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_37 = _GEN_8714 == 8'h4 ? _GEN_33 : phv_data_18; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_38 = _GEN_8714 == 8'h4 ? _GEN_34 : phv_data_17; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_39 = _GEN_8714 == 8'h4 ? _GEN_35 : phv_data_16; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_40 = mask_0[0] ? byte_ : phv_data_23; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_41 = mask_0[1] ? byte_1 : phv_data_22; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_42 = mask_0[2] ? byte_2 : phv_data_21; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_43 = mask_0[3] ? byte_3 : phv_data_20; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_44 = _GEN_8714 == 8'h5 ? _GEN_40 : phv_data_23; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_45 = _GEN_8714 == 8'h5 ? _GEN_41 : phv_data_22; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_46 = _GEN_8714 == 8'h5 ? _GEN_42 : phv_data_21; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_47 = _GEN_8714 == 8'h5 ? _GEN_43 : phv_data_20; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_48 = mask_0[0] ? byte_ : phv_data_27; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_49 = mask_0[1] ? byte_1 : phv_data_26; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_50 = mask_0[2] ? byte_2 : phv_data_25; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_51 = mask_0[3] ? byte_3 : phv_data_24; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_52 = _GEN_8714 == 8'h6 ? _GEN_48 : phv_data_27; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_53 = _GEN_8714 == 8'h6 ? _GEN_49 : phv_data_26; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_54 = _GEN_8714 == 8'h6 ? _GEN_50 : phv_data_25; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_55 = _GEN_8714 == 8'h6 ? _GEN_51 : phv_data_24; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_56 = mask_0[0] ? byte_ : phv_data_31; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_57 = mask_0[1] ? byte_1 : phv_data_30; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_58 = mask_0[2] ? byte_2 : phv_data_29; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_59 = mask_0[3] ? byte_3 : phv_data_28; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_60 = _GEN_8714 == 8'h7 ? _GEN_56 : phv_data_31; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_61 = _GEN_8714 == 8'h7 ? _GEN_57 : phv_data_30; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_62 = _GEN_8714 == 8'h7 ? _GEN_58 : phv_data_29; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_63 = _GEN_8714 == 8'h7 ? _GEN_59 : phv_data_28; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_64 = mask_0[0] ? byte_ : phv_data_35; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_65 = mask_0[1] ? byte_1 : phv_data_34; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_66 = mask_0[2] ? byte_2 : phv_data_33; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_67 = mask_0[3] ? byte_3 : phv_data_32; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_68 = _GEN_8714 == 8'h8 ? _GEN_64 : phv_data_35; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_69 = _GEN_8714 == 8'h8 ? _GEN_65 : phv_data_34; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_70 = _GEN_8714 == 8'h8 ? _GEN_66 : phv_data_33; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_71 = _GEN_8714 == 8'h8 ? _GEN_67 : phv_data_32; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_72 = mask_0[0] ? byte_ : phv_data_39; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_73 = mask_0[1] ? byte_1 : phv_data_38; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_74 = mask_0[2] ? byte_2 : phv_data_37; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_75 = mask_0[3] ? byte_3 : phv_data_36; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_76 = _GEN_8714 == 8'h9 ? _GEN_72 : phv_data_39; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_77 = _GEN_8714 == 8'h9 ? _GEN_73 : phv_data_38; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_78 = _GEN_8714 == 8'h9 ? _GEN_74 : phv_data_37; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_79 = _GEN_8714 == 8'h9 ? _GEN_75 : phv_data_36; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_80 = mask_0[0] ? byte_ : phv_data_43; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_81 = mask_0[1] ? byte_1 : phv_data_42; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_82 = mask_0[2] ? byte_2 : phv_data_41; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_83 = mask_0[3] ? byte_3 : phv_data_40; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_84 = _GEN_8714 == 8'ha ? _GEN_80 : phv_data_43; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_85 = _GEN_8714 == 8'ha ? _GEN_81 : phv_data_42; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_86 = _GEN_8714 == 8'ha ? _GEN_82 : phv_data_41; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_87 = _GEN_8714 == 8'ha ? _GEN_83 : phv_data_40; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_88 = mask_0[0] ? byte_ : phv_data_47; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_89 = mask_0[1] ? byte_1 : phv_data_46; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_90 = mask_0[2] ? byte_2 : phv_data_45; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_91 = mask_0[3] ? byte_3 : phv_data_44; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_92 = _GEN_8714 == 8'hb ? _GEN_88 : phv_data_47; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_93 = _GEN_8714 == 8'hb ? _GEN_89 : phv_data_46; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_94 = _GEN_8714 == 8'hb ? _GEN_90 : phv_data_45; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_95 = _GEN_8714 == 8'hb ? _GEN_91 : phv_data_44; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_96 = mask_0[0] ? byte_ : phv_data_51; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_97 = mask_0[1] ? byte_1 : phv_data_50; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_98 = mask_0[2] ? byte_2 : phv_data_49; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_99 = mask_0[3] ? byte_3 : phv_data_48; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_100 = _GEN_8714 == 8'hc ? _GEN_96 : phv_data_51; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_101 = _GEN_8714 == 8'hc ? _GEN_97 : phv_data_50; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_102 = _GEN_8714 == 8'hc ? _GEN_98 : phv_data_49; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_103 = _GEN_8714 == 8'hc ? _GEN_99 : phv_data_48; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_104 = mask_0[0] ? byte_ : phv_data_55; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_105 = mask_0[1] ? byte_1 : phv_data_54; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_106 = mask_0[2] ? byte_2 : phv_data_53; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_107 = mask_0[3] ? byte_3 : phv_data_52; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_108 = _GEN_8714 == 8'hd ? _GEN_104 : phv_data_55; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_109 = _GEN_8714 == 8'hd ? _GEN_105 : phv_data_54; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_110 = _GEN_8714 == 8'hd ? _GEN_106 : phv_data_53; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_111 = _GEN_8714 == 8'hd ? _GEN_107 : phv_data_52; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_112 = mask_0[0] ? byte_ : phv_data_59; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_113 = mask_0[1] ? byte_1 : phv_data_58; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_114 = mask_0[2] ? byte_2 : phv_data_57; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_115 = mask_0[3] ? byte_3 : phv_data_56; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_116 = _GEN_8714 == 8'he ? _GEN_112 : phv_data_59; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_117 = _GEN_8714 == 8'he ? _GEN_113 : phv_data_58; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_118 = _GEN_8714 == 8'he ? _GEN_114 : phv_data_57; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_119 = _GEN_8714 == 8'he ? _GEN_115 : phv_data_56; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_120 = mask_0[0] ? byte_ : phv_data_63; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_121 = mask_0[1] ? byte_1 : phv_data_62; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_122 = mask_0[2] ? byte_2 : phv_data_61; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_123 = mask_0[3] ? byte_3 : phv_data_60; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_124 = _GEN_8714 == 8'hf ? _GEN_120 : phv_data_63; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_125 = _GEN_8714 == 8'hf ? _GEN_121 : phv_data_62; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_126 = _GEN_8714 == 8'hf ? _GEN_122 : phv_data_61; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_127 = _GEN_8714 == 8'hf ? _GEN_123 : phv_data_60; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_128 = mask_0[0] ? byte_ : phv_data_67; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_129 = mask_0[1] ? byte_1 : phv_data_66; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_130 = mask_0[2] ? byte_2 : phv_data_65; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_131 = mask_0[3] ? byte_3 : phv_data_64; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_132 = _GEN_8714 == 8'h10 ? _GEN_128 : phv_data_67; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_133 = _GEN_8714 == 8'h10 ? _GEN_129 : phv_data_66; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_134 = _GEN_8714 == 8'h10 ? _GEN_130 : phv_data_65; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_135 = _GEN_8714 == 8'h10 ? _GEN_131 : phv_data_64; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_136 = mask_0[0] ? byte_ : phv_data_71; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_137 = mask_0[1] ? byte_1 : phv_data_70; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_138 = mask_0[2] ? byte_2 : phv_data_69; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_139 = mask_0[3] ? byte_3 : phv_data_68; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_140 = _GEN_8714 == 8'h11 ? _GEN_136 : phv_data_71; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_141 = _GEN_8714 == 8'h11 ? _GEN_137 : phv_data_70; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_142 = _GEN_8714 == 8'h11 ? _GEN_138 : phv_data_69; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_143 = _GEN_8714 == 8'h11 ? _GEN_139 : phv_data_68; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_144 = mask_0[0] ? byte_ : phv_data_75; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_145 = mask_0[1] ? byte_1 : phv_data_74; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_146 = mask_0[2] ? byte_2 : phv_data_73; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_147 = mask_0[3] ? byte_3 : phv_data_72; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_148 = _GEN_8714 == 8'h12 ? _GEN_144 : phv_data_75; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_149 = _GEN_8714 == 8'h12 ? _GEN_145 : phv_data_74; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_150 = _GEN_8714 == 8'h12 ? _GEN_146 : phv_data_73; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_151 = _GEN_8714 == 8'h12 ? _GEN_147 : phv_data_72; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_152 = mask_0[0] ? byte_ : phv_data_79; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_153 = mask_0[1] ? byte_1 : phv_data_78; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_154 = mask_0[2] ? byte_2 : phv_data_77; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_155 = mask_0[3] ? byte_3 : phv_data_76; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_156 = _GEN_8714 == 8'h13 ? _GEN_152 : phv_data_79; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_157 = _GEN_8714 == 8'h13 ? _GEN_153 : phv_data_78; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_158 = _GEN_8714 == 8'h13 ? _GEN_154 : phv_data_77; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_159 = _GEN_8714 == 8'h13 ? _GEN_155 : phv_data_76; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_160 = mask_0[0] ? byte_ : phv_data_83; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_161 = mask_0[1] ? byte_1 : phv_data_82; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_162 = mask_0[2] ? byte_2 : phv_data_81; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_163 = mask_0[3] ? byte_3 : phv_data_80; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_164 = _GEN_8714 == 8'h14 ? _GEN_160 : phv_data_83; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_165 = _GEN_8714 == 8'h14 ? _GEN_161 : phv_data_82; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_166 = _GEN_8714 == 8'h14 ? _GEN_162 : phv_data_81; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_167 = _GEN_8714 == 8'h14 ? _GEN_163 : phv_data_80; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_168 = mask_0[0] ? byte_ : phv_data_87; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_169 = mask_0[1] ? byte_1 : phv_data_86; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_170 = mask_0[2] ? byte_2 : phv_data_85; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_171 = mask_0[3] ? byte_3 : phv_data_84; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_172 = _GEN_8714 == 8'h15 ? _GEN_168 : phv_data_87; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_173 = _GEN_8714 == 8'h15 ? _GEN_169 : phv_data_86; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_174 = _GEN_8714 == 8'h15 ? _GEN_170 : phv_data_85; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_175 = _GEN_8714 == 8'h15 ? _GEN_171 : phv_data_84; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_176 = mask_0[0] ? byte_ : phv_data_91; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_177 = mask_0[1] ? byte_1 : phv_data_90; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_178 = mask_0[2] ? byte_2 : phv_data_89; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_179 = mask_0[3] ? byte_3 : phv_data_88; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_180 = _GEN_8714 == 8'h16 ? _GEN_176 : phv_data_91; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_181 = _GEN_8714 == 8'h16 ? _GEN_177 : phv_data_90; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_182 = _GEN_8714 == 8'h16 ? _GEN_178 : phv_data_89; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_183 = _GEN_8714 == 8'h16 ? _GEN_179 : phv_data_88; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_184 = mask_0[0] ? byte_ : phv_data_95; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_185 = mask_0[1] ? byte_1 : phv_data_94; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_186 = mask_0[2] ? byte_2 : phv_data_93; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_187 = mask_0[3] ? byte_3 : phv_data_92; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_188 = _GEN_8714 == 8'h17 ? _GEN_184 : phv_data_95; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_189 = _GEN_8714 == 8'h17 ? _GEN_185 : phv_data_94; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_190 = _GEN_8714 == 8'h17 ? _GEN_186 : phv_data_93; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_191 = _GEN_8714 == 8'h17 ? _GEN_187 : phv_data_92; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_192 = mask_0[0] ? byte_ : phv_data_99; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_193 = mask_0[1] ? byte_1 : phv_data_98; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_194 = mask_0[2] ? byte_2 : phv_data_97; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_195 = mask_0[3] ? byte_3 : phv_data_96; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_196 = _GEN_8714 == 8'h18 ? _GEN_192 : phv_data_99; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_197 = _GEN_8714 == 8'h18 ? _GEN_193 : phv_data_98; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_198 = _GEN_8714 == 8'h18 ? _GEN_194 : phv_data_97; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_199 = _GEN_8714 == 8'h18 ? _GEN_195 : phv_data_96; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_200 = mask_0[0] ? byte_ : phv_data_103; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_201 = mask_0[1] ? byte_1 : phv_data_102; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_202 = mask_0[2] ? byte_2 : phv_data_101; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_203 = mask_0[3] ? byte_3 : phv_data_100; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_204 = _GEN_8714 == 8'h19 ? _GEN_200 : phv_data_103; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_205 = _GEN_8714 == 8'h19 ? _GEN_201 : phv_data_102; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_206 = _GEN_8714 == 8'h19 ? _GEN_202 : phv_data_101; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_207 = _GEN_8714 == 8'h19 ? _GEN_203 : phv_data_100; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_208 = mask_0[0] ? byte_ : phv_data_107; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_209 = mask_0[1] ? byte_1 : phv_data_106; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_210 = mask_0[2] ? byte_2 : phv_data_105; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_211 = mask_0[3] ? byte_3 : phv_data_104; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_212 = _GEN_8714 == 8'h1a ? _GEN_208 : phv_data_107; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_213 = _GEN_8714 == 8'h1a ? _GEN_209 : phv_data_106; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_214 = _GEN_8714 == 8'h1a ? _GEN_210 : phv_data_105; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_215 = _GEN_8714 == 8'h1a ? _GEN_211 : phv_data_104; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_216 = mask_0[0] ? byte_ : phv_data_111; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_217 = mask_0[1] ? byte_1 : phv_data_110; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_218 = mask_0[2] ? byte_2 : phv_data_109; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_219 = mask_0[3] ? byte_3 : phv_data_108; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_220 = _GEN_8714 == 8'h1b ? _GEN_216 : phv_data_111; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_221 = _GEN_8714 == 8'h1b ? _GEN_217 : phv_data_110; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_222 = _GEN_8714 == 8'h1b ? _GEN_218 : phv_data_109; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_223 = _GEN_8714 == 8'h1b ? _GEN_219 : phv_data_108; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_224 = mask_0[0] ? byte_ : phv_data_115; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_225 = mask_0[1] ? byte_1 : phv_data_114; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_226 = mask_0[2] ? byte_2 : phv_data_113; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_227 = mask_0[3] ? byte_3 : phv_data_112; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_228 = _GEN_8714 == 8'h1c ? _GEN_224 : phv_data_115; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_229 = _GEN_8714 == 8'h1c ? _GEN_225 : phv_data_114; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_230 = _GEN_8714 == 8'h1c ? _GEN_226 : phv_data_113; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_231 = _GEN_8714 == 8'h1c ? _GEN_227 : phv_data_112; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_232 = mask_0[0] ? byte_ : phv_data_119; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_233 = mask_0[1] ? byte_1 : phv_data_118; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_234 = mask_0[2] ? byte_2 : phv_data_117; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_235 = mask_0[3] ? byte_3 : phv_data_116; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_236 = _GEN_8714 == 8'h1d ? _GEN_232 : phv_data_119; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_237 = _GEN_8714 == 8'h1d ? _GEN_233 : phv_data_118; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_238 = _GEN_8714 == 8'h1d ? _GEN_234 : phv_data_117; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_239 = _GEN_8714 == 8'h1d ? _GEN_235 : phv_data_116; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_240 = mask_0[0] ? byte_ : phv_data_123; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_241 = mask_0[1] ? byte_1 : phv_data_122; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_242 = mask_0[2] ? byte_2 : phv_data_121; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_243 = mask_0[3] ? byte_3 : phv_data_120; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_244 = _GEN_8714 == 8'h1e ? _GEN_240 : phv_data_123; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_245 = _GEN_8714 == 8'h1e ? _GEN_241 : phv_data_122; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_246 = _GEN_8714 == 8'h1e ? _GEN_242 : phv_data_121; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_247 = _GEN_8714 == 8'h1e ? _GEN_243 : phv_data_120; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_248 = mask_0[0] ? byte_ : phv_data_127; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_249 = mask_0[1] ? byte_1 : phv_data_126; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_250 = mask_0[2] ? byte_2 : phv_data_125; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_251 = mask_0[3] ? byte_3 : phv_data_124; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_252 = _GEN_8714 == 8'h1f ? _GEN_248 : phv_data_127; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_253 = _GEN_8714 == 8'h1f ? _GEN_249 : phv_data_126; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_254 = _GEN_8714 == 8'h1f ? _GEN_250 : phv_data_125; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_255 = _GEN_8714 == 8'h1f ? _GEN_251 : phv_data_124; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_256 = mask_0[0] ? byte_ : phv_data_131; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_257 = mask_0[1] ? byte_1 : phv_data_130; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_258 = mask_0[2] ? byte_2 : phv_data_129; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_259 = mask_0[3] ? byte_3 : phv_data_128; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_260 = _GEN_8714 == 8'h20 ? _GEN_256 : phv_data_131; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_261 = _GEN_8714 == 8'h20 ? _GEN_257 : phv_data_130; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_262 = _GEN_8714 == 8'h20 ? _GEN_258 : phv_data_129; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_263 = _GEN_8714 == 8'h20 ? _GEN_259 : phv_data_128; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_264 = mask_0[0] ? byte_ : phv_data_135; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_265 = mask_0[1] ? byte_1 : phv_data_134; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_266 = mask_0[2] ? byte_2 : phv_data_133; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_267 = mask_0[3] ? byte_3 : phv_data_132; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_268 = _GEN_8714 == 8'h21 ? _GEN_264 : phv_data_135; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_269 = _GEN_8714 == 8'h21 ? _GEN_265 : phv_data_134; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_270 = _GEN_8714 == 8'h21 ? _GEN_266 : phv_data_133; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_271 = _GEN_8714 == 8'h21 ? _GEN_267 : phv_data_132; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_272 = mask_0[0] ? byte_ : phv_data_139; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_273 = mask_0[1] ? byte_1 : phv_data_138; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_274 = mask_0[2] ? byte_2 : phv_data_137; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_275 = mask_0[3] ? byte_3 : phv_data_136; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_276 = _GEN_8714 == 8'h22 ? _GEN_272 : phv_data_139; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_277 = _GEN_8714 == 8'h22 ? _GEN_273 : phv_data_138; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_278 = _GEN_8714 == 8'h22 ? _GEN_274 : phv_data_137; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_279 = _GEN_8714 == 8'h22 ? _GEN_275 : phv_data_136; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_280 = mask_0[0] ? byte_ : phv_data_143; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_281 = mask_0[1] ? byte_1 : phv_data_142; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_282 = mask_0[2] ? byte_2 : phv_data_141; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_283 = mask_0[3] ? byte_3 : phv_data_140; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_284 = _GEN_8714 == 8'h23 ? _GEN_280 : phv_data_143; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_285 = _GEN_8714 == 8'h23 ? _GEN_281 : phv_data_142; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_286 = _GEN_8714 == 8'h23 ? _GEN_282 : phv_data_141; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_287 = _GEN_8714 == 8'h23 ? _GEN_283 : phv_data_140; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_288 = mask_0[0] ? byte_ : phv_data_147; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_289 = mask_0[1] ? byte_1 : phv_data_146; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_290 = mask_0[2] ? byte_2 : phv_data_145; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_291 = mask_0[3] ? byte_3 : phv_data_144; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_292 = _GEN_8714 == 8'h24 ? _GEN_288 : phv_data_147; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_293 = _GEN_8714 == 8'h24 ? _GEN_289 : phv_data_146; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_294 = _GEN_8714 == 8'h24 ? _GEN_290 : phv_data_145; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_295 = _GEN_8714 == 8'h24 ? _GEN_291 : phv_data_144; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_296 = mask_0[0] ? byte_ : phv_data_151; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_297 = mask_0[1] ? byte_1 : phv_data_150; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_298 = mask_0[2] ? byte_2 : phv_data_149; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_299 = mask_0[3] ? byte_3 : phv_data_148; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_300 = _GEN_8714 == 8'h25 ? _GEN_296 : phv_data_151; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_301 = _GEN_8714 == 8'h25 ? _GEN_297 : phv_data_150; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_302 = _GEN_8714 == 8'h25 ? _GEN_298 : phv_data_149; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_303 = _GEN_8714 == 8'h25 ? _GEN_299 : phv_data_148; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_304 = mask_0[0] ? byte_ : phv_data_155; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_305 = mask_0[1] ? byte_1 : phv_data_154; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_306 = mask_0[2] ? byte_2 : phv_data_153; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_307 = mask_0[3] ? byte_3 : phv_data_152; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_308 = _GEN_8714 == 8'h26 ? _GEN_304 : phv_data_155; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_309 = _GEN_8714 == 8'h26 ? _GEN_305 : phv_data_154; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_310 = _GEN_8714 == 8'h26 ? _GEN_306 : phv_data_153; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_311 = _GEN_8714 == 8'h26 ? _GEN_307 : phv_data_152; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_312 = mask_0[0] ? byte_ : phv_data_159; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_313 = mask_0[1] ? byte_1 : phv_data_158; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_314 = mask_0[2] ? byte_2 : phv_data_157; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_315 = mask_0[3] ? byte_3 : phv_data_156; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_316 = _GEN_8714 == 8'h27 ? _GEN_312 : phv_data_159; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_317 = _GEN_8714 == 8'h27 ? _GEN_313 : phv_data_158; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_318 = _GEN_8714 == 8'h27 ? _GEN_314 : phv_data_157; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_319 = _GEN_8714 == 8'h27 ? _GEN_315 : phv_data_156; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_320 = mask_0[0] ? byte_ : phv_data_163; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_321 = mask_0[1] ? byte_1 : phv_data_162; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_322 = mask_0[2] ? byte_2 : phv_data_161; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_323 = mask_0[3] ? byte_3 : phv_data_160; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_324 = _GEN_8714 == 8'h28 ? _GEN_320 : phv_data_163; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_325 = _GEN_8714 == 8'h28 ? _GEN_321 : phv_data_162; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_326 = _GEN_8714 == 8'h28 ? _GEN_322 : phv_data_161; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_327 = _GEN_8714 == 8'h28 ? _GEN_323 : phv_data_160; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_328 = mask_0[0] ? byte_ : phv_data_167; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_329 = mask_0[1] ? byte_1 : phv_data_166; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_330 = mask_0[2] ? byte_2 : phv_data_165; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_331 = mask_0[3] ? byte_3 : phv_data_164; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_332 = _GEN_8714 == 8'h29 ? _GEN_328 : phv_data_167; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_333 = _GEN_8714 == 8'h29 ? _GEN_329 : phv_data_166; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_334 = _GEN_8714 == 8'h29 ? _GEN_330 : phv_data_165; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_335 = _GEN_8714 == 8'h29 ? _GEN_331 : phv_data_164; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_336 = mask_0[0] ? byte_ : phv_data_171; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_337 = mask_0[1] ? byte_1 : phv_data_170; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_338 = mask_0[2] ? byte_2 : phv_data_169; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_339 = mask_0[3] ? byte_3 : phv_data_168; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_340 = _GEN_8714 == 8'h2a ? _GEN_336 : phv_data_171; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_341 = _GEN_8714 == 8'h2a ? _GEN_337 : phv_data_170; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_342 = _GEN_8714 == 8'h2a ? _GEN_338 : phv_data_169; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_343 = _GEN_8714 == 8'h2a ? _GEN_339 : phv_data_168; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_344 = mask_0[0] ? byte_ : phv_data_175; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_345 = mask_0[1] ? byte_1 : phv_data_174; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_346 = mask_0[2] ? byte_2 : phv_data_173; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_347 = mask_0[3] ? byte_3 : phv_data_172; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_348 = _GEN_8714 == 8'h2b ? _GEN_344 : phv_data_175; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_349 = _GEN_8714 == 8'h2b ? _GEN_345 : phv_data_174; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_350 = _GEN_8714 == 8'h2b ? _GEN_346 : phv_data_173; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_351 = _GEN_8714 == 8'h2b ? _GEN_347 : phv_data_172; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_352 = mask_0[0] ? byte_ : phv_data_179; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_353 = mask_0[1] ? byte_1 : phv_data_178; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_354 = mask_0[2] ? byte_2 : phv_data_177; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_355 = mask_0[3] ? byte_3 : phv_data_176; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_356 = _GEN_8714 == 8'h2c ? _GEN_352 : phv_data_179; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_357 = _GEN_8714 == 8'h2c ? _GEN_353 : phv_data_178; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_358 = _GEN_8714 == 8'h2c ? _GEN_354 : phv_data_177; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_359 = _GEN_8714 == 8'h2c ? _GEN_355 : phv_data_176; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_360 = mask_0[0] ? byte_ : phv_data_183; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_361 = mask_0[1] ? byte_1 : phv_data_182; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_362 = mask_0[2] ? byte_2 : phv_data_181; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_363 = mask_0[3] ? byte_3 : phv_data_180; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_364 = _GEN_8714 == 8'h2d ? _GEN_360 : phv_data_183; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_365 = _GEN_8714 == 8'h2d ? _GEN_361 : phv_data_182; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_366 = _GEN_8714 == 8'h2d ? _GEN_362 : phv_data_181; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_367 = _GEN_8714 == 8'h2d ? _GEN_363 : phv_data_180; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_368 = mask_0[0] ? byte_ : phv_data_187; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_369 = mask_0[1] ? byte_1 : phv_data_186; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_370 = mask_0[2] ? byte_2 : phv_data_185; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_371 = mask_0[3] ? byte_3 : phv_data_184; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_372 = _GEN_8714 == 8'h2e ? _GEN_368 : phv_data_187; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_373 = _GEN_8714 == 8'h2e ? _GEN_369 : phv_data_186; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_374 = _GEN_8714 == 8'h2e ? _GEN_370 : phv_data_185; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_375 = _GEN_8714 == 8'h2e ? _GEN_371 : phv_data_184; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_376 = mask_0[0] ? byte_ : phv_data_191; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_377 = mask_0[1] ? byte_1 : phv_data_190; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_378 = mask_0[2] ? byte_2 : phv_data_189; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_379 = mask_0[3] ? byte_3 : phv_data_188; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_380 = _GEN_8714 == 8'h2f ? _GEN_376 : phv_data_191; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_381 = _GEN_8714 == 8'h2f ? _GEN_377 : phv_data_190; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_382 = _GEN_8714 == 8'h2f ? _GEN_378 : phv_data_189; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_383 = _GEN_8714 == 8'h2f ? _GEN_379 : phv_data_188; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_384 = mask_0[0] ? byte_ : phv_data_195; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_385 = mask_0[1] ? byte_1 : phv_data_194; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_386 = mask_0[2] ? byte_2 : phv_data_193; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_387 = mask_0[3] ? byte_3 : phv_data_192; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_388 = _GEN_8714 == 8'h30 ? _GEN_384 : phv_data_195; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_389 = _GEN_8714 == 8'h30 ? _GEN_385 : phv_data_194; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_390 = _GEN_8714 == 8'h30 ? _GEN_386 : phv_data_193; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_391 = _GEN_8714 == 8'h30 ? _GEN_387 : phv_data_192; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_392 = mask_0[0] ? byte_ : phv_data_199; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_393 = mask_0[1] ? byte_1 : phv_data_198; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_394 = mask_0[2] ? byte_2 : phv_data_197; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_395 = mask_0[3] ? byte_3 : phv_data_196; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_396 = _GEN_8714 == 8'h31 ? _GEN_392 : phv_data_199; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_397 = _GEN_8714 == 8'h31 ? _GEN_393 : phv_data_198; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_398 = _GEN_8714 == 8'h31 ? _GEN_394 : phv_data_197; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_399 = _GEN_8714 == 8'h31 ? _GEN_395 : phv_data_196; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_400 = mask_0[0] ? byte_ : phv_data_203; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_401 = mask_0[1] ? byte_1 : phv_data_202; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_402 = mask_0[2] ? byte_2 : phv_data_201; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_403 = mask_0[3] ? byte_3 : phv_data_200; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_404 = _GEN_8714 == 8'h32 ? _GEN_400 : phv_data_203; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_405 = _GEN_8714 == 8'h32 ? _GEN_401 : phv_data_202; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_406 = _GEN_8714 == 8'h32 ? _GEN_402 : phv_data_201; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_407 = _GEN_8714 == 8'h32 ? _GEN_403 : phv_data_200; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_408 = mask_0[0] ? byte_ : phv_data_207; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_409 = mask_0[1] ? byte_1 : phv_data_206; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_410 = mask_0[2] ? byte_2 : phv_data_205; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_411 = mask_0[3] ? byte_3 : phv_data_204; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_412 = _GEN_8714 == 8'h33 ? _GEN_408 : phv_data_207; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_413 = _GEN_8714 == 8'h33 ? _GEN_409 : phv_data_206; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_414 = _GEN_8714 == 8'h33 ? _GEN_410 : phv_data_205; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_415 = _GEN_8714 == 8'h33 ? _GEN_411 : phv_data_204; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_416 = mask_0[0] ? byte_ : phv_data_211; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_417 = mask_0[1] ? byte_1 : phv_data_210; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_418 = mask_0[2] ? byte_2 : phv_data_209; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_419 = mask_0[3] ? byte_3 : phv_data_208; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_420 = _GEN_8714 == 8'h34 ? _GEN_416 : phv_data_211; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_421 = _GEN_8714 == 8'h34 ? _GEN_417 : phv_data_210; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_422 = _GEN_8714 == 8'h34 ? _GEN_418 : phv_data_209; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_423 = _GEN_8714 == 8'h34 ? _GEN_419 : phv_data_208; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_424 = mask_0[0] ? byte_ : phv_data_215; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_425 = mask_0[1] ? byte_1 : phv_data_214; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_426 = mask_0[2] ? byte_2 : phv_data_213; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_427 = mask_0[3] ? byte_3 : phv_data_212; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_428 = _GEN_8714 == 8'h35 ? _GEN_424 : phv_data_215; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_429 = _GEN_8714 == 8'h35 ? _GEN_425 : phv_data_214; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_430 = _GEN_8714 == 8'h35 ? _GEN_426 : phv_data_213; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_431 = _GEN_8714 == 8'h35 ? _GEN_427 : phv_data_212; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_432 = mask_0[0] ? byte_ : phv_data_219; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_433 = mask_0[1] ? byte_1 : phv_data_218; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_434 = mask_0[2] ? byte_2 : phv_data_217; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_435 = mask_0[3] ? byte_3 : phv_data_216; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_436 = _GEN_8714 == 8'h36 ? _GEN_432 : phv_data_219; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_437 = _GEN_8714 == 8'h36 ? _GEN_433 : phv_data_218; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_438 = _GEN_8714 == 8'h36 ? _GEN_434 : phv_data_217; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_439 = _GEN_8714 == 8'h36 ? _GEN_435 : phv_data_216; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_440 = mask_0[0] ? byte_ : phv_data_223; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_441 = mask_0[1] ? byte_1 : phv_data_222; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_442 = mask_0[2] ? byte_2 : phv_data_221; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_443 = mask_0[3] ? byte_3 : phv_data_220; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_444 = _GEN_8714 == 8'h37 ? _GEN_440 : phv_data_223; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_445 = _GEN_8714 == 8'h37 ? _GEN_441 : phv_data_222; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_446 = _GEN_8714 == 8'h37 ? _GEN_442 : phv_data_221; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_447 = _GEN_8714 == 8'h37 ? _GEN_443 : phv_data_220; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_448 = mask_0[0] ? byte_ : phv_data_227; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_449 = mask_0[1] ? byte_1 : phv_data_226; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_450 = mask_0[2] ? byte_2 : phv_data_225; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_451 = mask_0[3] ? byte_3 : phv_data_224; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_452 = _GEN_8714 == 8'h38 ? _GEN_448 : phv_data_227; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_453 = _GEN_8714 == 8'h38 ? _GEN_449 : phv_data_226; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_454 = _GEN_8714 == 8'h38 ? _GEN_450 : phv_data_225; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_455 = _GEN_8714 == 8'h38 ? _GEN_451 : phv_data_224; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_456 = mask_0[0] ? byte_ : phv_data_231; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_457 = mask_0[1] ? byte_1 : phv_data_230; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_458 = mask_0[2] ? byte_2 : phv_data_229; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_459 = mask_0[3] ? byte_3 : phv_data_228; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_460 = _GEN_8714 == 8'h39 ? _GEN_456 : phv_data_231; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_461 = _GEN_8714 == 8'h39 ? _GEN_457 : phv_data_230; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_462 = _GEN_8714 == 8'h39 ? _GEN_458 : phv_data_229; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_463 = _GEN_8714 == 8'h39 ? _GEN_459 : phv_data_228; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_464 = mask_0[0] ? byte_ : phv_data_235; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_465 = mask_0[1] ? byte_1 : phv_data_234; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_466 = mask_0[2] ? byte_2 : phv_data_233; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_467 = mask_0[3] ? byte_3 : phv_data_232; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_468 = _GEN_8714 == 8'h3a ? _GEN_464 : phv_data_235; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_469 = _GEN_8714 == 8'h3a ? _GEN_465 : phv_data_234; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_470 = _GEN_8714 == 8'h3a ? _GEN_466 : phv_data_233; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_471 = _GEN_8714 == 8'h3a ? _GEN_467 : phv_data_232; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_472 = mask_0[0] ? byte_ : phv_data_239; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_473 = mask_0[1] ? byte_1 : phv_data_238; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_474 = mask_0[2] ? byte_2 : phv_data_237; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_475 = mask_0[3] ? byte_3 : phv_data_236; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_476 = _GEN_8714 == 8'h3b ? _GEN_472 : phv_data_239; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_477 = _GEN_8714 == 8'h3b ? _GEN_473 : phv_data_238; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_478 = _GEN_8714 == 8'h3b ? _GEN_474 : phv_data_237; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_479 = _GEN_8714 == 8'h3b ? _GEN_475 : phv_data_236; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_480 = mask_0[0] ? byte_ : phv_data_243; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_481 = mask_0[1] ? byte_1 : phv_data_242; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_482 = mask_0[2] ? byte_2 : phv_data_241; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_483 = mask_0[3] ? byte_3 : phv_data_240; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_484 = _GEN_8714 == 8'h3c ? _GEN_480 : phv_data_243; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_485 = _GEN_8714 == 8'h3c ? _GEN_481 : phv_data_242; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_486 = _GEN_8714 == 8'h3c ? _GEN_482 : phv_data_241; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_487 = _GEN_8714 == 8'h3c ? _GEN_483 : phv_data_240; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_488 = mask_0[0] ? byte_ : phv_data_247; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_489 = mask_0[1] ? byte_1 : phv_data_246; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_490 = mask_0[2] ? byte_2 : phv_data_245; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_491 = mask_0[3] ? byte_3 : phv_data_244; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_492 = _GEN_8714 == 8'h3d ? _GEN_488 : phv_data_247; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_493 = _GEN_8714 == 8'h3d ? _GEN_489 : phv_data_246; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_494 = _GEN_8714 == 8'h3d ? _GEN_490 : phv_data_245; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_495 = _GEN_8714 == 8'h3d ? _GEN_491 : phv_data_244; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_496 = mask_0[0] ? byte_ : phv_data_251; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_497 = mask_0[1] ? byte_1 : phv_data_250; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_498 = mask_0[2] ? byte_2 : phv_data_249; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_499 = mask_0[3] ? byte_3 : phv_data_248; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_500 = _GEN_8714 == 8'h3e ? _GEN_496 : phv_data_251; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_501 = _GEN_8714 == 8'h3e ? _GEN_497 : phv_data_250; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_502 = _GEN_8714 == 8'h3e ? _GEN_498 : phv_data_249; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_503 = _GEN_8714 == 8'h3e ? _GEN_499 : phv_data_248; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_504 = mask_0[0] ? byte_ : phv_data_255; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_505 = mask_0[1] ? byte_1 : phv_data_254; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_506 = mask_0[2] ? byte_2 : phv_data_253; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_507 = mask_0[3] ? byte_3 : phv_data_252; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_508 = _GEN_8714 == 8'h3f ? _GEN_504 : phv_data_255; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_509 = _GEN_8714 == 8'h3f ? _GEN_505 : phv_data_254; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_510 = _GEN_8714 == 8'h3f ? _GEN_506 : phv_data_253; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_511 = _GEN_8714 == 8'h3f ? _GEN_507 : phv_data_252; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_512 = mask_0[0] ? byte_ : phv_data_259; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_513 = mask_0[1] ? byte_1 : phv_data_258; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_514 = mask_0[2] ? byte_2 : phv_data_257; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_515 = mask_0[3] ? byte_3 : phv_data_256; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_516 = _GEN_8714 == 8'h40 ? _GEN_512 : phv_data_259; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_517 = _GEN_8714 == 8'h40 ? _GEN_513 : phv_data_258; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_518 = _GEN_8714 == 8'h40 ? _GEN_514 : phv_data_257; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_519 = _GEN_8714 == 8'h40 ? _GEN_515 : phv_data_256; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_520 = mask_0[0] ? byte_ : phv_data_263; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_521 = mask_0[1] ? byte_1 : phv_data_262; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_522 = mask_0[2] ? byte_2 : phv_data_261; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_523 = mask_0[3] ? byte_3 : phv_data_260; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_524 = _GEN_8714 == 8'h41 ? _GEN_520 : phv_data_263; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_525 = _GEN_8714 == 8'h41 ? _GEN_521 : phv_data_262; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_526 = _GEN_8714 == 8'h41 ? _GEN_522 : phv_data_261; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_527 = _GEN_8714 == 8'h41 ? _GEN_523 : phv_data_260; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_528 = mask_0[0] ? byte_ : phv_data_267; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_529 = mask_0[1] ? byte_1 : phv_data_266; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_530 = mask_0[2] ? byte_2 : phv_data_265; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_531 = mask_0[3] ? byte_3 : phv_data_264; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_532 = _GEN_8714 == 8'h42 ? _GEN_528 : phv_data_267; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_533 = _GEN_8714 == 8'h42 ? _GEN_529 : phv_data_266; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_534 = _GEN_8714 == 8'h42 ? _GEN_530 : phv_data_265; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_535 = _GEN_8714 == 8'h42 ? _GEN_531 : phv_data_264; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_536 = mask_0[0] ? byte_ : phv_data_271; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_537 = mask_0[1] ? byte_1 : phv_data_270; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_538 = mask_0[2] ? byte_2 : phv_data_269; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_539 = mask_0[3] ? byte_3 : phv_data_268; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_540 = _GEN_8714 == 8'h43 ? _GEN_536 : phv_data_271; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_541 = _GEN_8714 == 8'h43 ? _GEN_537 : phv_data_270; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_542 = _GEN_8714 == 8'h43 ? _GEN_538 : phv_data_269; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_543 = _GEN_8714 == 8'h43 ? _GEN_539 : phv_data_268; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_544 = mask_0[0] ? byte_ : phv_data_275; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_545 = mask_0[1] ? byte_1 : phv_data_274; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_546 = mask_0[2] ? byte_2 : phv_data_273; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_547 = mask_0[3] ? byte_3 : phv_data_272; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_548 = _GEN_8714 == 8'h44 ? _GEN_544 : phv_data_275; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_549 = _GEN_8714 == 8'h44 ? _GEN_545 : phv_data_274; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_550 = _GEN_8714 == 8'h44 ? _GEN_546 : phv_data_273; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_551 = _GEN_8714 == 8'h44 ? _GEN_547 : phv_data_272; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_552 = mask_0[0] ? byte_ : phv_data_279; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_553 = mask_0[1] ? byte_1 : phv_data_278; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_554 = mask_0[2] ? byte_2 : phv_data_277; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_555 = mask_0[3] ? byte_3 : phv_data_276; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_556 = _GEN_8714 == 8'h45 ? _GEN_552 : phv_data_279; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_557 = _GEN_8714 == 8'h45 ? _GEN_553 : phv_data_278; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_558 = _GEN_8714 == 8'h45 ? _GEN_554 : phv_data_277; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_559 = _GEN_8714 == 8'h45 ? _GEN_555 : phv_data_276; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_560 = mask_0[0] ? byte_ : phv_data_283; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_561 = mask_0[1] ? byte_1 : phv_data_282; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_562 = mask_0[2] ? byte_2 : phv_data_281; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_563 = mask_0[3] ? byte_3 : phv_data_280; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_564 = _GEN_8714 == 8'h46 ? _GEN_560 : phv_data_283; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_565 = _GEN_8714 == 8'h46 ? _GEN_561 : phv_data_282; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_566 = _GEN_8714 == 8'h46 ? _GEN_562 : phv_data_281; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_567 = _GEN_8714 == 8'h46 ? _GEN_563 : phv_data_280; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_568 = mask_0[0] ? byte_ : phv_data_287; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_569 = mask_0[1] ? byte_1 : phv_data_286; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_570 = mask_0[2] ? byte_2 : phv_data_285; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_571 = mask_0[3] ? byte_3 : phv_data_284; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_572 = _GEN_8714 == 8'h47 ? _GEN_568 : phv_data_287; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_573 = _GEN_8714 == 8'h47 ? _GEN_569 : phv_data_286; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_574 = _GEN_8714 == 8'h47 ? _GEN_570 : phv_data_285; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_575 = _GEN_8714 == 8'h47 ? _GEN_571 : phv_data_284; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_576 = mask_0[0] ? byte_ : phv_data_291; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_577 = mask_0[1] ? byte_1 : phv_data_290; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_578 = mask_0[2] ? byte_2 : phv_data_289; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_579 = mask_0[3] ? byte_3 : phv_data_288; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_580 = _GEN_8714 == 8'h48 ? _GEN_576 : phv_data_291; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_581 = _GEN_8714 == 8'h48 ? _GEN_577 : phv_data_290; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_582 = _GEN_8714 == 8'h48 ? _GEN_578 : phv_data_289; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_583 = _GEN_8714 == 8'h48 ? _GEN_579 : phv_data_288; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_584 = mask_0[0] ? byte_ : phv_data_295; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_585 = mask_0[1] ? byte_1 : phv_data_294; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_586 = mask_0[2] ? byte_2 : phv_data_293; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_587 = mask_0[3] ? byte_3 : phv_data_292; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_588 = _GEN_8714 == 8'h49 ? _GEN_584 : phv_data_295; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_589 = _GEN_8714 == 8'h49 ? _GEN_585 : phv_data_294; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_590 = _GEN_8714 == 8'h49 ? _GEN_586 : phv_data_293; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_591 = _GEN_8714 == 8'h49 ? _GEN_587 : phv_data_292; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_592 = mask_0[0] ? byte_ : phv_data_299; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_593 = mask_0[1] ? byte_1 : phv_data_298; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_594 = mask_0[2] ? byte_2 : phv_data_297; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_595 = mask_0[3] ? byte_3 : phv_data_296; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_596 = _GEN_8714 == 8'h4a ? _GEN_592 : phv_data_299; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_597 = _GEN_8714 == 8'h4a ? _GEN_593 : phv_data_298; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_598 = _GEN_8714 == 8'h4a ? _GEN_594 : phv_data_297; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_599 = _GEN_8714 == 8'h4a ? _GEN_595 : phv_data_296; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_600 = mask_0[0] ? byte_ : phv_data_303; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_601 = mask_0[1] ? byte_1 : phv_data_302; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_602 = mask_0[2] ? byte_2 : phv_data_301; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_603 = mask_0[3] ? byte_3 : phv_data_300; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_604 = _GEN_8714 == 8'h4b ? _GEN_600 : phv_data_303; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_605 = _GEN_8714 == 8'h4b ? _GEN_601 : phv_data_302; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_606 = _GEN_8714 == 8'h4b ? _GEN_602 : phv_data_301; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_607 = _GEN_8714 == 8'h4b ? _GEN_603 : phv_data_300; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_608 = mask_0[0] ? byte_ : phv_data_307; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_609 = mask_0[1] ? byte_1 : phv_data_306; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_610 = mask_0[2] ? byte_2 : phv_data_305; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_611 = mask_0[3] ? byte_3 : phv_data_304; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_612 = _GEN_8714 == 8'h4c ? _GEN_608 : phv_data_307; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_613 = _GEN_8714 == 8'h4c ? _GEN_609 : phv_data_306; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_614 = _GEN_8714 == 8'h4c ? _GEN_610 : phv_data_305; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_615 = _GEN_8714 == 8'h4c ? _GEN_611 : phv_data_304; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_616 = mask_0[0] ? byte_ : phv_data_311; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_617 = mask_0[1] ? byte_1 : phv_data_310; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_618 = mask_0[2] ? byte_2 : phv_data_309; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_619 = mask_0[3] ? byte_3 : phv_data_308; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_620 = _GEN_8714 == 8'h4d ? _GEN_616 : phv_data_311; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_621 = _GEN_8714 == 8'h4d ? _GEN_617 : phv_data_310; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_622 = _GEN_8714 == 8'h4d ? _GEN_618 : phv_data_309; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_623 = _GEN_8714 == 8'h4d ? _GEN_619 : phv_data_308; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_624 = mask_0[0] ? byte_ : phv_data_315; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_625 = mask_0[1] ? byte_1 : phv_data_314; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_626 = mask_0[2] ? byte_2 : phv_data_313; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_627 = mask_0[3] ? byte_3 : phv_data_312; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_628 = _GEN_8714 == 8'h4e ? _GEN_624 : phv_data_315; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_629 = _GEN_8714 == 8'h4e ? _GEN_625 : phv_data_314; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_630 = _GEN_8714 == 8'h4e ? _GEN_626 : phv_data_313; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_631 = _GEN_8714 == 8'h4e ? _GEN_627 : phv_data_312; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_632 = mask_0[0] ? byte_ : phv_data_319; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_633 = mask_0[1] ? byte_1 : phv_data_318; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_634 = mask_0[2] ? byte_2 : phv_data_317; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_635 = mask_0[3] ? byte_3 : phv_data_316; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_636 = _GEN_8714 == 8'h4f ? _GEN_632 : phv_data_319; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_637 = _GEN_8714 == 8'h4f ? _GEN_633 : phv_data_318; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_638 = _GEN_8714 == 8'h4f ? _GEN_634 : phv_data_317; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_639 = _GEN_8714 == 8'h4f ? _GEN_635 : phv_data_316; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_640 = mask_0[0] ? byte_ : phv_data_323; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_641 = mask_0[1] ? byte_1 : phv_data_322; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_642 = mask_0[2] ? byte_2 : phv_data_321; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_643 = mask_0[3] ? byte_3 : phv_data_320; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_644 = _GEN_8714 == 8'h50 ? _GEN_640 : phv_data_323; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_645 = _GEN_8714 == 8'h50 ? _GEN_641 : phv_data_322; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_646 = _GEN_8714 == 8'h50 ? _GEN_642 : phv_data_321; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_647 = _GEN_8714 == 8'h50 ? _GEN_643 : phv_data_320; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_648 = mask_0[0] ? byte_ : phv_data_327; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_649 = mask_0[1] ? byte_1 : phv_data_326; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_650 = mask_0[2] ? byte_2 : phv_data_325; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_651 = mask_0[3] ? byte_3 : phv_data_324; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_652 = _GEN_8714 == 8'h51 ? _GEN_648 : phv_data_327; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_653 = _GEN_8714 == 8'h51 ? _GEN_649 : phv_data_326; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_654 = _GEN_8714 == 8'h51 ? _GEN_650 : phv_data_325; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_655 = _GEN_8714 == 8'h51 ? _GEN_651 : phv_data_324; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_656 = mask_0[0] ? byte_ : phv_data_331; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_657 = mask_0[1] ? byte_1 : phv_data_330; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_658 = mask_0[2] ? byte_2 : phv_data_329; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_659 = mask_0[3] ? byte_3 : phv_data_328; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_660 = _GEN_8714 == 8'h52 ? _GEN_656 : phv_data_331; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_661 = _GEN_8714 == 8'h52 ? _GEN_657 : phv_data_330; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_662 = _GEN_8714 == 8'h52 ? _GEN_658 : phv_data_329; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_663 = _GEN_8714 == 8'h52 ? _GEN_659 : phv_data_328; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_664 = mask_0[0] ? byte_ : phv_data_335; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_665 = mask_0[1] ? byte_1 : phv_data_334; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_666 = mask_0[2] ? byte_2 : phv_data_333; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_667 = mask_0[3] ? byte_3 : phv_data_332; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_668 = _GEN_8714 == 8'h53 ? _GEN_664 : phv_data_335; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_669 = _GEN_8714 == 8'h53 ? _GEN_665 : phv_data_334; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_670 = _GEN_8714 == 8'h53 ? _GEN_666 : phv_data_333; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_671 = _GEN_8714 == 8'h53 ? _GEN_667 : phv_data_332; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_672 = mask_0[0] ? byte_ : phv_data_339; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_673 = mask_0[1] ? byte_1 : phv_data_338; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_674 = mask_0[2] ? byte_2 : phv_data_337; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_675 = mask_0[3] ? byte_3 : phv_data_336; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_676 = _GEN_8714 == 8'h54 ? _GEN_672 : phv_data_339; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_677 = _GEN_8714 == 8'h54 ? _GEN_673 : phv_data_338; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_678 = _GEN_8714 == 8'h54 ? _GEN_674 : phv_data_337; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_679 = _GEN_8714 == 8'h54 ? _GEN_675 : phv_data_336; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_680 = mask_0[0] ? byte_ : phv_data_343; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_681 = mask_0[1] ? byte_1 : phv_data_342; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_682 = mask_0[2] ? byte_2 : phv_data_341; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_683 = mask_0[3] ? byte_3 : phv_data_340; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_684 = _GEN_8714 == 8'h55 ? _GEN_680 : phv_data_343; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_685 = _GEN_8714 == 8'h55 ? _GEN_681 : phv_data_342; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_686 = _GEN_8714 == 8'h55 ? _GEN_682 : phv_data_341; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_687 = _GEN_8714 == 8'h55 ? _GEN_683 : phv_data_340; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_688 = mask_0[0] ? byte_ : phv_data_347; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_689 = mask_0[1] ? byte_1 : phv_data_346; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_690 = mask_0[2] ? byte_2 : phv_data_345; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_691 = mask_0[3] ? byte_3 : phv_data_344; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_692 = _GEN_8714 == 8'h56 ? _GEN_688 : phv_data_347; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_693 = _GEN_8714 == 8'h56 ? _GEN_689 : phv_data_346; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_694 = _GEN_8714 == 8'h56 ? _GEN_690 : phv_data_345; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_695 = _GEN_8714 == 8'h56 ? _GEN_691 : phv_data_344; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_696 = mask_0[0] ? byte_ : phv_data_351; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_697 = mask_0[1] ? byte_1 : phv_data_350; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_698 = mask_0[2] ? byte_2 : phv_data_349; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_699 = mask_0[3] ? byte_3 : phv_data_348; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_700 = _GEN_8714 == 8'h57 ? _GEN_696 : phv_data_351; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_701 = _GEN_8714 == 8'h57 ? _GEN_697 : phv_data_350; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_702 = _GEN_8714 == 8'h57 ? _GEN_698 : phv_data_349; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_703 = _GEN_8714 == 8'h57 ? _GEN_699 : phv_data_348; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_704 = mask_0[0] ? byte_ : phv_data_355; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_705 = mask_0[1] ? byte_1 : phv_data_354; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_706 = mask_0[2] ? byte_2 : phv_data_353; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_707 = mask_0[3] ? byte_3 : phv_data_352; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_708 = _GEN_8714 == 8'h58 ? _GEN_704 : phv_data_355; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_709 = _GEN_8714 == 8'h58 ? _GEN_705 : phv_data_354; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_710 = _GEN_8714 == 8'h58 ? _GEN_706 : phv_data_353; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_711 = _GEN_8714 == 8'h58 ? _GEN_707 : phv_data_352; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_712 = mask_0[0] ? byte_ : phv_data_359; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_713 = mask_0[1] ? byte_1 : phv_data_358; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_714 = mask_0[2] ? byte_2 : phv_data_357; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_715 = mask_0[3] ? byte_3 : phv_data_356; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_716 = _GEN_8714 == 8'h59 ? _GEN_712 : phv_data_359; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_717 = _GEN_8714 == 8'h59 ? _GEN_713 : phv_data_358; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_718 = _GEN_8714 == 8'h59 ? _GEN_714 : phv_data_357; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_719 = _GEN_8714 == 8'h59 ? _GEN_715 : phv_data_356; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_720 = mask_0[0] ? byte_ : phv_data_363; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_721 = mask_0[1] ? byte_1 : phv_data_362; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_722 = mask_0[2] ? byte_2 : phv_data_361; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_723 = mask_0[3] ? byte_3 : phv_data_360; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_724 = _GEN_8714 == 8'h5a ? _GEN_720 : phv_data_363; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_725 = _GEN_8714 == 8'h5a ? _GEN_721 : phv_data_362; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_726 = _GEN_8714 == 8'h5a ? _GEN_722 : phv_data_361; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_727 = _GEN_8714 == 8'h5a ? _GEN_723 : phv_data_360; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_728 = mask_0[0] ? byte_ : phv_data_367; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_729 = mask_0[1] ? byte_1 : phv_data_366; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_730 = mask_0[2] ? byte_2 : phv_data_365; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_731 = mask_0[3] ? byte_3 : phv_data_364; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_732 = _GEN_8714 == 8'h5b ? _GEN_728 : phv_data_367; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_733 = _GEN_8714 == 8'h5b ? _GEN_729 : phv_data_366; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_734 = _GEN_8714 == 8'h5b ? _GEN_730 : phv_data_365; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_735 = _GEN_8714 == 8'h5b ? _GEN_731 : phv_data_364; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_736 = mask_0[0] ? byte_ : phv_data_371; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_737 = mask_0[1] ? byte_1 : phv_data_370; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_738 = mask_0[2] ? byte_2 : phv_data_369; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_739 = mask_0[3] ? byte_3 : phv_data_368; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_740 = _GEN_8714 == 8'h5c ? _GEN_736 : phv_data_371; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_741 = _GEN_8714 == 8'h5c ? _GEN_737 : phv_data_370; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_742 = _GEN_8714 == 8'h5c ? _GEN_738 : phv_data_369; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_743 = _GEN_8714 == 8'h5c ? _GEN_739 : phv_data_368; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_744 = mask_0[0] ? byte_ : phv_data_375; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_745 = mask_0[1] ? byte_1 : phv_data_374; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_746 = mask_0[2] ? byte_2 : phv_data_373; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_747 = mask_0[3] ? byte_3 : phv_data_372; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_748 = _GEN_8714 == 8'h5d ? _GEN_744 : phv_data_375; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_749 = _GEN_8714 == 8'h5d ? _GEN_745 : phv_data_374; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_750 = _GEN_8714 == 8'h5d ? _GEN_746 : phv_data_373; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_751 = _GEN_8714 == 8'h5d ? _GEN_747 : phv_data_372; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_752 = mask_0[0] ? byte_ : phv_data_379; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_753 = mask_0[1] ? byte_1 : phv_data_378; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_754 = mask_0[2] ? byte_2 : phv_data_377; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_755 = mask_0[3] ? byte_3 : phv_data_376; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_756 = _GEN_8714 == 8'h5e ? _GEN_752 : phv_data_379; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_757 = _GEN_8714 == 8'h5e ? _GEN_753 : phv_data_378; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_758 = _GEN_8714 == 8'h5e ? _GEN_754 : phv_data_377; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_759 = _GEN_8714 == 8'h5e ? _GEN_755 : phv_data_376; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_760 = mask_0[0] ? byte_ : phv_data_383; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_761 = mask_0[1] ? byte_1 : phv_data_382; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_762 = mask_0[2] ? byte_2 : phv_data_381; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_763 = mask_0[3] ? byte_3 : phv_data_380; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_764 = _GEN_8714 == 8'h5f ? _GEN_760 : phv_data_383; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_765 = _GEN_8714 == 8'h5f ? _GEN_761 : phv_data_382; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_766 = _GEN_8714 == 8'h5f ? _GEN_762 : phv_data_381; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_767 = _GEN_8714 == 8'h5f ? _GEN_763 : phv_data_380; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_768 = mask_0[0] ? byte_ : phv_data_387; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_769 = mask_0[1] ? byte_1 : phv_data_386; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_770 = mask_0[2] ? byte_2 : phv_data_385; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_771 = mask_0[3] ? byte_3 : phv_data_384; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_772 = _GEN_8714 == 8'h60 ? _GEN_768 : phv_data_387; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_773 = _GEN_8714 == 8'h60 ? _GEN_769 : phv_data_386; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_774 = _GEN_8714 == 8'h60 ? _GEN_770 : phv_data_385; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_775 = _GEN_8714 == 8'h60 ? _GEN_771 : phv_data_384; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_776 = mask_0[0] ? byte_ : phv_data_391; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_777 = mask_0[1] ? byte_1 : phv_data_390; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_778 = mask_0[2] ? byte_2 : phv_data_389; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_779 = mask_0[3] ? byte_3 : phv_data_388; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_780 = _GEN_8714 == 8'h61 ? _GEN_776 : phv_data_391; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_781 = _GEN_8714 == 8'h61 ? _GEN_777 : phv_data_390; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_782 = _GEN_8714 == 8'h61 ? _GEN_778 : phv_data_389; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_783 = _GEN_8714 == 8'h61 ? _GEN_779 : phv_data_388; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_784 = mask_0[0] ? byte_ : phv_data_395; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_785 = mask_0[1] ? byte_1 : phv_data_394; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_786 = mask_0[2] ? byte_2 : phv_data_393; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_787 = mask_0[3] ? byte_3 : phv_data_392; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_788 = _GEN_8714 == 8'h62 ? _GEN_784 : phv_data_395; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_789 = _GEN_8714 == 8'h62 ? _GEN_785 : phv_data_394; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_790 = _GEN_8714 == 8'h62 ? _GEN_786 : phv_data_393; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_791 = _GEN_8714 == 8'h62 ? _GEN_787 : phv_data_392; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_792 = mask_0[0] ? byte_ : phv_data_399; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_793 = mask_0[1] ? byte_1 : phv_data_398; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_794 = mask_0[2] ? byte_2 : phv_data_397; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_795 = mask_0[3] ? byte_3 : phv_data_396; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_796 = _GEN_8714 == 8'h63 ? _GEN_792 : phv_data_399; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_797 = _GEN_8714 == 8'h63 ? _GEN_793 : phv_data_398; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_798 = _GEN_8714 == 8'h63 ? _GEN_794 : phv_data_397; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_799 = _GEN_8714 == 8'h63 ? _GEN_795 : phv_data_396; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_800 = mask_0[0] ? byte_ : phv_data_403; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_801 = mask_0[1] ? byte_1 : phv_data_402; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_802 = mask_0[2] ? byte_2 : phv_data_401; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_803 = mask_0[3] ? byte_3 : phv_data_400; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_804 = _GEN_8714 == 8'h64 ? _GEN_800 : phv_data_403; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_805 = _GEN_8714 == 8'h64 ? _GEN_801 : phv_data_402; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_806 = _GEN_8714 == 8'h64 ? _GEN_802 : phv_data_401; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_807 = _GEN_8714 == 8'h64 ? _GEN_803 : phv_data_400; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_808 = mask_0[0] ? byte_ : phv_data_407; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_809 = mask_0[1] ? byte_1 : phv_data_406; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_810 = mask_0[2] ? byte_2 : phv_data_405; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_811 = mask_0[3] ? byte_3 : phv_data_404; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_812 = _GEN_8714 == 8'h65 ? _GEN_808 : phv_data_407; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_813 = _GEN_8714 == 8'h65 ? _GEN_809 : phv_data_406; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_814 = _GEN_8714 == 8'h65 ? _GEN_810 : phv_data_405; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_815 = _GEN_8714 == 8'h65 ? _GEN_811 : phv_data_404; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_816 = mask_0[0] ? byte_ : phv_data_411; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_817 = mask_0[1] ? byte_1 : phv_data_410; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_818 = mask_0[2] ? byte_2 : phv_data_409; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_819 = mask_0[3] ? byte_3 : phv_data_408; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_820 = _GEN_8714 == 8'h66 ? _GEN_816 : phv_data_411; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_821 = _GEN_8714 == 8'h66 ? _GEN_817 : phv_data_410; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_822 = _GEN_8714 == 8'h66 ? _GEN_818 : phv_data_409; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_823 = _GEN_8714 == 8'h66 ? _GEN_819 : phv_data_408; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_824 = mask_0[0] ? byte_ : phv_data_415; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_825 = mask_0[1] ? byte_1 : phv_data_414; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_826 = mask_0[2] ? byte_2 : phv_data_413; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_827 = mask_0[3] ? byte_3 : phv_data_412; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_828 = _GEN_8714 == 8'h67 ? _GEN_824 : phv_data_415; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_829 = _GEN_8714 == 8'h67 ? _GEN_825 : phv_data_414; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_830 = _GEN_8714 == 8'h67 ? _GEN_826 : phv_data_413; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_831 = _GEN_8714 == 8'h67 ? _GEN_827 : phv_data_412; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_832 = mask_0[0] ? byte_ : phv_data_419; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_833 = mask_0[1] ? byte_1 : phv_data_418; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_834 = mask_0[2] ? byte_2 : phv_data_417; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_835 = mask_0[3] ? byte_3 : phv_data_416; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_836 = _GEN_8714 == 8'h68 ? _GEN_832 : phv_data_419; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_837 = _GEN_8714 == 8'h68 ? _GEN_833 : phv_data_418; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_838 = _GEN_8714 == 8'h68 ? _GEN_834 : phv_data_417; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_839 = _GEN_8714 == 8'h68 ? _GEN_835 : phv_data_416; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_840 = mask_0[0] ? byte_ : phv_data_423; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_841 = mask_0[1] ? byte_1 : phv_data_422; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_842 = mask_0[2] ? byte_2 : phv_data_421; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_843 = mask_0[3] ? byte_3 : phv_data_420; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_844 = _GEN_8714 == 8'h69 ? _GEN_840 : phv_data_423; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_845 = _GEN_8714 == 8'h69 ? _GEN_841 : phv_data_422; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_846 = _GEN_8714 == 8'h69 ? _GEN_842 : phv_data_421; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_847 = _GEN_8714 == 8'h69 ? _GEN_843 : phv_data_420; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_848 = mask_0[0] ? byte_ : phv_data_427; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_849 = mask_0[1] ? byte_1 : phv_data_426; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_850 = mask_0[2] ? byte_2 : phv_data_425; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_851 = mask_0[3] ? byte_3 : phv_data_424; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_852 = _GEN_8714 == 8'h6a ? _GEN_848 : phv_data_427; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_853 = _GEN_8714 == 8'h6a ? _GEN_849 : phv_data_426; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_854 = _GEN_8714 == 8'h6a ? _GEN_850 : phv_data_425; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_855 = _GEN_8714 == 8'h6a ? _GEN_851 : phv_data_424; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_856 = mask_0[0] ? byte_ : phv_data_431; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_857 = mask_0[1] ? byte_1 : phv_data_430; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_858 = mask_0[2] ? byte_2 : phv_data_429; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_859 = mask_0[3] ? byte_3 : phv_data_428; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_860 = _GEN_8714 == 8'h6b ? _GEN_856 : phv_data_431; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_861 = _GEN_8714 == 8'h6b ? _GEN_857 : phv_data_430; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_862 = _GEN_8714 == 8'h6b ? _GEN_858 : phv_data_429; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_863 = _GEN_8714 == 8'h6b ? _GEN_859 : phv_data_428; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_864 = mask_0[0] ? byte_ : phv_data_435; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_865 = mask_0[1] ? byte_1 : phv_data_434; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_866 = mask_0[2] ? byte_2 : phv_data_433; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_867 = mask_0[3] ? byte_3 : phv_data_432; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_868 = _GEN_8714 == 8'h6c ? _GEN_864 : phv_data_435; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_869 = _GEN_8714 == 8'h6c ? _GEN_865 : phv_data_434; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_870 = _GEN_8714 == 8'h6c ? _GEN_866 : phv_data_433; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_871 = _GEN_8714 == 8'h6c ? _GEN_867 : phv_data_432; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_872 = mask_0[0] ? byte_ : phv_data_439; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_873 = mask_0[1] ? byte_1 : phv_data_438; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_874 = mask_0[2] ? byte_2 : phv_data_437; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_875 = mask_0[3] ? byte_3 : phv_data_436; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_876 = _GEN_8714 == 8'h6d ? _GEN_872 : phv_data_439; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_877 = _GEN_8714 == 8'h6d ? _GEN_873 : phv_data_438; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_878 = _GEN_8714 == 8'h6d ? _GEN_874 : phv_data_437; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_879 = _GEN_8714 == 8'h6d ? _GEN_875 : phv_data_436; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_880 = mask_0[0] ? byte_ : phv_data_443; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_881 = mask_0[1] ? byte_1 : phv_data_442; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_882 = mask_0[2] ? byte_2 : phv_data_441; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_883 = mask_0[3] ? byte_3 : phv_data_440; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_884 = _GEN_8714 == 8'h6e ? _GEN_880 : phv_data_443; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_885 = _GEN_8714 == 8'h6e ? _GEN_881 : phv_data_442; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_886 = _GEN_8714 == 8'h6e ? _GEN_882 : phv_data_441; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_887 = _GEN_8714 == 8'h6e ? _GEN_883 : phv_data_440; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_888 = mask_0[0] ? byte_ : phv_data_447; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_889 = mask_0[1] ? byte_1 : phv_data_446; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_890 = mask_0[2] ? byte_2 : phv_data_445; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_891 = mask_0[3] ? byte_3 : phv_data_444; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_892 = _GEN_8714 == 8'h6f ? _GEN_888 : phv_data_447; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_893 = _GEN_8714 == 8'h6f ? _GEN_889 : phv_data_446; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_894 = _GEN_8714 == 8'h6f ? _GEN_890 : phv_data_445; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_895 = _GEN_8714 == 8'h6f ? _GEN_891 : phv_data_444; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_896 = mask_0[0] ? byte_ : phv_data_451; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_897 = mask_0[1] ? byte_1 : phv_data_450; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_898 = mask_0[2] ? byte_2 : phv_data_449; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_899 = mask_0[3] ? byte_3 : phv_data_448; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_900 = _GEN_8714 == 8'h70 ? _GEN_896 : phv_data_451; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_901 = _GEN_8714 == 8'h70 ? _GEN_897 : phv_data_450; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_902 = _GEN_8714 == 8'h70 ? _GEN_898 : phv_data_449; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_903 = _GEN_8714 == 8'h70 ? _GEN_899 : phv_data_448; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_904 = mask_0[0] ? byte_ : phv_data_455; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_905 = mask_0[1] ? byte_1 : phv_data_454; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_906 = mask_0[2] ? byte_2 : phv_data_453; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_907 = mask_0[3] ? byte_3 : phv_data_452; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_908 = _GEN_8714 == 8'h71 ? _GEN_904 : phv_data_455; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_909 = _GEN_8714 == 8'h71 ? _GEN_905 : phv_data_454; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_910 = _GEN_8714 == 8'h71 ? _GEN_906 : phv_data_453; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_911 = _GEN_8714 == 8'h71 ? _GEN_907 : phv_data_452; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_912 = mask_0[0] ? byte_ : phv_data_459; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_913 = mask_0[1] ? byte_1 : phv_data_458; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_914 = mask_0[2] ? byte_2 : phv_data_457; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_915 = mask_0[3] ? byte_3 : phv_data_456; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_916 = _GEN_8714 == 8'h72 ? _GEN_912 : phv_data_459; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_917 = _GEN_8714 == 8'h72 ? _GEN_913 : phv_data_458; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_918 = _GEN_8714 == 8'h72 ? _GEN_914 : phv_data_457; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_919 = _GEN_8714 == 8'h72 ? _GEN_915 : phv_data_456; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_920 = mask_0[0] ? byte_ : phv_data_463; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_921 = mask_0[1] ? byte_1 : phv_data_462; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_922 = mask_0[2] ? byte_2 : phv_data_461; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_923 = mask_0[3] ? byte_3 : phv_data_460; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_924 = _GEN_8714 == 8'h73 ? _GEN_920 : phv_data_463; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_925 = _GEN_8714 == 8'h73 ? _GEN_921 : phv_data_462; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_926 = _GEN_8714 == 8'h73 ? _GEN_922 : phv_data_461; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_927 = _GEN_8714 == 8'h73 ? _GEN_923 : phv_data_460; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_928 = mask_0[0] ? byte_ : phv_data_467; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_929 = mask_0[1] ? byte_1 : phv_data_466; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_930 = mask_0[2] ? byte_2 : phv_data_465; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_931 = mask_0[3] ? byte_3 : phv_data_464; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_932 = _GEN_8714 == 8'h74 ? _GEN_928 : phv_data_467; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_933 = _GEN_8714 == 8'h74 ? _GEN_929 : phv_data_466; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_934 = _GEN_8714 == 8'h74 ? _GEN_930 : phv_data_465; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_935 = _GEN_8714 == 8'h74 ? _GEN_931 : phv_data_464; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_936 = mask_0[0] ? byte_ : phv_data_471; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_937 = mask_0[1] ? byte_1 : phv_data_470; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_938 = mask_0[2] ? byte_2 : phv_data_469; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_939 = mask_0[3] ? byte_3 : phv_data_468; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_940 = _GEN_8714 == 8'h75 ? _GEN_936 : phv_data_471; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_941 = _GEN_8714 == 8'h75 ? _GEN_937 : phv_data_470; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_942 = _GEN_8714 == 8'h75 ? _GEN_938 : phv_data_469; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_943 = _GEN_8714 == 8'h75 ? _GEN_939 : phv_data_468; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_944 = mask_0[0] ? byte_ : phv_data_475; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_945 = mask_0[1] ? byte_1 : phv_data_474; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_946 = mask_0[2] ? byte_2 : phv_data_473; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_947 = mask_0[3] ? byte_3 : phv_data_472; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_948 = _GEN_8714 == 8'h76 ? _GEN_944 : phv_data_475; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_949 = _GEN_8714 == 8'h76 ? _GEN_945 : phv_data_474; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_950 = _GEN_8714 == 8'h76 ? _GEN_946 : phv_data_473; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_951 = _GEN_8714 == 8'h76 ? _GEN_947 : phv_data_472; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_952 = mask_0[0] ? byte_ : phv_data_479; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_953 = mask_0[1] ? byte_1 : phv_data_478; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_954 = mask_0[2] ? byte_2 : phv_data_477; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_955 = mask_0[3] ? byte_3 : phv_data_476; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_956 = _GEN_8714 == 8'h77 ? _GEN_952 : phv_data_479; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_957 = _GEN_8714 == 8'h77 ? _GEN_953 : phv_data_478; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_958 = _GEN_8714 == 8'h77 ? _GEN_954 : phv_data_477; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_959 = _GEN_8714 == 8'h77 ? _GEN_955 : phv_data_476; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_960 = mask_0[0] ? byte_ : phv_data_483; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_961 = mask_0[1] ? byte_1 : phv_data_482; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_962 = mask_0[2] ? byte_2 : phv_data_481; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_963 = mask_0[3] ? byte_3 : phv_data_480; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_964 = _GEN_8714 == 8'h78 ? _GEN_960 : phv_data_483; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_965 = _GEN_8714 == 8'h78 ? _GEN_961 : phv_data_482; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_966 = _GEN_8714 == 8'h78 ? _GEN_962 : phv_data_481; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_967 = _GEN_8714 == 8'h78 ? _GEN_963 : phv_data_480; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_968 = mask_0[0] ? byte_ : phv_data_487; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_969 = mask_0[1] ? byte_1 : phv_data_486; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_970 = mask_0[2] ? byte_2 : phv_data_485; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_971 = mask_0[3] ? byte_3 : phv_data_484; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_972 = _GEN_8714 == 8'h79 ? _GEN_968 : phv_data_487; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_973 = _GEN_8714 == 8'h79 ? _GEN_969 : phv_data_486; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_974 = _GEN_8714 == 8'h79 ? _GEN_970 : phv_data_485; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_975 = _GEN_8714 == 8'h79 ? _GEN_971 : phv_data_484; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_976 = mask_0[0] ? byte_ : phv_data_491; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_977 = mask_0[1] ? byte_1 : phv_data_490; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_978 = mask_0[2] ? byte_2 : phv_data_489; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_979 = mask_0[3] ? byte_3 : phv_data_488; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_980 = _GEN_8714 == 8'h7a ? _GEN_976 : phv_data_491; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_981 = _GEN_8714 == 8'h7a ? _GEN_977 : phv_data_490; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_982 = _GEN_8714 == 8'h7a ? _GEN_978 : phv_data_489; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_983 = _GEN_8714 == 8'h7a ? _GEN_979 : phv_data_488; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_984 = mask_0[0] ? byte_ : phv_data_495; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_985 = mask_0[1] ? byte_1 : phv_data_494; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_986 = mask_0[2] ? byte_2 : phv_data_493; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_987 = mask_0[3] ? byte_3 : phv_data_492; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_988 = _GEN_8714 == 8'h7b ? _GEN_984 : phv_data_495; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_989 = _GEN_8714 == 8'h7b ? _GEN_985 : phv_data_494; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_990 = _GEN_8714 == 8'h7b ? _GEN_986 : phv_data_493; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_991 = _GEN_8714 == 8'h7b ? _GEN_987 : phv_data_492; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_992 = mask_0[0] ? byte_ : phv_data_499; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_993 = mask_0[1] ? byte_1 : phv_data_498; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_994 = mask_0[2] ? byte_2 : phv_data_497; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_995 = mask_0[3] ? byte_3 : phv_data_496; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_996 = _GEN_8714 == 8'h7c ? _GEN_992 : phv_data_499; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_997 = _GEN_8714 == 8'h7c ? _GEN_993 : phv_data_498; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_998 = _GEN_8714 == 8'h7c ? _GEN_994 : phv_data_497; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_999 = _GEN_8714 == 8'h7c ? _GEN_995 : phv_data_496; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1000 = mask_0[0] ? byte_ : phv_data_503; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1001 = mask_0[1] ? byte_1 : phv_data_502; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1002 = mask_0[2] ? byte_2 : phv_data_501; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1003 = mask_0[3] ? byte_3 : phv_data_500; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1004 = _GEN_8714 == 8'h7d ? _GEN_1000 : phv_data_503; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1005 = _GEN_8714 == 8'h7d ? _GEN_1001 : phv_data_502; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1006 = _GEN_8714 == 8'h7d ? _GEN_1002 : phv_data_501; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1007 = _GEN_8714 == 8'h7d ? _GEN_1003 : phv_data_500; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1008 = mask_0[0] ? byte_ : phv_data_507; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1009 = mask_0[1] ? byte_1 : phv_data_506; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1010 = mask_0[2] ? byte_2 : phv_data_505; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1011 = mask_0[3] ? byte_3 : phv_data_504; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1012 = _GEN_8714 == 8'h7e ? _GEN_1008 : phv_data_507; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1013 = _GEN_8714 == 8'h7e ? _GEN_1009 : phv_data_506; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1014 = _GEN_8714 == 8'h7e ? _GEN_1010 : phv_data_505; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1015 = _GEN_8714 == 8'h7e ? _GEN_1011 : phv_data_504; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1016 = mask_0[0] ? byte_ : phv_data_511; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1017 = mask_0[1] ? byte_1 : phv_data_510; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1018 = mask_0[2] ? byte_2 : phv_data_509; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1019 = mask_0[3] ? byte_3 : phv_data_508; // @[executor.scala 476:55 executor.scala 477:71 executor.scala 450:25]
  wire [7:0] _GEN_1020 = _GEN_8714 == 8'h7f ? _GEN_1016 : phv_data_511; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1021 = _GEN_8714 == 8'h7f ? _GEN_1017 : phv_data_510; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1022 = _GEN_8714 == 8'h7f ? _GEN_1018 : phv_data_509; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1023 = _GEN_8714 == 8'h7f ? _GEN_1019 : phv_data_508; // @[executor.scala 473:84 executor.scala 450:25]
  wire [7:0] _GEN_1024 = opcode != 4'h0 ? _GEN_4 : phv_data_3; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1025 = opcode != 4'h0 ? _GEN_5 : phv_data_2; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1026 = opcode != 4'h0 ? _GEN_6 : phv_data_1; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1027 = opcode != 4'h0 ? _GEN_7 : phv_data_0; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1028 = opcode != 4'h0 ? _GEN_12 : phv_data_7; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1029 = opcode != 4'h0 ? _GEN_13 : phv_data_6; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1030 = opcode != 4'h0 ? _GEN_14 : phv_data_5; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1031 = opcode != 4'h0 ? _GEN_15 : phv_data_4; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1032 = opcode != 4'h0 ? _GEN_20 : phv_data_11; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1033 = opcode != 4'h0 ? _GEN_21 : phv_data_10; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1034 = opcode != 4'h0 ? _GEN_22 : phv_data_9; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1035 = opcode != 4'h0 ? _GEN_23 : phv_data_8; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1036 = opcode != 4'h0 ? _GEN_28 : phv_data_15; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1037 = opcode != 4'h0 ? _GEN_29 : phv_data_14; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1038 = opcode != 4'h0 ? _GEN_30 : phv_data_13; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1039 = opcode != 4'h0 ? _GEN_31 : phv_data_12; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1040 = opcode != 4'h0 ? _GEN_36 : phv_data_19; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1041 = opcode != 4'h0 ? _GEN_37 : phv_data_18; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1042 = opcode != 4'h0 ? _GEN_38 : phv_data_17; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1043 = opcode != 4'h0 ? _GEN_39 : phv_data_16; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1044 = opcode != 4'h0 ? _GEN_44 : phv_data_23; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1045 = opcode != 4'h0 ? _GEN_45 : phv_data_22; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1046 = opcode != 4'h0 ? _GEN_46 : phv_data_21; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1047 = opcode != 4'h0 ? _GEN_47 : phv_data_20; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1048 = opcode != 4'h0 ? _GEN_52 : phv_data_27; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1049 = opcode != 4'h0 ? _GEN_53 : phv_data_26; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1050 = opcode != 4'h0 ? _GEN_54 : phv_data_25; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1051 = opcode != 4'h0 ? _GEN_55 : phv_data_24; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1052 = opcode != 4'h0 ? _GEN_60 : phv_data_31; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1053 = opcode != 4'h0 ? _GEN_61 : phv_data_30; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1054 = opcode != 4'h0 ? _GEN_62 : phv_data_29; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1055 = opcode != 4'h0 ? _GEN_63 : phv_data_28; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1056 = opcode != 4'h0 ? _GEN_68 : phv_data_35; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1057 = opcode != 4'h0 ? _GEN_69 : phv_data_34; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1058 = opcode != 4'h0 ? _GEN_70 : phv_data_33; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1059 = opcode != 4'h0 ? _GEN_71 : phv_data_32; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1060 = opcode != 4'h0 ? _GEN_76 : phv_data_39; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1061 = opcode != 4'h0 ? _GEN_77 : phv_data_38; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1062 = opcode != 4'h0 ? _GEN_78 : phv_data_37; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1063 = opcode != 4'h0 ? _GEN_79 : phv_data_36; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1064 = opcode != 4'h0 ? _GEN_84 : phv_data_43; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1065 = opcode != 4'h0 ? _GEN_85 : phv_data_42; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1066 = opcode != 4'h0 ? _GEN_86 : phv_data_41; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1067 = opcode != 4'h0 ? _GEN_87 : phv_data_40; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1068 = opcode != 4'h0 ? _GEN_92 : phv_data_47; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1069 = opcode != 4'h0 ? _GEN_93 : phv_data_46; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1070 = opcode != 4'h0 ? _GEN_94 : phv_data_45; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1071 = opcode != 4'h0 ? _GEN_95 : phv_data_44; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1072 = opcode != 4'h0 ? _GEN_100 : phv_data_51; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1073 = opcode != 4'h0 ? _GEN_101 : phv_data_50; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1074 = opcode != 4'h0 ? _GEN_102 : phv_data_49; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1075 = opcode != 4'h0 ? _GEN_103 : phv_data_48; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1076 = opcode != 4'h0 ? _GEN_108 : phv_data_55; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1077 = opcode != 4'h0 ? _GEN_109 : phv_data_54; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1078 = opcode != 4'h0 ? _GEN_110 : phv_data_53; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1079 = opcode != 4'h0 ? _GEN_111 : phv_data_52; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1080 = opcode != 4'h0 ? _GEN_116 : phv_data_59; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1081 = opcode != 4'h0 ? _GEN_117 : phv_data_58; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1082 = opcode != 4'h0 ? _GEN_118 : phv_data_57; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1083 = opcode != 4'h0 ? _GEN_119 : phv_data_56; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1084 = opcode != 4'h0 ? _GEN_124 : phv_data_63; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1085 = opcode != 4'h0 ? _GEN_125 : phv_data_62; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1086 = opcode != 4'h0 ? _GEN_126 : phv_data_61; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1087 = opcode != 4'h0 ? _GEN_127 : phv_data_60; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1088 = opcode != 4'h0 ? _GEN_132 : phv_data_67; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1089 = opcode != 4'h0 ? _GEN_133 : phv_data_66; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1090 = opcode != 4'h0 ? _GEN_134 : phv_data_65; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1091 = opcode != 4'h0 ? _GEN_135 : phv_data_64; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1092 = opcode != 4'h0 ? _GEN_140 : phv_data_71; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1093 = opcode != 4'h0 ? _GEN_141 : phv_data_70; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1094 = opcode != 4'h0 ? _GEN_142 : phv_data_69; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1095 = opcode != 4'h0 ? _GEN_143 : phv_data_68; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1096 = opcode != 4'h0 ? _GEN_148 : phv_data_75; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1097 = opcode != 4'h0 ? _GEN_149 : phv_data_74; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1098 = opcode != 4'h0 ? _GEN_150 : phv_data_73; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1099 = opcode != 4'h0 ? _GEN_151 : phv_data_72; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1100 = opcode != 4'h0 ? _GEN_156 : phv_data_79; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1101 = opcode != 4'h0 ? _GEN_157 : phv_data_78; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1102 = opcode != 4'h0 ? _GEN_158 : phv_data_77; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1103 = opcode != 4'h0 ? _GEN_159 : phv_data_76; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1104 = opcode != 4'h0 ? _GEN_164 : phv_data_83; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1105 = opcode != 4'h0 ? _GEN_165 : phv_data_82; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1106 = opcode != 4'h0 ? _GEN_166 : phv_data_81; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1107 = opcode != 4'h0 ? _GEN_167 : phv_data_80; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1108 = opcode != 4'h0 ? _GEN_172 : phv_data_87; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1109 = opcode != 4'h0 ? _GEN_173 : phv_data_86; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1110 = opcode != 4'h0 ? _GEN_174 : phv_data_85; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1111 = opcode != 4'h0 ? _GEN_175 : phv_data_84; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1112 = opcode != 4'h0 ? _GEN_180 : phv_data_91; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1113 = opcode != 4'h0 ? _GEN_181 : phv_data_90; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1114 = opcode != 4'h0 ? _GEN_182 : phv_data_89; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1115 = opcode != 4'h0 ? _GEN_183 : phv_data_88; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1116 = opcode != 4'h0 ? _GEN_188 : phv_data_95; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1117 = opcode != 4'h0 ? _GEN_189 : phv_data_94; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1118 = opcode != 4'h0 ? _GEN_190 : phv_data_93; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1119 = opcode != 4'h0 ? _GEN_191 : phv_data_92; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1120 = opcode != 4'h0 ? _GEN_196 : phv_data_99; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1121 = opcode != 4'h0 ? _GEN_197 : phv_data_98; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1122 = opcode != 4'h0 ? _GEN_198 : phv_data_97; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1123 = opcode != 4'h0 ? _GEN_199 : phv_data_96; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1124 = opcode != 4'h0 ? _GEN_204 : phv_data_103; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1125 = opcode != 4'h0 ? _GEN_205 : phv_data_102; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1126 = opcode != 4'h0 ? _GEN_206 : phv_data_101; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1127 = opcode != 4'h0 ? _GEN_207 : phv_data_100; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1128 = opcode != 4'h0 ? _GEN_212 : phv_data_107; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1129 = opcode != 4'h0 ? _GEN_213 : phv_data_106; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1130 = opcode != 4'h0 ? _GEN_214 : phv_data_105; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1131 = opcode != 4'h0 ? _GEN_215 : phv_data_104; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1132 = opcode != 4'h0 ? _GEN_220 : phv_data_111; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1133 = opcode != 4'h0 ? _GEN_221 : phv_data_110; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1134 = opcode != 4'h0 ? _GEN_222 : phv_data_109; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1135 = opcode != 4'h0 ? _GEN_223 : phv_data_108; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1136 = opcode != 4'h0 ? _GEN_228 : phv_data_115; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1137 = opcode != 4'h0 ? _GEN_229 : phv_data_114; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1138 = opcode != 4'h0 ? _GEN_230 : phv_data_113; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1139 = opcode != 4'h0 ? _GEN_231 : phv_data_112; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1140 = opcode != 4'h0 ? _GEN_236 : phv_data_119; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1141 = opcode != 4'h0 ? _GEN_237 : phv_data_118; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1142 = opcode != 4'h0 ? _GEN_238 : phv_data_117; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1143 = opcode != 4'h0 ? _GEN_239 : phv_data_116; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1144 = opcode != 4'h0 ? _GEN_244 : phv_data_123; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1145 = opcode != 4'h0 ? _GEN_245 : phv_data_122; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1146 = opcode != 4'h0 ? _GEN_246 : phv_data_121; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1147 = opcode != 4'h0 ? _GEN_247 : phv_data_120; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1148 = opcode != 4'h0 ? _GEN_252 : phv_data_127; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1149 = opcode != 4'h0 ? _GEN_253 : phv_data_126; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1150 = opcode != 4'h0 ? _GEN_254 : phv_data_125; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1151 = opcode != 4'h0 ? _GEN_255 : phv_data_124; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1152 = opcode != 4'h0 ? _GEN_260 : phv_data_131; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1153 = opcode != 4'h0 ? _GEN_261 : phv_data_130; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1154 = opcode != 4'h0 ? _GEN_262 : phv_data_129; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1155 = opcode != 4'h0 ? _GEN_263 : phv_data_128; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1156 = opcode != 4'h0 ? _GEN_268 : phv_data_135; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1157 = opcode != 4'h0 ? _GEN_269 : phv_data_134; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1158 = opcode != 4'h0 ? _GEN_270 : phv_data_133; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1159 = opcode != 4'h0 ? _GEN_271 : phv_data_132; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1160 = opcode != 4'h0 ? _GEN_276 : phv_data_139; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1161 = opcode != 4'h0 ? _GEN_277 : phv_data_138; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1162 = opcode != 4'h0 ? _GEN_278 : phv_data_137; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1163 = opcode != 4'h0 ? _GEN_279 : phv_data_136; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1164 = opcode != 4'h0 ? _GEN_284 : phv_data_143; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1165 = opcode != 4'h0 ? _GEN_285 : phv_data_142; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1166 = opcode != 4'h0 ? _GEN_286 : phv_data_141; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1167 = opcode != 4'h0 ? _GEN_287 : phv_data_140; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1168 = opcode != 4'h0 ? _GEN_292 : phv_data_147; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1169 = opcode != 4'h0 ? _GEN_293 : phv_data_146; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1170 = opcode != 4'h0 ? _GEN_294 : phv_data_145; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1171 = opcode != 4'h0 ? _GEN_295 : phv_data_144; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1172 = opcode != 4'h0 ? _GEN_300 : phv_data_151; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1173 = opcode != 4'h0 ? _GEN_301 : phv_data_150; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1174 = opcode != 4'h0 ? _GEN_302 : phv_data_149; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1175 = opcode != 4'h0 ? _GEN_303 : phv_data_148; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1176 = opcode != 4'h0 ? _GEN_308 : phv_data_155; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1177 = opcode != 4'h0 ? _GEN_309 : phv_data_154; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1178 = opcode != 4'h0 ? _GEN_310 : phv_data_153; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1179 = opcode != 4'h0 ? _GEN_311 : phv_data_152; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1180 = opcode != 4'h0 ? _GEN_316 : phv_data_159; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1181 = opcode != 4'h0 ? _GEN_317 : phv_data_158; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1182 = opcode != 4'h0 ? _GEN_318 : phv_data_157; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1183 = opcode != 4'h0 ? _GEN_319 : phv_data_156; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1184 = opcode != 4'h0 ? _GEN_324 : phv_data_163; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1185 = opcode != 4'h0 ? _GEN_325 : phv_data_162; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1186 = opcode != 4'h0 ? _GEN_326 : phv_data_161; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1187 = opcode != 4'h0 ? _GEN_327 : phv_data_160; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1188 = opcode != 4'h0 ? _GEN_332 : phv_data_167; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1189 = opcode != 4'h0 ? _GEN_333 : phv_data_166; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1190 = opcode != 4'h0 ? _GEN_334 : phv_data_165; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1191 = opcode != 4'h0 ? _GEN_335 : phv_data_164; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1192 = opcode != 4'h0 ? _GEN_340 : phv_data_171; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1193 = opcode != 4'h0 ? _GEN_341 : phv_data_170; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1194 = opcode != 4'h0 ? _GEN_342 : phv_data_169; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1195 = opcode != 4'h0 ? _GEN_343 : phv_data_168; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1196 = opcode != 4'h0 ? _GEN_348 : phv_data_175; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1197 = opcode != 4'h0 ? _GEN_349 : phv_data_174; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1198 = opcode != 4'h0 ? _GEN_350 : phv_data_173; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1199 = opcode != 4'h0 ? _GEN_351 : phv_data_172; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1200 = opcode != 4'h0 ? _GEN_356 : phv_data_179; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1201 = opcode != 4'h0 ? _GEN_357 : phv_data_178; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1202 = opcode != 4'h0 ? _GEN_358 : phv_data_177; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1203 = opcode != 4'h0 ? _GEN_359 : phv_data_176; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1204 = opcode != 4'h0 ? _GEN_364 : phv_data_183; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1205 = opcode != 4'h0 ? _GEN_365 : phv_data_182; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1206 = opcode != 4'h0 ? _GEN_366 : phv_data_181; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1207 = opcode != 4'h0 ? _GEN_367 : phv_data_180; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1208 = opcode != 4'h0 ? _GEN_372 : phv_data_187; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1209 = opcode != 4'h0 ? _GEN_373 : phv_data_186; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1210 = opcode != 4'h0 ? _GEN_374 : phv_data_185; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1211 = opcode != 4'h0 ? _GEN_375 : phv_data_184; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1212 = opcode != 4'h0 ? _GEN_380 : phv_data_191; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1213 = opcode != 4'h0 ? _GEN_381 : phv_data_190; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1214 = opcode != 4'h0 ? _GEN_382 : phv_data_189; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1215 = opcode != 4'h0 ? _GEN_383 : phv_data_188; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1216 = opcode != 4'h0 ? _GEN_388 : phv_data_195; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1217 = opcode != 4'h0 ? _GEN_389 : phv_data_194; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1218 = opcode != 4'h0 ? _GEN_390 : phv_data_193; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1219 = opcode != 4'h0 ? _GEN_391 : phv_data_192; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1220 = opcode != 4'h0 ? _GEN_396 : phv_data_199; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1221 = opcode != 4'h0 ? _GEN_397 : phv_data_198; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1222 = opcode != 4'h0 ? _GEN_398 : phv_data_197; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1223 = opcode != 4'h0 ? _GEN_399 : phv_data_196; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1224 = opcode != 4'h0 ? _GEN_404 : phv_data_203; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1225 = opcode != 4'h0 ? _GEN_405 : phv_data_202; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1226 = opcode != 4'h0 ? _GEN_406 : phv_data_201; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1227 = opcode != 4'h0 ? _GEN_407 : phv_data_200; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1228 = opcode != 4'h0 ? _GEN_412 : phv_data_207; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1229 = opcode != 4'h0 ? _GEN_413 : phv_data_206; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1230 = opcode != 4'h0 ? _GEN_414 : phv_data_205; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1231 = opcode != 4'h0 ? _GEN_415 : phv_data_204; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1232 = opcode != 4'h0 ? _GEN_420 : phv_data_211; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1233 = opcode != 4'h0 ? _GEN_421 : phv_data_210; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1234 = opcode != 4'h0 ? _GEN_422 : phv_data_209; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1235 = opcode != 4'h0 ? _GEN_423 : phv_data_208; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1236 = opcode != 4'h0 ? _GEN_428 : phv_data_215; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1237 = opcode != 4'h0 ? _GEN_429 : phv_data_214; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1238 = opcode != 4'h0 ? _GEN_430 : phv_data_213; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1239 = opcode != 4'h0 ? _GEN_431 : phv_data_212; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1240 = opcode != 4'h0 ? _GEN_436 : phv_data_219; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1241 = opcode != 4'h0 ? _GEN_437 : phv_data_218; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1242 = opcode != 4'h0 ? _GEN_438 : phv_data_217; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1243 = opcode != 4'h0 ? _GEN_439 : phv_data_216; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1244 = opcode != 4'h0 ? _GEN_444 : phv_data_223; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1245 = opcode != 4'h0 ? _GEN_445 : phv_data_222; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1246 = opcode != 4'h0 ? _GEN_446 : phv_data_221; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1247 = opcode != 4'h0 ? _GEN_447 : phv_data_220; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1248 = opcode != 4'h0 ? _GEN_452 : phv_data_227; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1249 = opcode != 4'h0 ? _GEN_453 : phv_data_226; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1250 = opcode != 4'h0 ? _GEN_454 : phv_data_225; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1251 = opcode != 4'h0 ? _GEN_455 : phv_data_224; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1252 = opcode != 4'h0 ? _GEN_460 : phv_data_231; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1253 = opcode != 4'h0 ? _GEN_461 : phv_data_230; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1254 = opcode != 4'h0 ? _GEN_462 : phv_data_229; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1255 = opcode != 4'h0 ? _GEN_463 : phv_data_228; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1256 = opcode != 4'h0 ? _GEN_468 : phv_data_235; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1257 = opcode != 4'h0 ? _GEN_469 : phv_data_234; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1258 = opcode != 4'h0 ? _GEN_470 : phv_data_233; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1259 = opcode != 4'h0 ? _GEN_471 : phv_data_232; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1260 = opcode != 4'h0 ? _GEN_476 : phv_data_239; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1261 = opcode != 4'h0 ? _GEN_477 : phv_data_238; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1262 = opcode != 4'h0 ? _GEN_478 : phv_data_237; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1263 = opcode != 4'h0 ? _GEN_479 : phv_data_236; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1264 = opcode != 4'h0 ? _GEN_484 : phv_data_243; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1265 = opcode != 4'h0 ? _GEN_485 : phv_data_242; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1266 = opcode != 4'h0 ? _GEN_486 : phv_data_241; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1267 = opcode != 4'h0 ? _GEN_487 : phv_data_240; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1268 = opcode != 4'h0 ? _GEN_492 : phv_data_247; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1269 = opcode != 4'h0 ? _GEN_493 : phv_data_246; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1270 = opcode != 4'h0 ? _GEN_494 : phv_data_245; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1271 = opcode != 4'h0 ? _GEN_495 : phv_data_244; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1272 = opcode != 4'h0 ? _GEN_500 : phv_data_251; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1273 = opcode != 4'h0 ? _GEN_501 : phv_data_250; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1274 = opcode != 4'h0 ? _GEN_502 : phv_data_249; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1275 = opcode != 4'h0 ? _GEN_503 : phv_data_248; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1276 = opcode != 4'h0 ? _GEN_508 : phv_data_255; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1277 = opcode != 4'h0 ? _GEN_509 : phv_data_254; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1278 = opcode != 4'h0 ? _GEN_510 : phv_data_253; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1279 = opcode != 4'h0 ? _GEN_511 : phv_data_252; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1280 = opcode != 4'h0 ? _GEN_516 : phv_data_259; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1281 = opcode != 4'h0 ? _GEN_517 : phv_data_258; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1282 = opcode != 4'h0 ? _GEN_518 : phv_data_257; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1283 = opcode != 4'h0 ? _GEN_519 : phv_data_256; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1284 = opcode != 4'h0 ? _GEN_524 : phv_data_263; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1285 = opcode != 4'h0 ? _GEN_525 : phv_data_262; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1286 = opcode != 4'h0 ? _GEN_526 : phv_data_261; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1287 = opcode != 4'h0 ? _GEN_527 : phv_data_260; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1288 = opcode != 4'h0 ? _GEN_532 : phv_data_267; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1289 = opcode != 4'h0 ? _GEN_533 : phv_data_266; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1290 = opcode != 4'h0 ? _GEN_534 : phv_data_265; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1291 = opcode != 4'h0 ? _GEN_535 : phv_data_264; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1292 = opcode != 4'h0 ? _GEN_540 : phv_data_271; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1293 = opcode != 4'h0 ? _GEN_541 : phv_data_270; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1294 = opcode != 4'h0 ? _GEN_542 : phv_data_269; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1295 = opcode != 4'h0 ? _GEN_543 : phv_data_268; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1296 = opcode != 4'h0 ? _GEN_548 : phv_data_275; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1297 = opcode != 4'h0 ? _GEN_549 : phv_data_274; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1298 = opcode != 4'h0 ? _GEN_550 : phv_data_273; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1299 = opcode != 4'h0 ? _GEN_551 : phv_data_272; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1300 = opcode != 4'h0 ? _GEN_556 : phv_data_279; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1301 = opcode != 4'h0 ? _GEN_557 : phv_data_278; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1302 = opcode != 4'h0 ? _GEN_558 : phv_data_277; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1303 = opcode != 4'h0 ? _GEN_559 : phv_data_276; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1304 = opcode != 4'h0 ? _GEN_564 : phv_data_283; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1305 = opcode != 4'h0 ? _GEN_565 : phv_data_282; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1306 = opcode != 4'h0 ? _GEN_566 : phv_data_281; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1307 = opcode != 4'h0 ? _GEN_567 : phv_data_280; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1308 = opcode != 4'h0 ? _GEN_572 : phv_data_287; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1309 = opcode != 4'h0 ? _GEN_573 : phv_data_286; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1310 = opcode != 4'h0 ? _GEN_574 : phv_data_285; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1311 = opcode != 4'h0 ? _GEN_575 : phv_data_284; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1312 = opcode != 4'h0 ? _GEN_580 : phv_data_291; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1313 = opcode != 4'h0 ? _GEN_581 : phv_data_290; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1314 = opcode != 4'h0 ? _GEN_582 : phv_data_289; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1315 = opcode != 4'h0 ? _GEN_583 : phv_data_288; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1316 = opcode != 4'h0 ? _GEN_588 : phv_data_295; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1317 = opcode != 4'h0 ? _GEN_589 : phv_data_294; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1318 = opcode != 4'h0 ? _GEN_590 : phv_data_293; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1319 = opcode != 4'h0 ? _GEN_591 : phv_data_292; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1320 = opcode != 4'h0 ? _GEN_596 : phv_data_299; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1321 = opcode != 4'h0 ? _GEN_597 : phv_data_298; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1322 = opcode != 4'h0 ? _GEN_598 : phv_data_297; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1323 = opcode != 4'h0 ? _GEN_599 : phv_data_296; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1324 = opcode != 4'h0 ? _GEN_604 : phv_data_303; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1325 = opcode != 4'h0 ? _GEN_605 : phv_data_302; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1326 = opcode != 4'h0 ? _GEN_606 : phv_data_301; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1327 = opcode != 4'h0 ? _GEN_607 : phv_data_300; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1328 = opcode != 4'h0 ? _GEN_612 : phv_data_307; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1329 = opcode != 4'h0 ? _GEN_613 : phv_data_306; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1330 = opcode != 4'h0 ? _GEN_614 : phv_data_305; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1331 = opcode != 4'h0 ? _GEN_615 : phv_data_304; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1332 = opcode != 4'h0 ? _GEN_620 : phv_data_311; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1333 = opcode != 4'h0 ? _GEN_621 : phv_data_310; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1334 = opcode != 4'h0 ? _GEN_622 : phv_data_309; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1335 = opcode != 4'h0 ? _GEN_623 : phv_data_308; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1336 = opcode != 4'h0 ? _GEN_628 : phv_data_315; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1337 = opcode != 4'h0 ? _GEN_629 : phv_data_314; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1338 = opcode != 4'h0 ? _GEN_630 : phv_data_313; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1339 = opcode != 4'h0 ? _GEN_631 : phv_data_312; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1340 = opcode != 4'h0 ? _GEN_636 : phv_data_319; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1341 = opcode != 4'h0 ? _GEN_637 : phv_data_318; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1342 = opcode != 4'h0 ? _GEN_638 : phv_data_317; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1343 = opcode != 4'h0 ? _GEN_639 : phv_data_316; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1344 = opcode != 4'h0 ? _GEN_644 : phv_data_323; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1345 = opcode != 4'h0 ? _GEN_645 : phv_data_322; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1346 = opcode != 4'h0 ? _GEN_646 : phv_data_321; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1347 = opcode != 4'h0 ? _GEN_647 : phv_data_320; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1348 = opcode != 4'h0 ? _GEN_652 : phv_data_327; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1349 = opcode != 4'h0 ? _GEN_653 : phv_data_326; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1350 = opcode != 4'h0 ? _GEN_654 : phv_data_325; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1351 = opcode != 4'h0 ? _GEN_655 : phv_data_324; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1352 = opcode != 4'h0 ? _GEN_660 : phv_data_331; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1353 = opcode != 4'h0 ? _GEN_661 : phv_data_330; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1354 = opcode != 4'h0 ? _GEN_662 : phv_data_329; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1355 = opcode != 4'h0 ? _GEN_663 : phv_data_328; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1356 = opcode != 4'h0 ? _GEN_668 : phv_data_335; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1357 = opcode != 4'h0 ? _GEN_669 : phv_data_334; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1358 = opcode != 4'h0 ? _GEN_670 : phv_data_333; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1359 = opcode != 4'h0 ? _GEN_671 : phv_data_332; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1360 = opcode != 4'h0 ? _GEN_676 : phv_data_339; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1361 = opcode != 4'h0 ? _GEN_677 : phv_data_338; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1362 = opcode != 4'h0 ? _GEN_678 : phv_data_337; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1363 = opcode != 4'h0 ? _GEN_679 : phv_data_336; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1364 = opcode != 4'h0 ? _GEN_684 : phv_data_343; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1365 = opcode != 4'h0 ? _GEN_685 : phv_data_342; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1366 = opcode != 4'h0 ? _GEN_686 : phv_data_341; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1367 = opcode != 4'h0 ? _GEN_687 : phv_data_340; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1368 = opcode != 4'h0 ? _GEN_692 : phv_data_347; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1369 = opcode != 4'h0 ? _GEN_693 : phv_data_346; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1370 = opcode != 4'h0 ? _GEN_694 : phv_data_345; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1371 = opcode != 4'h0 ? _GEN_695 : phv_data_344; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1372 = opcode != 4'h0 ? _GEN_700 : phv_data_351; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1373 = opcode != 4'h0 ? _GEN_701 : phv_data_350; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1374 = opcode != 4'h0 ? _GEN_702 : phv_data_349; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1375 = opcode != 4'h0 ? _GEN_703 : phv_data_348; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1376 = opcode != 4'h0 ? _GEN_708 : phv_data_355; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1377 = opcode != 4'h0 ? _GEN_709 : phv_data_354; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1378 = opcode != 4'h0 ? _GEN_710 : phv_data_353; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1379 = opcode != 4'h0 ? _GEN_711 : phv_data_352; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1380 = opcode != 4'h0 ? _GEN_716 : phv_data_359; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1381 = opcode != 4'h0 ? _GEN_717 : phv_data_358; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1382 = opcode != 4'h0 ? _GEN_718 : phv_data_357; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1383 = opcode != 4'h0 ? _GEN_719 : phv_data_356; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1384 = opcode != 4'h0 ? _GEN_724 : phv_data_363; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1385 = opcode != 4'h0 ? _GEN_725 : phv_data_362; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1386 = opcode != 4'h0 ? _GEN_726 : phv_data_361; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1387 = opcode != 4'h0 ? _GEN_727 : phv_data_360; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1388 = opcode != 4'h0 ? _GEN_732 : phv_data_367; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1389 = opcode != 4'h0 ? _GEN_733 : phv_data_366; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1390 = opcode != 4'h0 ? _GEN_734 : phv_data_365; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1391 = opcode != 4'h0 ? _GEN_735 : phv_data_364; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1392 = opcode != 4'h0 ? _GEN_740 : phv_data_371; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1393 = opcode != 4'h0 ? _GEN_741 : phv_data_370; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1394 = opcode != 4'h0 ? _GEN_742 : phv_data_369; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1395 = opcode != 4'h0 ? _GEN_743 : phv_data_368; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1396 = opcode != 4'h0 ? _GEN_748 : phv_data_375; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1397 = opcode != 4'h0 ? _GEN_749 : phv_data_374; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1398 = opcode != 4'h0 ? _GEN_750 : phv_data_373; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1399 = opcode != 4'h0 ? _GEN_751 : phv_data_372; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1400 = opcode != 4'h0 ? _GEN_756 : phv_data_379; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1401 = opcode != 4'h0 ? _GEN_757 : phv_data_378; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1402 = opcode != 4'h0 ? _GEN_758 : phv_data_377; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1403 = opcode != 4'h0 ? _GEN_759 : phv_data_376; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1404 = opcode != 4'h0 ? _GEN_764 : phv_data_383; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1405 = opcode != 4'h0 ? _GEN_765 : phv_data_382; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1406 = opcode != 4'h0 ? _GEN_766 : phv_data_381; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1407 = opcode != 4'h0 ? _GEN_767 : phv_data_380; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1408 = opcode != 4'h0 ? _GEN_772 : phv_data_387; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1409 = opcode != 4'h0 ? _GEN_773 : phv_data_386; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1410 = opcode != 4'h0 ? _GEN_774 : phv_data_385; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1411 = opcode != 4'h0 ? _GEN_775 : phv_data_384; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1412 = opcode != 4'h0 ? _GEN_780 : phv_data_391; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1413 = opcode != 4'h0 ? _GEN_781 : phv_data_390; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1414 = opcode != 4'h0 ? _GEN_782 : phv_data_389; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1415 = opcode != 4'h0 ? _GEN_783 : phv_data_388; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1416 = opcode != 4'h0 ? _GEN_788 : phv_data_395; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1417 = opcode != 4'h0 ? _GEN_789 : phv_data_394; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1418 = opcode != 4'h0 ? _GEN_790 : phv_data_393; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1419 = opcode != 4'h0 ? _GEN_791 : phv_data_392; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1420 = opcode != 4'h0 ? _GEN_796 : phv_data_399; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1421 = opcode != 4'h0 ? _GEN_797 : phv_data_398; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1422 = opcode != 4'h0 ? _GEN_798 : phv_data_397; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1423 = opcode != 4'h0 ? _GEN_799 : phv_data_396; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1424 = opcode != 4'h0 ? _GEN_804 : phv_data_403; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1425 = opcode != 4'h0 ? _GEN_805 : phv_data_402; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1426 = opcode != 4'h0 ? _GEN_806 : phv_data_401; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1427 = opcode != 4'h0 ? _GEN_807 : phv_data_400; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1428 = opcode != 4'h0 ? _GEN_812 : phv_data_407; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1429 = opcode != 4'h0 ? _GEN_813 : phv_data_406; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1430 = opcode != 4'h0 ? _GEN_814 : phv_data_405; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1431 = opcode != 4'h0 ? _GEN_815 : phv_data_404; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1432 = opcode != 4'h0 ? _GEN_820 : phv_data_411; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1433 = opcode != 4'h0 ? _GEN_821 : phv_data_410; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1434 = opcode != 4'h0 ? _GEN_822 : phv_data_409; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1435 = opcode != 4'h0 ? _GEN_823 : phv_data_408; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1436 = opcode != 4'h0 ? _GEN_828 : phv_data_415; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1437 = opcode != 4'h0 ? _GEN_829 : phv_data_414; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1438 = opcode != 4'h0 ? _GEN_830 : phv_data_413; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1439 = opcode != 4'h0 ? _GEN_831 : phv_data_412; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1440 = opcode != 4'h0 ? _GEN_836 : phv_data_419; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1441 = opcode != 4'h0 ? _GEN_837 : phv_data_418; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1442 = opcode != 4'h0 ? _GEN_838 : phv_data_417; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1443 = opcode != 4'h0 ? _GEN_839 : phv_data_416; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1444 = opcode != 4'h0 ? _GEN_844 : phv_data_423; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1445 = opcode != 4'h0 ? _GEN_845 : phv_data_422; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1446 = opcode != 4'h0 ? _GEN_846 : phv_data_421; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1447 = opcode != 4'h0 ? _GEN_847 : phv_data_420; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1448 = opcode != 4'h0 ? _GEN_852 : phv_data_427; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1449 = opcode != 4'h0 ? _GEN_853 : phv_data_426; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1450 = opcode != 4'h0 ? _GEN_854 : phv_data_425; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1451 = opcode != 4'h0 ? _GEN_855 : phv_data_424; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1452 = opcode != 4'h0 ? _GEN_860 : phv_data_431; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1453 = opcode != 4'h0 ? _GEN_861 : phv_data_430; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1454 = opcode != 4'h0 ? _GEN_862 : phv_data_429; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1455 = opcode != 4'h0 ? _GEN_863 : phv_data_428; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1456 = opcode != 4'h0 ? _GEN_868 : phv_data_435; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1457 = opcode != 4'h0 ? _GEN_869 : phv_data_434; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1458 = opcode != 4'h0 ? _GEN_870 : phv_data_433; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1459 = opcode != 4'h0 ? _GEN_871 : phv_data_432; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1460 = opcode != 4'h0 ? _GEN_876 : phv_data_439; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1461 = opcode != 4'h0 ? _GEN_877 : phv_data_438; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1462 = opcode != 4'h0 ? _GEN_878 : phv_data_437; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1463 = opcode != 4'h0 ? _GEN_879 : phv_data_436; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1464 = opcode != 4'h0 ? _GEN_884 : phv_data_443; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1465 = opcode != 4'h0 ? _GEN_885 : phv_data_442; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1466 = opcode != 4'h0 ? _GEN_886 : phv_data_441; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1467 = opcode != 4'h0 ? _GEN_887 : phv_data_440; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1468 = opcode != 4'h0 ? _GEN_892 : phv_data_447; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1469 = opcode != 4'h0 ? _GEN_893 : phv_data_446; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1470 = opcode != 4'h0 ? _GEN_894 : phv_data_445; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1471 = opcode != 4'h0 ? _GEN_895 : phv_data_444; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1472 = opcode != 4'h0 ? _GEN_900 : phv_data_451; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1473 = opcode != 4'h0 ? _GEN_901 : phv_data_450; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1474 = opcode != 4'h0 ? _GEN_902 : phv_data_449; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1475 = opcode != 4'h0 ? _GEN_903 : phv_data_448; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1476 = opcode != 4'h0 ? _GEN_908 : phv_data_455; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1477 = opcode != 4'h0 ? _GEN_909 : phv_data_454; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1478 = opcode != 4'h0 ? _GEN_910 : phv_data_453; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1479 = opcode != 4'h0 ? _GEN_911 : phv_data_452; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1480 = opcode != 4'h0 ? _GEN_916 : phv_data_459; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1481 = opcode != 4'h0 ? _GEN_917 : phv_data_458; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1482 = opcode != 4'h0 ? _GEN_918 : phv_data_457; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1483 = opcode != 4'h0 ? _GEN_919 : phv_data_456; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1484 = opcode != 4'h0 ? _GEN_924 : phv_data_463; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1485 = opcode != 4'h0 ? _GEN_925 : phv_data_462; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1486 = opcode != 4'h0 ? _GEN_926 : phv_data_461; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1487 = opcode != 4'h0 ? _GEN_927 : phv_data_460; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1488 = opcode != 4'h0 ? _GEN_932 : phv_data_467; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1489 = opcode != 4'h0 ? _GEN_933 : phv_data_466; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1490 = opcode != 4'h0 ? _GEN_934 : phv_data_465; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1491 = opcode != 4'h0 ? _GEN_935 : phv_data_464; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1492 = opcode != 4'h0 ? _GEN_940 : phv_data_471; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1493 = opcode != 4'h0 ? _GEN_941 : phv_data_470; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1494 = opcode != 4'h0 ? _GEN_942 : phv_data_469; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1495 = opcode != 4'h0 ? _GEN_943 : phv_data_468; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1496 = opcode != 4'h0 ? _GEN_948 : phv_data_475; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1497 = opcode != 4'h0 ? _GEN_949 : phv_data_474; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1498 = opcode != 4'h0 ? _GEN_950 : phv_data_473; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1499 = opcode != 4'h0 ? _GEN_951 : phv_data_472; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1500 = opcode != 4'h0 ? _GEN_956 : phv_data_479; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1501 = opcode != 4'h0 ? _GEN_957 : phv_data_478; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1502 = opcode != 4'h0 ? _GEN_958 : phv_data_477; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1503 = opcode != 4'h0 ? _GEN_959 : phv_data_476; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1504 = opcode != 4'h0 ? _GEN_964 : phv_data_483; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1505 = opcode != 4'h0 ? _GEN_965 : phv_data_482; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1506 = opcode != 4'h0 ? _GEN_966 : phv_data_481; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1507 = opcode != 4'h0 ? _GEN_967 : phv_data_480; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1508 = opcode != 4'h0 ? _GEN_972 : phv_data_487; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1509 = opcode != 4'h0 ? _GEN_973 : phv_data_486; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1510 = opcode != 4'h0 ? _GEN_974 : phv_data_485; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1511 = opcode != 4'h0 ? _GEN_975 : phv_data_484; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1512 = opcode != 4'h0 ? _GEN_980 : phv_data_491; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1513 = opcode != 4'h0 ? _GEN_981 : phv_data_490; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1514 = opcode != 4'h0 ? _GEN_982 : phv_data_489; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1515 = opcode != 4'h0 ? _GEN_983 : phv_data_488; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1516 = opcode != 4'h0 ? _GEN_988 : phv_data_495; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1517 = opcode != 4'h0 ? _GEN_989 : phv_data_494; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1518 = opcode != 4'h0 ? _GEN_990 : phv_data_493; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1519 = opcode != 4'h0 ? _GEN_991 : phv_data_492; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1520 = opcode != 4'h0 ? _GEN_996 : phv_data_499; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1521 = opcode != 4'h0 ? _GEN_997 : phv_data_498; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1522 = opcode != 4'h0 ? _GEN_998 : phv_data_497; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1523 = opcode != 4'h0 ? _GEN_999 : phv_data_496; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1524 = opcode != 4'h0 ? _GEN_1004 : phv_data_503; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1525 = opcode != 4'h0 ? _GEN_1005 : phv_data_502; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1526 = opcode != 4'h0 ? _GEN_1006 : phv_data_501; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1527 = opcode != 4'h0 ? _GEN_1007 : phv_data_500; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1528 = opcode != 4'h0 ? _GEN_1012 : phv_data_507; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1529 = opcode != 4'h0 ? _GEN_1013 : phv_data_506; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1530 = opcode != 4'h0 ? _GEN_1014 : phv_data_505; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1531 = opcode != 4'h0 ? _GEN_1015 : phv_data_504; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1532 = opcode != 4'h0 ? _GEN_1020 : phv_data_511; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1533 = opcode != 4'h0 ? _GEN_1021 : phv_data_510; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1534 = opcode != 4'h0 ? _GEN_1022 : phv_data_509; // @[executor.scala 470:55 executor.scala 450:25]
  wire [7:0] _GEN_1535 = opcode != 4'h0 ? _GEN_1023 : phv_data_508; // @[executor.scala 470:55 executor.scala 450:25]
  wire [3:0] _GEN_1536 = opcode == 4'hf ? parameter_2[13:10] : phv_next_processor_id; // @[executor.scala 466:52 executor.scala 467:55 executor.scala 450:25]
  wire  _GEN_1537 = opcode == 4'hf ? parameter_2[0] : phv_next_config_id; // @[executor.scala 466:52 executor.scala 468:55 executor.scala 450:25]
  wire [7:0] _GEN_1538 = opcode == 4'hf ? phv_data_3 : _GEN_1024; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1539 = opcode == 4'hf ? phv_data_2 : _GEN_1025; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1540 = opcode == 4'hf ? phv_data_1 : _GEN_1026; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1541 = opcode == 4'hf ? phv_data_0 : _GEN_1027; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1542 = opcode == 4'hf ? phv_data_7 : _GEN_1028; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1543 = opcode == 4'hf ? phv_data_6 : _GEN_1029; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1544 = opcode == 4'hf ? phv_data_5 : _GEN_1030; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1545 = opcode == 4'hf ? phv_data_4 : _GEN_1031; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1546 = opcode == 4'hf ? phv_data_11 : _GEN_1032; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1547 = opcode == 4'hf ? phv_data_10 : _GEN_1033; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1548 = opcode == 4'hf ? phv_data_9 : _GEN_1034; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1549 = opcode == 4'hf ? phv_data_8 : _GEN_1035; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1550 = opcode == 4'hf ? phv_data_15 : _GEN_1036; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1551 = opcode == 4'hf ? phv_data_14 : _GEN_1037; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1552 = opcode == 4'hf ? phv_data_13 : _GEN_1038; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1553 = opcode == 4'hf ? phv_data_12 : _GEN_1039; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1554 = opcode == 4'hf ? phv_data_19 : _GEN_1040; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1555 = opcode == 4'hf ? phv_data_18 : _GEN_1041; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1556 = opcode == 4'hf ? phv_data_17 : _GEN_1042; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1557 = opcode == 4'hf ? phv_data_16 : _GEN_1043; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1558 = opcode == 4'hf ? phv_data_23 : _GEN_1044; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1559 = opcode == 4'hf ? phv_data_22 : _GEN_1045; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1560 = opcode == 4'hf ? phv_data_21 : _GEN_1046; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1561 = opcode == 4'hf ? phv_data_20 : _GEN_1047; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1562 = opcode == 4'hf ? phv_data_27 : _GEN_1048; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1563 = opcode == 4'hf ? phv_data_26 : _GEN_1049; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1564 = opcode == 4'hf ? phv_data_25 : _GEN_1050; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1565 = opcode == 4'hf ? phv_data_24 : _GEN_1051; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1566 = opcode == 4'hf ? phv_data_31 : _GEN_1052; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1567 = opcode == 4'hf ? phv_data_30 : _GEN_1053; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1568 = opcode == 4'hf ? phv_data_29 : _GEN_1054; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1569 = opcode == 4'hf ? phv_data_28 : _GEN_1055; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1570 = opcode == 4'hf ? phv_data_35 : _GEN_1056; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1571 = opcode == 4'hf ? phv_data_34 : _GEN_1057; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1572 = opcode == 4'hf ? phv_data_33 : _GEN_1058; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1573 = opcode == 4'hf ? phv_data_32 : _GEN_1059; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1574 = opcode == 4'hf ? phv_data_39 : _GEN_1060; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1575 = opcode == 4'hf ? phv_data_38 : _GEN_1061; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1576 = opcode == 4'hf ? phv_data_37 : _GEN_1062; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1577 = opcode == 4'hf ? phv_data_36 : _GEN_1063; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1578 = opcode == 4'hf ? phv_data_43 : _GEN_1064; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1579 = opcode == 4'hf ? phv_data_42 : _GEN_1065; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1580 = opcode == 4'hf ? phv_data_41 : _GEN_1066; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1581 = opcode == 4'hf ? phv_data_40 : _GEN_1067; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1582 = opcode == 4'hf ? phv_data_47 : _GEN_1068; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1583 = opcode == 4'hf ? phv_data_46 : _GEN_1069; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1584 = opcode == 4'hf ? phv_data_45 : _GEN_1070; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1585 = opcode == 4'hf ? phv_data_44 : _GEN_1071; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1586 = opcode == 4'hf ? phv_data_51 : _GEN_1072; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1587 = opcode == 4'hf ? phv_data_50 : _GEN_1073; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1588 = opcode == 4'hf ? phv_data_49 : _GEN_1074; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1589 = opcode == 4'hf ? phv_data_48 : _GEN_1075; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1590 = opcode == 4'hf ? phv_data_55 : _GEN_1076; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1591 = opcode == 4'hf ? phv_data_54 : _GEN_1077; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1592 = opcode == 4'hf ? phv_data_53 : _GEN_1078; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1593 = opcode == 4'hf ? phv_data_52 : _GEN_1079; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1594 = opcode == 4'hf ? phv_data_59 : _GEN_1080; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1595 = opcode == 4'hf ? phv_data_58 : _GEN_1081; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1596 = opcode == 4'hf ? phv_data_57 : _GEN_1082; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1597 = opcode == 4'hf ? phv_data_56 : _GEN_1083; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1598 = opcode == 4'hf ? phv_data_63 : _GEN_1084; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1599 = opcode == 4'hf ? phv_data_62 : _GEN_1085; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1600 = opcode == 4'hf ? phv_data_61 : _GEN_1086; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1601 = opcode == 4'hf ? phv_data_60 : _GEN_1087; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1602 = opcode == 4'hf ? phv_data_67 : _GEN_1088; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1603 = opcode == 4'hf ? phv_data_66 : _GEN_1089; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1604 = opcode == 4'hf ? phv_data_65 : _GEN_1090; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1605 = opcode == 4'hf ? phv_data_64 : _GEN_1091; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1606 = opcode == 4'hf ? phv_data_71 : _GEN_1092; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1607 = opcode == 4'hf ? phv_data_70 : _GEN_1093; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1608 = opcode == 4'hf ? phv_data_69 : _GEN_1094; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1609 = opcode == 4'hf ? phv_data_68 : _GEN_1095; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1610 = opcode == 4'hf ? phv_data_75 : _GEN_1096; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1611 = opcode == 4'hf ? phv_data_74 : _GEN_1097; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1612 = opcode == 4'hf ? phv_data_73 : _GEN_1098; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1613 = opcode == 4'hf ? phv_data_72 : _GEN_1099; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1614 = opcode == 4'hf ? phv_data_79 : _GEN_1100; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1615 = opcode == 4'hf ? phv_data_78 : _GEN_1101; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1616 = opcode == 4'hf ? phv_data_77 : _GEN_1102; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1617 = opcode == 4'hf ? phv_data_76 : _GEN_1103; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1618 = opcode == 4'hf ? phv_data_83 : _GEN_1104; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1619 = opcode == 4'hf ? phv_data_82 : _GEN_1105; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1620 = opcode == 4'hf ? phv_data_81 : _GEN_1106; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1621 = opcode == 4'hf ? phv_data_80 : _GEN_1107; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1622 = opcode == 4'hf ? phv_data_87 : _GEN_1108; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1623 = opcode == 4'hf ? phv_data_86 : _GEN_1109; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1624 = opcode == 4'hf ? phv_data_85 : _GEN_1110; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1625 = opcode == 4'hf ? phv_data_84 : _GEN_1111; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1626 = opcode == 4'hf ? phv_data_91 : _GEN_1112; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1627 = opcode == 4'hf ? phv_data_90 : _GEN_1113; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1628 = opcode == 4'hf ? phv_data_89 : _GEN_1114; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1629 = opcode == 4'hf ? phv_data_88 : _GEN_1115; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1630 = opcode == 4'hf ? phv_data_95 : _GEN_1116; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1631 = opcode == 4'hf ? phv_data_94 : _GEN_1117; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1632 = opcode == 4'hf ? phv_data_93 : _GEN_1118; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1633 = opcode == 4'hf ? phv_data_92 : _GEN_1119; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1634 = opcode == 4'hf ? phv_data_99 : _GEN_1120; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1635 = opcode == 4'hf ? phv_data_98 : _GEN_1121; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1636 = opcode == 4'hf ? phv_data_97 : _GEN_1122; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1637 = opcode == 4'hf ? phv_data_96 : _GEN_1123; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1638 = opcode == 4'hf ? phv_data_103 : _GEN_1124; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1639 = opcode == 4'hf ? phv_data_102 : _GEN_1125; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1640 = opcode == 4'hf ? phv_data_101 : _GEN_1126; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1641 = opcode == 4'hf ? phv_data_100 : _GEN_1127; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1642 = opcode == 4'hf ? phv_data_107 : _GEN_1128; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1643 = opcode == 4'hf ? phv_data_106 : _GEN_1129; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1644 = opcode == 4'hf ? phv_data_105 : _GEN_1130; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1645 = opcode == 4'hf ? phv_data_104 : _GEN_1131; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1646 = opcode == 4'hf ? phv_data_111 : _GEN_1132; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1647 = opcode == 4'hf ? phv_data_110 : _GEN_1133; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1648 = opcode == 4'hf ? phv_data_109 : _GEN_1134; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1649 = opcode == 4'hf ? phv_data_108 : _GEN_1135; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1650 = opcode == 4'hf ? phv_data_115 : _GEN_1136; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1651 = opcode == 4'hf ? phv_data_114 : _GEN_1137; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1652 = opcode == 4'hf ? phv_data_113 : _GEN_1138; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1653 = opcode == 4'hf ? phv_data_112 : _GEN_1139; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1654 = opcode == 4'hf ? phv_data_119 : _GEN_1140; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1655 = opcode == 4'hf ? phv_data_118 : _GEN_1141; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1656 = opcode == 4'hf ? phv_data_117 : _GEN_1142; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1657 = opcode == 4'hf ? phv_data_116 : _GEN_1143; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1658 = opcode == 4'hf ? phv_data_123 : _GEN_1144; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1659 = opcode == 4'hf ? phv_data_122 : _GEN_1145; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1660 = opcode == 4'hf ? phv_data_121 : _GEN_1146; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1661 = opcode == 4'hf ? phv_data_120 : _GEN_1147; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1662 = opcode == 4'hf ? phv_data_127 : _GEN_1148; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1663 = opcode == 4'hf ? phv_data_126 : _GEN_1149; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1664 = opcode == 4'hf ? phv_data_125 : _GEN_1150; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1665 = opcode == 4'hf ? phv_data_124 : _GEN_1151; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1666 = opcode == 4'hf ? phv_data_131 : _GEN_1152; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1667 = opcode == 4'hf ? phv_data_130 : _GEN_1153; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1668 = opcode == 4'hf ? phv_data_129 : _GEN_1154; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1669 = opcode == 4'hf ? phv_data_128 : _GEN_1155; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1670 = opcode == 4'hf ? phv_data_135 : _GEN_1156; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1671 = opcode == 4'hf ? phv_data_134 : _GEN_1157; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1672 = opcode == 4'hf ? phv_data_133 : _GEN_1158; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1673 = opcode == 4'hf ? phv_data_132 : _GEN_1159; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1674 = opcode == 4'hf ? phv_data_139 : _GEN_1160; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1675 = opcode == 4'hf ? phv_data_138 : _GEN_1161; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1676 = opcode == 4'hf ? phv_data_137 : _GEN_1162; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1677 = opcode == 4'hf ? phv_data_136 : _GEN_1163; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1678 = opcode == 4'hf ? phv_data_143 : _GEN_1164; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1679 = opcode == 4'hf ? phv_data_142 : _GEN_1165; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1680 = opcode == 4'hf ? phv_data_141 : _GEN_1166; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1681 = opcode == 4'hf ? phv_data_140 : _GEN_1167; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1682 = opcode == 4'hf ? phv_data_147 : _GEN_1168; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1683 = opcode == 4'hf ? phv_data_146 : _GEN_1169; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1684 = opcode == 4'hf ? phv_data_145 : _GEN_1170; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1685 = opcode == 4'hf ? phv_data_144 : _GEN_1171; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1686 = opcode == 4'hf ? phv_data_151 : _GEN_1172; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1687 = opcode == 4'hf ? phv_data_150 : _GEN_1173; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1688 = opcode == 4'hf ? phv_data_149 : _GEN_1174; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1689 = opcode == 4'hf ? phv_data_148 : _GEN_1175; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1690 = opcode == 4'hf ? phv_data_155 : _GEN_1176; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1691 = opcode == 4'hf ? phv_data_154 : _GEN_1177; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1692 = opcode == 4'hf ? phv_data_153 : _GEN_1178; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1693 = opcode == 4'hf ? phv_data_152 : _GEN_1179; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1694 = opcode == 4'hf ? phv_data_159 : _GEN_1180; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1695 = opcode == 4'hf ? phv_data_158 : _GEN_1181; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1696 = opcode == 4'hf ? phv_data_157 : _GEN_1182; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1697 = opcode == 4'hf ? phv_data_156 : _GEN_1183; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1698 = opcode == 4'hf ? phv_data_163 : _GEN_1184; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1699 = opcode == 4'hf ? phv_data_162 : _GEN_1185; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1700 = opcode == 4'hf ? phv_data_161 : _GEN_1186; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1701 = opcode == 4'hf ? phv_data_160 : _GEN_1187; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1702 = opcode == 4'hf ? phv_data_167 : _GEN_1188; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1703 = opcode == 4'hf ? phv_data_166 : _GEN_1189; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1704 = opcode == 4'hf ? phv_data_165 : _GEN_1190; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1705 = opcode == 4'hf ? phv_data_164 : _GEN_1191; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1706 = opcode == 4'hf ? phv_data_171 : _GEN_1192; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1707 = opcode == 4'hf ? phv_data_170 : _GEN_1193; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1708 = opcode == 4'hf ? phv_data_169 : _GEN_1194; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1709 = opcode == 4'hf ? phv_data_168 : _GEN_1195; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1710 = opcode == 4'hf ? phv_data_175 : _GEN_1196; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1711 = opcode == 4'hf ? phv_data_174 : _GEN_1197; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1712 = opcode == 4'hf ? phv_data_173 : _GEN_1198; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1713 = opcode == 4'hf ? phv_data_172 : _GEN_1199; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1714 = opcode == 4'hf ? phv_data_179 : _GEN_1200; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1715 = opcode == 4'hf ? phv_data_178 : _GEN_1201; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1716 = opcode == 4'hf ? phv_data_177 : _GEN_1202; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1717 = opcode == 4'hf ? phv_data_176 : _GEN_1203; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1718 = opcode == 4'hf ? phv_data_183 : _GEN_1204; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1719 = opcode == 4'hf ? phv_data_182 : _GEN_1205; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1720 = opcode == 4'hf ? phv_data_181 : _GEN_1206; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1721 = opcode == 4'hf ? phv_data_180 : _GEN_1207; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1722 = opcode == 4'hf ? phv_data_187 : _GEN_1208; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1723 = opcode == 4'hf ? phv_data_186 : _GEN_1209; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1724 = opcode == 4'hf ? phv_data_185 : _GEN_1210; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1725 = opcode == 4'hf ? phv_data_184 : _GEN_1211; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1726 = opcode == 4'hf ? phv_data_191 : _GEN_1212; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1727 = opcode == 4'hf ? phv_data_190 : _GEN_1213; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1728 = opcode == 4'hf ? phv_data_189 : _GEN_1214; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1729 = opcode == 4'hf ? phv_data_188 : _GEN_1215; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1730 = opcode == 4'hf ? phv_data_195 : _GEN_1216; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1731 = opcode == 4'hf ? phv_data_194 : _GEN_1217; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1732 = opcode == 4'hf ? phv_data_193 : _GEN_1218; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1733 = opcode == 4'hf ? phv_data_192 : _GEN_1219; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1734 = opcode == 4'hf ? phv_data_199 : _GEN_1220; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1735 = opcode == 4'hf ? phv_data_198 : _GEN_1221; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1736 = opcode == 4'hf ? phv_data_197 : _GEN_1222; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1737 = opcode == 4'hf ? phv_data_196 : _GEN_1223; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1738 = opcode == 4'hf ? phv_data_203 : _GEN_1224; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1739 = opcode == 4'hf ? phv_data_202 : _GEN_1225; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1740 = opcode == 4'hf ? phv_data_201 : _GEN_1226; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1741 = opcode == 4'hf ? phv_data_200 : _GEN_1227; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1742 = opcode == 4'hf ? phv_data_207 : _GEN_1228; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1743 = opcode == 4'hf ? phv_data_206 : _GEN_1229; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1744 = opcode == 4'hf ? phv_data_205 : _GEN_1230; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1745 = opcode == 4'hf ? phv_data_204 : _GEN_1231; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1746 = opcode == 4'hf ? phv_data_211 : _GEN_1232; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1747 = opcode == 4'hf ? phv_data_210 : _GEN_1233; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1748 = opcode == 4'hf ? phv_data_209 : _GEN_1234; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1749 = opcode == 4'hf ? phv_data_208 : _GEN_1235; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1750 = opcode == 4'hf ? phv_data_215 : _GEN_1236; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1751 = opcode == 4'hf ? phv_data_214 : _GEN_1237; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1752 = opcode == 4'hf ? phv_data_213 : _GEN_1238; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1753 = opcode == 4'hf ? phv_data_212 : _GEN_1239; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1754 = opcode == 4'hf ? phv_data_219 : _GEN_1240; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1755 = opcode == 4'hf ? phv_data_218 : _GEN_1241; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1756 = opcode == 4'hf ? phv_data_217 : _GEN_1242; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1757 = opcode == 4'hf ? phv_data_216 : _GEN_1243; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1758 = opcode == 4'hf ? phv_data_223 : _GEN_1244; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1759 = opcode == 4'hf ? phv_data_222 : _GEN_1245; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1760 = opcode == 4'hf ? phv_data_221 : _GEN_1246; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1761 = opcode == 4'hf ? phv_data_220 : _GEN_1247; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1762 = opcode == 4'hf ? phv_data_227 : _GEN_1248; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1763 = opcode == 4'hf ? phv_data_226 : _GEN_1249; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1764 = opcode == 4'hf ? phv_data_225 : _GEN_1250; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1765 = opcode == 4'hf ? phv_data_224 : _GEN_1251; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1766 = opcode == 4'hf ? phv_data_231 : _GEN_1252; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1767 = opcode == 4'hf ? phv_data_230 : _GEN_1253; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1768 = opcode == 4'hf ? phv_data_229 : _GEN_1254; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1769 = opcode == 4'hf ? phv_data_228 : _GEN_1255; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1770 = opcode == 4'hf ? phv_data_235 : _GEN_1256; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1771 = opcode == 4'hf ? phv_data_234 : _GEN_1257; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1772 = opcode == 4'hf ? phv_data_233 : _GEN_1258; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1773 = opcode == 4'hf ? phv_data_232 : _GEN_1259; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1774 = opcode == 4'hf ? phv_data_239 : _GEN_1260; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1775 = opcode == 4'hf ? phv_data_238 : _GEN_1261; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1776 = opcode == 4'hf ? phv_data_237 : _GEN_1262; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1777 = opcode == 4'hf ? phv_data_236 : _GEN_1263; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1778 = opcode == 4'hf ? phv_data_243 : _GEN_1264; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1779 = opcode == 4'hf ? phv_data_242 : _GEN_1265; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1780 = opcode == 4'hf ? phv_data_241 : _GEN_1266; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1781 = opcode == 4'hf ? phv_data_240 : _GEN_1267; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1782 = opcode == 4'hf ? phv_data_247 : _GEN_1268; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1783 = opcode == 4'hf ? phv_data_246 : _GEN_1269; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1784 = opcode == 4'hf ? phv_data_245 : _GEN_1270; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1785 = opcode == 4'hf ? phv_data_244 : _GEN_1271; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1786 = opcode == 4'hf ? phv_data_251 : _GEN_1272; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1787 = opcode == 4'hf ? phv_data_250 : _GEN_1273; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1788 = opcode == 4'hf ? phv_data_249 : _GEN_1274; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1789 = opcode == 4'hf ? phv_data_248 : _GEN_1275; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1790 = opcode == 4'hf ? phv_data_255 : _GEN_1276; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1791 = opcode == 4'hf ? phv_data_254 : _GEN_1277; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1792 = opcode == 4'hf ? phv_data_253 : _GEN_1278; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1793 = opcode == 4'hf ? phv_data_252 : _GEN_1279; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1794 = opcode == 4'hf ? phv_data_259 : _GEN_1280; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1795 = opcode == 4'hf ? phv_data_258 : _GEN_1281; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1796 = opcode == 4'hf ? phv_data_257 : _GEN_1282; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1797 = opcode == 4'hf ? phv_data_256 : _GEN_1283; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1798 = opcode == 4'hf ? phv_data_263 : _GEN_1284; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1799 = opcode == 4'hf ? phv_data_262 : _GEN_1285; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1800 = opcode == 4'hf ? phv_data_261 : _GEN_1286; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1801 = opcode == 4'hf ? phv_data_260 : _GEN_1287; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1802 = opcode == 4'hf ? phv_data_267 : _GEN_1288; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1803 = opcode == 4'hf ? phv_data_266 : _GEN_1289; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1804 = opcode == 4'hf ? phv_data_265 : _GEN_1290; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1805 = opcode == 4'hf ? phv_data_264 : _GEN_1291; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1806 = opcode == 4'hf ? phv_data_271 : _GEN_1292; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1807 = opcode == 4'hf ? phv_data_270 : _GEN_1293; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1808 = opcode == 4'hf ? phv_data_269 : _GEN_1294; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1809 = opcode == 4'hf ? phv_data_268 : _GEN_1295; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1810 = opcode == 4'hf ? phv_data_275 : _GEN_1296; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1811 = opcode == 4'hf ? phv_data_274 : _GEN_1297; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1812 = opcode == 4'hf ? phv_data_273 : _GEN_1298; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1813 = opcode == 4'hf ? phv_data_272 : _GEN_1299; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1814 = opcode == 4'hf ? phv_data_279 : _GEN_1300; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1815 = opcode == 4'hf ? phv_data_278 : _GEN_1301; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1816 = opcode == 4'hf ? phv_data_277 : _GEN_1302; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1817 = opcode == 4'hf ? phv_data_276 : _GEN_1303; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1818 = opcode == 4'hf ? phv_data_283 : _GEN_1304; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1819 = opcode == 4'hf ? phv_data_282 : _GEN_1305; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1820 = opcode == 4'hf ? phv_data_281 : _GEN_1306; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1821 = opcode == 4'hf ? phv_data_280 : _GEN_1307; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1822 = opcode == 4'hf ? phv_data_287 : _GEN_1308; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1823 = opcode == 4'hf ? phv_data_286 : _GEN_1309; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1824 = opcode == 4'hf ? phv_data_285 : _GEN_1310; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1825 = opcode == 4'hf ? phv_data_284 : _GEN_1311; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1826 = opcode == 4'hf ? phv_data_291 : _GEN_1312; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1827 = opcode == 4'hf ? phv_data_290 : _GEN_1313; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1828 = opcode == 4'hf ? phv_data_289 : _GEN_1314; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1829 = opcode == 4'hf ? phv_data_288 : _GEN_1315; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1830 = opcode == 4'hf ? phv_data_295 : _GEN_1316; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1831 = opcode == 4'hf ? phv_data_294 : _GEN_1317; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1832 = opcode == 4'hf ? phv_data_293 : _GEN_1318; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1833 = opcode == 4'hf ? phv_data_292 : _GEN_1319; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1834 = opcode == 4'hf ? phv_data_299 : _GEN_1320; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1835 = opcode == 4'hf ? phv_data_298 : _GEN_1321; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1836 = opcode == 4'hf ? phv_data_297 : _GEN_1322; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1837 = opcode == 4'hf ? phv_data_296 : _GEN_1323; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1838 = opcode == 4'hf ? phv_data_303 : _GEN_1324; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1839 = opcode == 4'hf ? phv_data_302 : _GEN_1325; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1840 = opcode == 4'hf ? phv_data_301 : _GEN_1326; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1841 = opcode == 4'hf ? phv_data_300 : _GEN_1327; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1842 = opcode == 4'hf ? phv_data_307 : _GEN_1328; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1843 = opcode == 4'hf ? phv_data_306 : _GEN_1329; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1844 = opcode == 4'hf ? phv_data_305 : _GEN_1330; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1845 = opcode == 4'hf ? phv_data_304 : _GEN_1331; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1846 = opcode == 4'hf ? phv_data_311 : _GEN_1332; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1847 = opcode == 4'hf ? phv_data_310 : _GEN_1333; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1848 = opcode == 4'hf ? phv_data_309 : _GEN_1334; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1849 = opcode == 4'hf ? phv_data_308 : _GEN_1335; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1850 = opcode == 4'hf ? phv_data_315 : _GEN_1336; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1851 = opcode == 4'hf ? phv_data_314 : _GEN_1337; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1852 = opcode == 4'hf ? phv_data_313 : _GEN_1338; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1853 = opcode == 4'hf ? phv_data_312 : _GEN_1339; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1854 = opcode == 4'hf ? phv_data_319 : _GEN_1340; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1855 = opcode == 4'hf ? phv_data_318 : _GEN_1341; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1856 = opcode == 4'hf ? phv_data_317 : _GEN_1342; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1857 = opcode == 4'hf ? phv_data_316 : _GEN_1343; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1858 = opcode == 4'hf ? phv_data_323 : _GEN_1344; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1859 = opcode == 4'hf ? phv_data_322 : _GEN_1345; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1860 = opcode == 4'hf ? phv_data_321 : _GEN_1346; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1861 = opcode == 4'hf ? phv_data_320 : _GEN_1347; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1862 = opcode == 4'hf ? phv_data_327 : _GEN_1348; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1863 = opcode == 4'hf ? phv_data_326 : _GEN_1349; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1864 = opcode == 4'hf ? phv_data_325 : _GEN_1350; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1865 = opcode == 4'hf ? phv_data_324 : _GEN_1351; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1866 = opcode == 4'hf ? phv_data_331 : _GEN_1352; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1867 = opcode == 4'hf ? phv_data_330 : _GEN_1353; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1868 = opcode == 4'hf ? phv_data_329 : _GEN_1354; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1869 = opcode == 4'hf ? phv_data_328 : _GEN_1355; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1870 = opcode == 4'hf ? phv_data_335 : _GEN_1356; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1871 = opcode == 4'hf ? phv_data_334 : _GEN_1357; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1872 = opcode == 4'hf ? phv_data_333 : _GEN_1358; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1873 = opcode == 4'hf ? phv_data_332 : _GEN_1359; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1874 = opcode == 4'hf ? phv_data_339 : _GEN_1360; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1875 = opcode == 4'hf ? phv_data_338 : _GEN_1361; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1876 = opcode == 4'hf ? phv_data_337 : _GEN_1362; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1877 = opcode == 4'hf ? phv_data_336 : _GEN_1363; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1878 = opcode == 4'hf ? phv_data_343 : _GEN_1364; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1879 = opcode == 4'hf ? phv_data_342 : _GEN_1365; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1880 = opcode == 4'hf ? phv_data_341 : _GEN_1366; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1881 = opcode == 4'hf ? phv_data_340 : _GEN_1367; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1882 = opcode == 4'hf ? phv_data_347 : _GEN_1368; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1883 = opcode == 4'hf ? phv_data_346 : _GEN_1369; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1884 = opcode == 4'hf ? phv_data_345 : _GEN_1370; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1885 = opcode == 4'hf ? phv_data_344 : _GEN_1371; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1886 = opcode == 4'hf ? phv_data_351 : _GEN_1372; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1887 = opcode == 4'hf ? phv_data_350 : _GEN_1373; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1888 = opcode == 4'hf ? phv_data_349 : _GEN_1374; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1889 = opcode == 4'hf ? phv_data_348 : _GEN_1375; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1890 = opcode == 4'hf ? phv_data_355 : _GEN_1376; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1891 = opcode == 4'hf ? phv_data_354 : _GEN_1377; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1892 = opcode == 4'hf ? phv_data_353 : _GEN_1378; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1893 = opcode == 4'hf ? phv_data_352 : _GEN_1379; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1894 = opcode == 4'hf ? phv_data_359 : _GEN_1380; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1895 = opcode == 4'hf ? phv_data_358 : _GEN_1381; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1896 = opcode == 4'hf ? phv_data_357 : _GEN_1382; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1897 = opcode == 4'hf ? phv_data_356 : _GEN_1383; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1898 = opcode == 4'hf ? phv_data_363 : _GEN_1384; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1899 = opcode == 4'hf ? phv_data_362 : _GEN_1385; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1900 = opcode == 4'hf ? phv_data_361 : _GEN_1386; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1901 = opcode == 4'hf ? phv_data_360 : _GEN_1387; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1902 = opcode == 4'hf ? phv_data_367 : _GEN_1388; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1903 = opcode == 4'hf ? phv_data_366 : _GEN_1389; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1904 = opcode == 4'hf ? phv_data_365 : _GEN_1390; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1905 = opcode == 4'hf ? phv_data_364 : _GEN_1391; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1906 = opcode == 4'hf ? phv_data_371 : _GEN_1392; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1907 = opcode == 4'hf ? phv_data_370 : _GEN_1393; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1908 = opcode == 4'hf ? phv_data_369 : _GEN_1394; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1909 = opcode == 4'hf ? phv_data_368 : _GEN_1395; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1910 = opcode == 4'hf ? phv_data_375 : _GEN_1396; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1911 = opcode == 4'hf ? phv_data_374 : _GEN_1397; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1912 = opcode == 4'hf ? phv_data_373 : _GEN_1398; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1913 = opcode == 4'hf ? phv_data_372 : _GEN_1399; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1914 = opcode == 4'hf ? phv_data_379 : _GEN_1400; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1915 = opcode == 4'hf ? phv_data_378 : _GEN_1401; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1916 = opcode == 4'hf ? phv_data_377 : _GEN_1402; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1917 = opcode == 4'hf ? phv_data_376 : _GEN_1403; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1918 = opcode == 4'hf ? phv_data_383 : _GEN_1404; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1919 = opcode == 4'hf ? phv_data_382 : _GEN_1405; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1920 = opcode == 4'hf ? phv_data_381 : _GEN_1406; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1921 = opcode == 4'hf ? phv_data_380 : _GEN_1407; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1922 = opcode == 4'hf ? phv_data_387 : _GEN_1408; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1923 = opcode == 4'hf ? phv_data_386 : _GEN_1409; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1924 = opcode == 4'hf ? phv_data_385 : _GEN_1410; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1925 = opcode == 4'hf ? phv_data_384 : _GEN_1411; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1926 = opcode == 4'hf ? phv_data_391 : _GEN_1412; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1927 = opcode == 4'hf ? phv_data_390 : _GEN_1413; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1928 = opcode == 4'hf ? phv_data_389 : _GEN_1414; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1929 = opcode == 4'hf ? phv_data_388 : _GEN_1415; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1930 = opcode == 4'hf ? phv_data_395 : _GEN_1416; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1931 = opcode == 4'hf ? phv_data_394 : _GEN_1417; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1932 = opcode == 4'hf ? phv_data_393 : _GEN_1418; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1933 = opcode == 4'hf ? phv_data_392 : _GEN_1419; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1934 = opcode == 4'hf ? phv_data_399 : _GEN_1420; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1935 = opcode == 4'hf ? phv_data_398 : _GEN_1421; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1936 = opcode == 4'hf ? phv_data_397 : _GEN_1422; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1937 = opcode == 4'hf ? phv_data_396 : _GEN_1423; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1938 = opcode == 4'hf ? phv_data_403 : _GEN_1424; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1939 = opcode == 4'hf ? phv_data_402 : _GEN_1425; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1940 = opcode == 4'hf ? phv_data_401 : _GEN_1426; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1941 = opcode == 4'hf ? phv_data_400 : _GEN_1427; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1942 = opcode == 4'hf ? phv_data_407 : _GEN_1428; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1943 = opcode == 4'hf ? phv_data_406 : _GEN_1429; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1944 = opcode == 4'hf ? phv_data_405 : _GEN_1430; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1945 = opcode == 4'hf ? phv_data_404 : _GEN_1431; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1946 = opcode == 4'hf ? phv_data_411 : _GEN_1432; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1947 = opcode == 4'hf ? phv_data_410 : _GEN_1433; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1948 = opcode == 4'hf ? phv_data_409 : _GEN_1434; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1949 = opcode == 4'hf ? phv_data_408 : _GEN_1435; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1950 = opcode == 4'hf ? phv_data_415 : _GEN_1436; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1951 = opcode == 4'hf ? phv_data_414 : _GEN_1437; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1952 = opcode == 4'hf ? phv_data_413 : _GEN_1438; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1953 = opcode == 4'hf ? phv_data_412 : _GEN_1439; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1954 = opcode == 4'hf ? phv_data_419 : _GEN_1440; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1955 = opcode == 4'hf ? phv_data_418 : _GEN_1441; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1956 = opcode == 4'hf ? phv_data_417 : _GEN_1442; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1957 = opcode == 4'hf ? phv_data_416 : _GEN_1443; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1958 = opcode == 4'hf ? phv_data_423 : _GEN_1444; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1959 = opcode == 4'hf ? phv_data_422 : _GEN_1445; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1960 = opcode == 4'hf ? phv_data_421 : _GEN_1446; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1961 = opcode == 4'hf ? phv_data_420 : _GEN_1447; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1962 = opcode == 4'hf ? phv_data_427 : _GEN_1448; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1963 = opcode == 4'hf ? phv_data_426 : _GEN_1449; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1964 = opcode == 4'hf ? phv_data_425 : _GEN_1450; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1965 = opcode == 4'hf ? phv_data_424 : _GEN_1451; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1966 = opcode == 4'hf ? phv_data_431 : _GEN_1452; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1967 = opcode == 4'hf ? phv_data_430 : _GEN_1453; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1968 = opcode == 4'hf ? phv_data_429 : _GEN_1454; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1969 = opcode == 4'hf ? phv_data_428 : _GEN_1455; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1970 = opcode == 4'hf ? phv_data_435 : _GEN_1456; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1971 = opcode == 4'hf ? phv_data_434 : _GEN_1457; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1972 = opcode == 4'hf ? phv_data_433 : _GEN_1458; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1973 = opcode == 4'hf ? phv_data_432 : _GEN_1459; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1974 = opcode == 4'hf ? phv_data_439 : _GEN_1460; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1975 = opcode == 4'hf ? phv_data_438 : _GEN_1461; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1976 = opcode == 4'hf ? phv_data_437 : _GEN_1462; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1977 = opcode == 4'hf ? phv_data_436 : _GEN_1463; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1978 = opcode == 4'hf ? phv_data_443 : _GEN_1464; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1979 = opcode == 4'hf ? phv_data_442 : _GEN_1465; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1980 = opcode == 4'hf ? phv_data_441 : _GEN_1466; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1981 = opcode == 4'hf ? phv_data_440 : _GEN_1467; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1982 = opcode == 4'hf ? phv_data_447 : _GEN_1468; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1983 = opcode == 4'hf ? phv_data_446 : _GEN_1469; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1984 = opcode == 4'hf ? phv_data_445 : _GEN_1470; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1985 = opcode == 4'hf ? phv_data_444 : _GEN_1471; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1986 = opcode == 4'hf ? phv_data_451 : _GEN_1472; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1987 = opcode == 4'hf ? phv_data_450 : _GEN_1473; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1988 = opcode == 4'hf ? phv_data_449 : _GEN_1474; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1989 = opcode == 4'hf ? phv_data_448 : _GEN_1475; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1990 = opcode == 4'hf ? phv_data_455 : _GEN_1476; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1991 = opcode == 4'hf ? phv_data_454 : _GEN_1477; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1992 = opcode == 4'hf ? phv_data_453 : _GEN_1478; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1993 = opcode == 4'hf ? phv_data_452 : _GEN_1479; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1994 = opcode == 4'hf ? phv_data_459 : _GEN_1480; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1995 = opcode == 4'hf ? phv_data_458 : _GEN_1481; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1996 = opcode == 4'hf ? phv_data_457 : _GEN_1482; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1997 = opcode == 4'hf ? phv_data_456 : _GEN_1483; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1998 = opcode == 4'hf ? phv_data_463 : _GEN_1484; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_1999 = opcode == 4'hf ? phv_data_462 : _GEN_1485; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2000 = opcode == 4'hf ? phv_data_461 : _GEN_1486; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2001 = opcode == 4'hf ? phv_data_460 : _GEN_1487; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2002 = opcode == 4'hf ? phv_data_467 : _GEN_1488; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2003 = opcode == 4'hf ? phv_data_466 : _GEN_1489; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2004 = opcode == 4'hf ? phv_data_465 : _GEN_1490; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2005 = opcode == 4'hf ? phv_data_464 : _GEN_1491; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2006 = opcode == 4'hf ? phv_data_471 : _GEN_1492; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2007 = opcode == 4'hf ? phv_data_470 : _GEN_1493; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2008 = opcode == 4'hf ? phv_data_469 : _GEN_1494; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2009 = opcode == 4'hf ? phv_data_468 : _GEN_1495; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2010 = opcode == 4'hf ? phv_data_475 : _GEN_1496; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2011 = opcode == 4'hf ? phv_data_474 : _GEN_1497; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2012 = opcode == 4'hf ? phv_data_473 : _GEN_1498; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2013 = opcode == 4'hf ? phv_data_472 : _GEN_1499; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2014 = opcode == 4'hf ? phv_data_479 : _GEN_1500; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2015 = opcode == 4'hf ? phv_data_478 : _GEN_1501; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2016 = opcode == 4'hf ? phv_data_477 : _GEN_1502; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2017 = opcode == 4'hf ? phv_data_476 : _GEN_1503; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2018 = opcode == 4'hf ? phv_data_483 : _GEN_1504; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2019 = opcode == 4'hf ? phv_data_482 : _GEN_1505; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2020 = opcode == 4'hf ? phv_data_481 : _GEN_1506; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2021 = opcode == 4'hf ? phv_data_480 : _GEN_1507; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2022 = opcode == 4'hf ? phv_data_487 : _GEN_1508; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2023 = opcode == 4'hf ? phv_data_486 : _GEN_1509; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2024 = opcode == 4'hf ? phv_data_485 : _GEN_1510; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2025 = opcode == 4'hf ? phv_data_484 : _GEN_1511; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2026 = opcode == 4'hf ? phv_data_491 : _GEN_1512; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2027 = opcode == 4'hf ? phv_data_490 : _GEN_1513; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2028 = opcode == 4'hf ? phv_data_489 : _GEN_1514; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2029 = opcode == 4'hf ? phv_data_488 : _GEN_1515; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2030 = opcode == 4'hf ? phv_data_495 : _GEN_1516; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2031 = opcode == 4'hf ? phv_data_494 : _GEN_1517; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2032 = opcode == 4'hf ? phv_data_493 : _GEN_1518; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2033 = opcode == 4'hf ? phv_data_492 : _GEN_1519; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2034 = opcode == 4'hf ? phv_data_499 : _GEN_1520; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2035 = opcode == 4'hf ? phv_data_498 : _GEN_1521; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2036 = opcode == 4'hf ? phv_data_497 : _GEN_1522; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2037 = opcode == 4'hf ? phv_data_496 : _GEN_1523; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2038 = opcode == 4'hf ? phv_data_503 : _GEN_1524; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2039 = opcode == 4'hf ? phv_data_502 : _GEN_1525; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2040 = opcode == 4'hf ? phv_data_501 : _GEN_1526; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2041 = opcode == 4'hf ? phv_data_500 : _GEN_1527; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2042 = opcode == 4'hf ? phv_data_507 : _GEN_1528; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2043 = opcode == 4'hf ? phv_data_506 : _GEN_1529; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2044 = opcode == 4'hf ? phv_data_505 : _GEN_1530; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2045 = opcode == 4'hf ? phv_data_504 : _GEN_1531; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2046 = opcode == 4'hf ? phv_data_511 : _GEN_1532; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2047 = opcode == 4'hf ? phv_data_510 : _GEN_1533; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2048 = opcode == 4'hf ? phv_data_509 : _GEN_1534; // @[executor.scala 466:52 executor.scala 450:25]
  wire [7:0] _GEN_2049 = opcode == 4'hf ? phv_data_508 : _GEN_1535; // @[executor.scala 466:52 executor.scala 450:25]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_1 = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8842 = {{2'd0}, dst_offset_1}; // @[executor.scala 473:49]
  wire [7:0] byte_512 = field_1[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2050 = mask_1[0] ? byte_512 : _GEN_1538; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_513 = field_1[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2051 = mask_1[1] ? byte_513 : _GEN_1539; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_514 = field_1[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2052 = mask_1[2] ? byte_514 : _GEN_1540; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_515 = field_1[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_2053 = mask_1[3] ? byte_515 : _GEN_1541; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2054 = _GEN_8842 == 8'h0 ? _GEN_2050 : _GEN_1538; // @[executor.scala 473:84]
  wire [7:0] _GEN_2055 = _GEN_8842 == 8'h0 ? _GEN_2051 : _GEN_1539; // @[executor.scala 473:84]
  wire [7:0] _GEN_2056 = _GEN_8842 == 8'h0 ? _GEN_2052 : _GEN_1540; // @[executor.scala 473:84]
  wire [7:0] _GEN_2057 = _GEN_8842 == 8'h0 ? _GEN_2053 : _GEN_1541; // @[executor.scala 473:84]
  wire [7:0] _GEN_2058 = mask_1[0] ? byte_512 : _GEN_1542; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2059 = mask_1[1] ? byte_513 : _GEN_1543; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2060 = mask_1[2] ? byte_514 : _GEN_1544; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2061 = mask_1[3] ? byte_515 : _GEN_1545; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2062 = _GEN_8842 == 8'h1 ? _GEN_2058 : _GEN_1542; // @[executor.scala 473:84]
  wire [7:0] _GEN_2063 = _GEN_8842 == 8'h1 ? _GEN_2059 : _GEN_1543; // @[executor.scala 473:84]
  wire [7:0] _GEN_2064 = _GEN_8842 == 8'h1 ? _GEN_2060 : _GEN_1544; // @[executor.scala 473:84]
  wire [7:0] _GEN_2065 = _GEN_8842 == 8'h1 ? _GEN_2061 : _GEN_1545; // @[executor.scala 473:84]
  wire [7:0] _GEN_2066 = mask_1[0] ? byte_512 : _GEN_1546; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2067 = mask_1[1] ? byte_513 : _GEN_1547; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2068 = mask_1[2] ? byte_514 : _GEN_1548; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2069 = mask_1[3] ? byte_515 : _GEN_1549; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2070 = _GEN_8842 == 8'h2 ? _GEN_2066 : _GEN_1546; // @[executor.scala 473:84]
  wire [7:0] _GEN_2071 = _GEN_8842 == 8'h2 ? _GEN_2067 : _GEN_1547; // @[executor.scala 473:84]
  wire [7:0] _GEN_2072 = _GEN_8842 == 8'h2 ? _GEN_2068 : _GEN_1548; // @[executor.scala 473:84]
  wire [7:0] _GEN_2073 = _GEN_8842 == 8'h2 ? _GEN_2069 : _GEN_1549; // @[executor.scala 473:84]
  wire [7:0] _GEN_2074 = mask_1[0] ? byte_512 : _GEN_1550; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2075 = mask_1[1] ? byte_513 : _GEN_1551; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2076 = mask_1[2] ? byte_514 : _GEN_1552; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2077 = mask_1[3] ? byte_515 : _GEN_1553; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2078 = _GEN_8842 == 8'h3 ? _GEN_2074 : _GEN_1550; // @[executor.scala 473:84]
  wire [7:0] _GEN_2079 = _GEN_8842 == 8'h3 ? _GEN_2075 : _GEN_1551; // @[executor.scala 473:84]
  wire [7:0] _GEN_2080 = _GEN_8842 == 8'h3 ? _GEN_2076 : _GEN_1552; // @[executor.scala 473:84]
  wire [7:0] _GEN_2081 = _GEN_8842 == 8'h3 ? _GEN_2077 : _GEN_1553; // @[executor.scala 473:84]
  wire [7:0] _GEN_2082 = mask_1[0] ? byte_512 : _GEN_1554; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2083 = mask_1[1] ? byte_513 : _GEN_1555; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2084 = mask_1[2] ? byte_514 : _GEN_1556; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2085 = mask_1[3] ? byte_515 : _GEN_1557; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2086 = _GEN_8842 == 8'h4 ? _GEN_2082 : _GEN_1554; // @[executor.scala 473:84]
  wire [7:0] _GEN_2087 = _GEN_8842 == 8'h4 ? _GEN_2083 : _GEN_1555; // @[executor.scala 473:84]
  wire [7:0] _GEN_2088 = _GEN_8842 == 8'h4 ? _GEN_2084 : _GEN_1556; // @[executor.scala 473:84]
  wire [7:0] _GEN_2089 = _GEN_8842 == 8'h4 ? _GEN_2085 : _GEN_1557; // @[executor.scala 473:84]
  wire [7:0] _GEN_2090 = mask_1[0] ? byte_512 : _GEN_1558; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2091 = mask_1[1] ? byte_513 : _GEN_1559; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2092 = mask_1[2] ? byte_514 : _GEN_1560; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2093 = mask_1[3] ? byte_515 : _GEN_1561; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2094 = _GEN_8842 == 8'h5 ? _GEN_2090 : _GEN_1558; // @[executor.scala 473:84]
  wire [7:0] _GEN_2095 = _GEN_8842 == 8'h5 ? _GEN_2091 : _GEN_1559; // @[executor.scala 473:84]
  wire [7:0] _GEN_2096 = _GEN_8842 == 8'h5 ? _GEN_2092 : _GEN_1560; // @[executor.scala 473:84]
  wire [7:0] _GEN_2097 = _GEN_8842 == 8'h5 ? _GEN_2093 : _GEN_1561; // @[executor.scala 473:84]
  wire [7:0] _GEN_2098 = mask_1[0] ? byte_512 : _GEN_1562; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2099 = mask_1[1] ? byte_513 : _GEN_1563; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2100 = mask_1[2] ? byte_514 : _GEN_1564; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2101 = mask_1[3] ? byte_515 : _GEN_1565; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2102 = _GEN_8842 == 8'h6 ? _GEN_2098 : _GEN_1562; // @[executor.scala 473:84]
  wire [7:0] _GEN_2103 = _GEN_8842 == 8'h6 ? _GEN_2099 : _GEN_1563; // @[executor.scala 473:84]
  wire [7:0] _GEN_2104 = _GEN_8842 == 8'h6 ? _GEN_2100 : _GEN_1564; // @[executor.scala 473:84]
  wire [7:0] _GEN_2105 = _GEN_8842 == 8'h6 ? _GEN_2101 : _GEN_1565; // @[executor.scala 473:84]
  wire [7:0] _GEN_2106 = mask_1[0] ? byte_512 : _GEN_1566; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2107 = mask_1[1] ? byte_513 : _GEN_1567; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2108 = mask_1[2] ? byte_514 : _GEN_1568; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2109 = mask_1[3] ? byte_515 : _GEN_1569; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2110 = _GEN_8842 == 8'h7 ? _GEN_2106 : _GEN_1566; // @[executor.scala 473:84]
  wire [7:0] _GEN_2111 = _GEN_8842 == 8'h7 ? _GEN_2107 : _GEN_1567; // @[executor.scala 473:84]
  wire [7:0] _GEN_2112 = _GEN_8842 == 8'h7 ? _GEN_2108 : _GEN_1568; // @[executor.scala 473:84]
  wire [7:0] _GEN_2113 = _GEN_8842 == 8'h7 ? _GEN_2109 : _GEN_1569; // @[executor.scala 473:84]
  wire [7:0] _GEN_2114 = mask_1[0] ? byte_512 : _GEN_1570; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2115 = mask_1[1] ? byte_513 : _GEN_1571; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2116 = mask_1[2] ? byte_514 : _GEN_1572; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2117 = mask_1[3] ? byte_515 : _GEN_1573; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2118 = _GEN_8842 == 8'h8 ? _GEN_2114 : _GEN_1570; // @[executor.scala 473:84]
  wire [7:0] _GEN_2119 = _GEN_8842 == 8'h8 ? _GEN_2115 : _GEN_1571; // @[executor.scala 473:84]
  wire [7:0] _GEN_2120 = _GEN_8842 == 8'h8 ? _GEN_2116 : _GEN_1572; // @[executor.scala 473:84]
  wire [7:0] _GEN_2121 = _GEN_8842 == 8'h8 ? _GEN_2117 : _GEN_1573; // @[executor.scala 473:84]
  wire [7:0] _GEN_2122 = mask_1[0] ? byte_512 : _GEN_1574; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2123 = mask_1[1] ? byte_513 : _GEN_1575; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2124 = mask_1[2] ? byte_514 : _GEN_1576; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2125 = mask_1[3] ? byte_515 : _GEN_1577; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2126 = _GEN_8842 == 8'h9 ? _GEN_2122 : _GEN_1574; // @[executor.scala 473:84]
  wire [7:0] _GEN_2127 = _GEN_8842 == 8'h9 ? _GEN_2123 : _GEN_1575; // @[executor.scala 473:84]
  wire [7:0] _GEN_2128 = _GEN_8842 == 8'h9 ? _GEN_2124 : _GEN_1576; // @[executor.scala 473:84]
  wire [7:0] _GEN_2129 = _GEN_8842 == 8'h9 ? _GEN_2125 : _GEN_1577; // @[executor.scala 473:84]
  wire [7:0] _GEN_2130 = mask_1[0] ? byte_512 : _GEN_1578; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2131 = mask_1[1] ? byte_513 : _GEN_1579; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2132 = mask_1[2] ? byte_514 : _GEN_1580; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2133 = mask_1[3] ? byte_515 : _GEN_1581; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2134 = _GEN_8842 == 8'ha ? _GEN_2130 : _GEN_1578; // @[executor.scala 473:84]
  wire [7:0] _GEN_2135 = _GEN_8842 == 8'ha ? _GEN_2131 : _GEN_1579; // @[executor.scala 473:84]
  wire [7:0] _GEN_2136 = _GEN_8842 == 8'ha ? _GEN_2132 : _GEN_1580; // @[executor.scala 473:84]
  wire [7:0] _GEN_2137 = _GEN_8842 == 8'ha ? _GEN_2133 : _GEN_1581; // @[executor.scala 473:84]
  wire [7:0] _GEN_2138 = mask_1[0] ? byte_512 : _GEN_1582; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2139 = mask_1[1] ? byte_513 : _GEN_1583; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2140 = mask_1[2] ? byte_514 : _GEN_1584; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2141 = mask_1[3] ? byte_515 : _GEN_1585; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2142 = _GEN_8842 == 8'hb ? _GEN_2138 : _GEN_1582; // @[executor.scala 473:84]
  wire [7:0] _GEN_2143 = _GEN_8842 == 8'hb ? _GEN_2139 : _GEN_1583; // @[executor.scala 473:84]
  wire [7:0] _GEN_2144 = _GEN_8842 == 8'hb ? _GEN_2140 : _GEN_1584; // @[executor.scala 473:84]
  wire [7:0] _GEN_2145 = _GEN_8842 == 8'hb ? _GEN_2141 : _GEN_1585; // @[executor.scala 473:84]
  wire [7:0] _GEN_2146 = mask_1[0] ? byte_512 : _GEN_1586; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2147 = mask_1[1] ? byte_513 : _GEN_1587; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2148 = mask_1[2] ? byte_514 : _GEN_1588; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2149 = mask_1[3] ? byte_515 : _GEN_1589; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2150 = _GEN_8842 == 8'hc ? _GEN_2146 : _GEN_1586; // @[executor.scala 473:84]
  wire [7:0] _GEN_2151 = _GEN_8842 == 8'hc ? _GEN_2147 : _GEN_1587; // @[executor.scala 473:84]
  wire [7:0] _GEN_2152 = _GEN_8842 == 8'hc ? _GEN_2148 : _GEN_1588; // @[executor.scala 473:84]
  wire [7:0] _GEN_2153 = _GEN_8842 == 8'hc ? _GEN_2149 : _GEN_1589; // @[executor.scala 473:84]
  wire [7:0] _GEN_2154 = mask_1[0] ? byte_512 : _GEN_1590; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2155 = mask_1[1] ? byte_513 : _GEN_1591; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2156 = mask_1[2] ? byte_514 : _GEN_1592; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2157 = mask_1[3] ? byte_515 : _GEN_1593; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2158 = _GEN_8842 == 8'hd ? _GEN_2154 : _GEN_1590; // @[executor.scala 473:84]
  wire [7:0] _GEN_2159 = _GEN_8842 == 8'hd ? _GEN_2155 : _GEN_1591; // @[executor.scala 473:84]
  wire [7:0] _GEN_2160 = _GEN_8842 == 8'hd ? _GEN_2156 : _GEN_1592; // @[executor.scala 473:84]
  wire [7:0] _GEN_2161 = _GEN_8842 == 8'hd ? _GEN_2157 : _GEN_1593; // @[executor.scala 473:84]
  wire [7:0] _GEN_2162 = mask_1[0] ? byte_512 : _GEN_1594; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2163 = mask_1[1] ? byte_513 : _GEN_1595; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2164 = mask_1[2] ? byte_514 : _GEN_1596; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2165 = mask_1[3] ? byte_515 : _GEN_1597; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2166 = _GEN_8842 == 8'he ? _GEN_2162 : _GEN_1594; // @[executor.scala 473:84]
  wire [7:0] _GEN_2167 = _GEN_8842 == 8'he ? _GEN_2163 : _GEN_1595; // @[executor.scala 473:84]
  wire [7:0] _GEN_2168 = _GEN_8842 == 8'he ? _GEN_2164 : _GEN_1596; // @[executor.scala 473:84]
  wire [7:0] _GEN_2169 = _GEN_8842 == 8'he ? _GEN_2165 : _GEN_1597; // @[executor.scala 473:84]
  wire [7:0] _GEN_2170 = mask_1[0] ? byte_512 : _GEN_1598; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2171 = mask_1[1] ? byte_513 : _GEN_1599; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2172 = mask_1[2] ? byte_514 : _GEN_1600; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2173 = mask_1[3] ? byte_515 : _GEN_1601; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2174 = _GEN_8842 == 8'hf ? _GEN_2170 : _GEN_1598; // @[executor.scala 473:84]
  wire [7:0] _GEN_2175 = _GEN_8842 == 8'hf ? _GEN_2171 : _GEN_1599; // @[executor.scala 473:84]
  wire [7:0] _GEN_2176 = _GEN_8842 == 8'hf ? _GEN_2172 : _GEN_1600; // @[executor.scala 473:84]
  wire [7:0] _GEN_2177 = _GEN_8842 == 8'hf ? _GEN_2173 : _GEN_1601; // @[executor.scala 473:84]
  wire [7:0] _GEN_2178 = mask_1[0] ? byte_512 : _GEN_1602; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2179 = mask_1[1] ? byte_513 : _GEN_1603; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2180 = mask_1[2] ? byte_514 : _GEN_1604; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2181 = mask_1[3] ? byte_515 : _GEN_1605; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2182 = _GEN_8842 == 8'h10 ? _GEN_2178 : _GEN_1602; // @[executor.scala 473:84]
  wire [7:0] _GEN_2183 = _GEN_8842 == 8'h10 ? _GEN_2179 : _GEN_1603; // @[executor.scala 473:84]
  wire [7:0] _GEN_2184 = _GEN_8842 == 8'h10 ? _GEN_2180 : _GEN_1604; // @[executor.scala 473:84]
  wire [7:0] _GEN_2185 = _GEN_8842 == 8'h10 ? _GEN_2181 : _GEN_1605; // @[executor.scala 473:84]
  wire [7:0] _GEN_2186 = mask_1[0] ? byte_512 : _GEN_1606; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2187 = mask_1[1] ? byte_513 : _GEN_1607; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2188 = mask_1[2] ? byte_514 : _GEN_1608; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2189 = mask_1[3] ? byte_515 : _GEN_1609; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2190 = _GEN_8842 == 8'h11 ? _GEN_2186 : _GEN_1606; // @[executor.scala 473:84]
  wire [7:0] _GEN_2191 = _GEN_8842 == 8'h11 ? _GEN_2187 : _GEN_1607; // @[executor.scala 473:84]
  wire [7:0] _GEN_2192 = _GEN_8842 == 8'h11 ? _GEN_2188 : _GEN_1608; // @[executor.scala 473:84]
  wire [7:0] _GEN_2193 = _GEN_8842 == 8'h11 ? _GEN_2189 : _GEN_1609; // @[executor.scala 473:84]
  wire [7:0] _GEN_2194 = mask_1[0] ? byte_512 : _GEN_1610; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2195 = mask_1[1] ? byte_513 : _GEN_1611; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2196 = mask_1[2] ? byte_514 : _GEN_1612; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2197 = mask_1[3] ? byte_515 : _GEN_1613; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2198 = _GEN_8842 == 8'h12 ? _GEN_2194 : _GEN_1610; // @[executor.scala 473:84]
  wire [7:0] _GEN_2199 = _GEN_8842 == 8'h12 ? _GEN_2195 : _GEN_1611; // @[executor.scala 473:84]
  wire [7:0] _GEN_2200 = _GEN_8842 == 8'h12 ? _GEN_2196 : _GEN_1612; // @[executor.scala 473:84]
  wire [7:0] _GEN_2201 = _GEN_8842 == 8'h12 ? _GEN_2197 : _GEN_1613; // @[executor.scala 473:84]
  wire [7:0] _GEN_2202 = mask_1[0] ? byte_512 : _GEN_1614; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2203 = mask_1[1] ? byte_513 : _GEN_1615; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2204 = mask_1[2] ? byte_514 : _GEN_1616; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2205 = mask_1[3] ? byte_515 : _GEN_1617; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2206 = _GEN_8842 == 8'h13 ? _GEN_2202 : _GEN_1614; // @[executor.scala 473:84]
  wire [7:0] _GEN_2207 = _GEN_8842 == 8'h13 ? _GEN_2203 : _GEN_1615; // @[executor.scala 473:84]
  wire [7:0] _GEN_2208 = _GEN_8842 == 8'h13 ? _GEN_2204 : _GEN_1616; // @[executor.scala 473:84]
  wire [7:0] _GEN_2209 = _GEN_8842 == 8'h13 ? _GEN_2205 : _GEN_1617; // @[executor.scala 473:84]
  wire [7:0] _GEN_2210 = mask_1[0] ? byte_512 : _GEN_1618; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2211 = mask_1[1] ? byte_513 : _GEN_1619; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2212 = mask_1[2] ? byte_514 : _GEN_1620; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2213 = mask_1[3] ? byte_515 : _GEN_1621; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2214 = _GEN_8842 == 8'h14 ? _GEN_2210 : _GEN_1618; // @[executor.scala 473:84]
  wire [7:0] _GEN_2215 = _GEN_8842 == 8'h14 ? _GEN_2211 : _GEN_1619; // @[executor.scala 473:84]
  wire [7:0] _GEN_2216 = _GEN_8842 == 8'h14 ? _GEN_2212 : _GEN_1620; // @[executor.scala 473:84]
  wire [7:0] _GEN_2217 = _GEN_8842 == 8'h14 ? _GEN_2213 : _GEN_1621; // @[executor.scala 473:84]
  wire [7:0] _GEN_2218 = mask_1[0] ? byte_512 : _GEN_1622; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2219 = mask_1[1] ? byte_513 : _GEN_1623; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2220 = mask_1[2] ? byte_514 : _GEN_1624; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2221 = mask_1[3] ? byte_515 : _GEN_1625; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2222 = _GEN_8842 == 8'h15 ? _GEN_2218 : _GEN_1622; // @[executor.scala 473:84]
  wire [7:0] _GEN_2223 = _GEN_8842 == 8'h15 ? _GEN_2219 : _GEN_1623; // @[executor.scala 473:84]
  wire [7:0] _GEN_2224 = _GEN_8842 == 8'h15 ? _GEN_2220 : _GEN_1624; // @[executor.scala 473:84]
  wire [7:0] _GEN_2225 = _GEN_8842 == 8'h15 ? _GEN_2221 : _GEN_1625; // @[executor.scala 473:84]
  wire [7:0] _GEN_2226 = mask_1[0] ? byte_512 : _GEN_1626; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2227 = mask_1[1] ? byte_513 : _GEN_1627; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2228 = mask_1[2] ? byte_514 : _GEN_1628; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2229 = mask_1[3] ? byte_515 : _GEN_1629; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2230 = _GEN_8842 == 8'h16 ? _GEN_2226 : _GEN_1626; // @[executor.scala 473:84]
  wire [7:0] _GEN_2231 = _GEN_8842 == 8'h16 ? _GEN_2227 : _GEN_1627; // @[executor.scala 473:84]
  wire [7:0] _GEN_2232 = _GEN_8842 == 8'h16 ? _GEN_2228 : _GEN_1628; // @[executor.scala 473:84]
  wire [7:0] _GEN_2233 = _GEN_8842 == 8'h16 ? _GEN_2229 : _GEN_1629; // @[executor.scala 473:84]
  wire [7:0] _GEN_2234 = mask_1[0] ? byte_512 : _GEN_1630; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2235 = mask_1[1] ? byte_513 : _GEN_1631; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2236 = mask_1[2] ? byte_514 : _GEN_1632; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2237 = mask_1[3] ? byte_515 : _GEN_1633; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2238 = _GEN_8842 == 8'h17 ? _GEN_2234 : _GEN_1630; // @[executor.scala 473:84]
  wire [7:0] _GEN_2239 = _GEN_8842 == 8'h17 ? _GEN_2235 : _GEN_1631; // @[executor.scala 473:84]
  wire [7:0] _GEN_2240 = _GEN_8842 == 8'h17 ? _GEN_2236 : _GEN_1632; // @[executor.scala 473:84]
  wire [7:0] _GEN_2241 = _GEN_8842 == 8'h17 ? _GEN_2237 : _GEN_1633; // @[executor.scala 473:84]
  wire [7:0] _GEN_2242 = mask_1[0] ? byte_512 : _GEN_1634; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2243 = mask_1[1] ? byte_513 : _GEN_1635; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2244 = mask_1[2] ? byte_514 : _GEN_1636; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2245 = mask_1[3] ? byte_515 : _GEN_1637; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2246 = _GEN_8842 == 8'h18 ? _GEN_2242 : _GEN_1634; // @[executor.scala 473:84]
  wire [7:0] _GEN_2247 = _GEN_8842 == 8'h18 ? _GEN_2243 : _GEN_1635; // @[executor.scala 473:84]
  wire [7:0] _GEN_2248 = _GEN_8842 == 8'h18 ? _GEN_2244 : _GEN_1636; // @[executor.scala 473:84]
  wire [7:0] _GEN_2249 = _GEN_8842 == 8'h18 ? _GEN_2245 : _GEN_1637; // @[executor.scala 473:84]
  wire [7:0] _GEN_2250 = mask_1[0] ? byte_512 : _GEN_1638; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2251 = mask_1[1] ? byte_513 : _GEN_1639; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2252 = mask_1[2] ? byte_514 : _GEN_1640; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2253 = mask_1[3] ? byte_515 : _GEN_1641; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2254 = _GEN_8842 == 8'h19 ? _GEN_2250 : _GEN_1638; // @[executor.scala 473:84]
  wire [7:0] _GEN_2255 = _GEN_8842 == 8'h19 ? _GEN_2251 : _GEN_1639; // @[executor.scala 473:84]
  wire [7:0] _GEN_2256 = _GEN_8842 == 8'h19 ? _GEN_2252 : _GEN_1640; // @[executor.scala 473:84]
  wire [7:0] _GEN_2257 = _GEN_8842 == 8'h19 ? _GEN_2253 : _GEN_1641; // @[executor.scala 473:84]
  wire [7:0] _GEN_2258 = mask_1[0] ? byte_512 : _GEN_1642; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2259 = mask_1[1] ? byte_513 : _GEN_1643; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2260 = mask_1[2] ? byte_514 : _GEN_1644; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2261 = mask_1[3] ? byte_515 : _GEN_1645; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2262 = _GEN_8842 == 8'h1a ? _GEN_2258 : _GEN_1642; // @[executor.scala 473:84]
  wire [7:0] _GEN_2263 = _GEN_8842 == 8'h1a ? _GEN_2259 : _GEN_1643; // @[executor.scala 473:84]
  wire [7:0] _GEN_2264 = _GEN_8842 == 8'h1a ? _GEN_2260 : _GEN_1644; // @[executor.scala 473:84]
  wire [7:0] _GEN_2265 = _GEN_8842 == 8'h1a ? _GEN_2261 : _GEN_1645; // @[executor.scala 473:84]
  wire [7:0] _GEN_2266 = mask_1[0] ? byte_512 : _GEN_1646; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2267 = mask_1[1] ? byte_513 : _GEN_1647; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2268 = mask_1[2] ? byte_514 : _GEN_1648; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2269 = mask_1[3] ? byte_515 : _GEN_1649; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2270 = _GEN_8842 == 8'h1b ? _GEN_2266 : _GEN_1646; // @[executor.scala 473:84]
  wire [7:0] _GEN_2271 = _GEN_8842 == 8'h1b ? _GEN_2267 : _GEN_1647; // @[executor.scala 473:84]
  wire [7:0] _GEN_2272 = _GEN_8842 == 8'h1b ? _GEN_2268 : _GEN_1648; // @[executor.scala 473:84]
  wire [7:0] _GEN_2273 = _GEN_8842 == 8'h1b ? _GEN_2269 : _GEN_1649; // @[executor.scala 473:84]
  wire [7:0] _GEN_2274 = mask_1[0] ? byte_512 : _GEN_1650; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2275 = mask_1[1] ? byte_513 : _GEN_1651; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2276 = mask_1[2] ? byte_514 : _GEN_1652; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2277 = mask_1[3] ? byte_515 : _GEN_1653; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2278 = _GEN_8842 == 8'h1c ? _GEN_2274 : _GEN_1650; // @[executor.scala 473:84]
  wire [7:0] _GEN_2279 = _GEN_8842 == 8'h1c ? _GEN_2275 : _GEN_1651; // @[executor.scala 473:84]
  wire [7:0] _GEN_2280 = _GEN_8842 == 8'h1c ? _GEN_2276 : _GEN_1652; // @[executor.scala 473:84]
  wire [7:0] _GEN_2281 = _GEN_8842 == 8'h1c ? _GEN_2277 : _GEN_1653; // @[executor.scala 473:84]
  wire [7:0] _GEN_2282 = mask_1[0] ? byte_512 : _GEN_1654; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2283 = mask_1[1] ? byte_513 : _GEN_1655; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2284 = mask_1[2] ? byte_514 : _GEN_1656; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2285 = mask_1[3] ? byte_515 : _GEN_1657; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2286 = _GEN_8842 == 8'h1d ? _GEN_2282 : _GEN_1654; // @[executor.scala 473:84]
  wire [7:0] _GEN_2287 = _GEN_8842 == 8'h1d ? _GEN_2283 : _GEN_1655; // @[executor.scala 473:84]
  wire [7:0] _GEN_2288 = _GEN_8842 == 8'h1d ? _GEN_2284 : _GEN_1656; // @[executor.scala 473:84]
  wire [7:0] _GEN_2289 = _GEN_8842 == 8'h1d ? _GEN_2285 : _GEN_1657; // @[executor.scala 473:84]
  wire [7:0] _GEN_2290 = mask_1[0] ? byte_512 : _GEN_1658; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2291 = mask_1[1] ? byte_513 : _GEN_1659; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2292 = mask_1[2] ? byte_514 : _GEN_1660; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2293 = mask_1[3] ? byte_515 : _GEN_1661; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2294 = _GEN_8842 == 8'h1e ? _GEN_2290 : _GEN_1658; // @[executor.scala 473:84]
  wire [7:0] _GEN_2295 = _GEN_8842 == 8'h1e ? _GEN_2291 : _GEN_1659; // @[executor.scala 473:84]
  wire [7:0] _GEN_2296 = _GEN_8842 == 8'h1e ? _GEN_2292 : _GEN_1660; // @[executor.scala 473:84]
  wire [7:0] _GEN_2297 = _GEN_8842 == 8'h1e ? _GEN_2293 : _GEN_1661; // @[executor.scala 473:84]
  wire [7:0] _GEN_2298 = mask_1[0] ? byte_512 : _GEN_1662; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2299 = mask_1[1] ? byte_513 : _GEN_1663; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2300 = mask_1[2] ? byte_514 : _GEN_1664; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2301 = mask_1[3] ? byte_515 : _GEN_1665; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2302 = _GEN_8842 == 8'h1f ? _GEN_2298 : _GEN_1662; // @[executor.scala 473:84]
  wire [7:0] _GEN_2303 = _GEN_8842 == 8'h1f ? _GEN_2299 : _GEN_1663; // @[executor.scala 473:84]
  wire [7:0] _GEN_2304 = _GEN_8842 == 8'h1f ? _GEN_2300 : _GEN_1664; // @[executor.scala 473:84]
  wire [7:0] _GEN_2305 = _GEN_8842 == 8'h1f ? _GEN_2301 : _GEN_1665; // @[executor.scala 473:84]
  wire [7:0] _GEN_2306 = mask_1[0] ? byte_512 : _GEN_1666; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2307 = mask_1[1] ? byte_513 : _GEN_1667; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2308 = mask_1[2] ? byte_514 : _GEN_1668; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2309 = mask_1[3] ? byte_515 : _GEN_1669; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2310 = _GEN_8842 == 8'h20 ? _GEN_2306 : _GEN_1666; // @[executor.scala 473:84]
  wire [7:0] _GEN_2311 = _GEN_8842 == 8'h20 ? _GEN_2307 : _GEN_1667; // @[executor.scala 473:84]
  wire [7:0] _GEN_2312 = _GEN_8842 == 8'h20 ? _GEN_2308 : _GEN_1668; // @[executor.scala 473:84]
  wire [7:0] _GEN_2313 = _GEN_8842 == 8'h20 ? _GEN_2309 : _GEN_1669; // @[executor.scala 473:84]
  wire [7:0] _GEN_2314 = mask_1[0] ? byte_512 : _GEN_1670; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2315 = mask_1[1] ? byte_513 : _GEN_1671; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2316 = mask_1[2] ? byte_514 : _GEN_1672; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2317 = mask_1[3] ? byte_515 : _GEN_1673; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2318 = _GEN_8842 == 8'h21 ? _GEN_2314 : _GEN_1670; // @[executor.scala 473:84]
  wire [7:0] _GEN_2319 = _GEN_8842 == 8'h21 ? _GEN_2315 : _GEN_1671; // @[executor.scala 473:84]
  wire [7:0] _GEN_2320 = _GEN_8842 == 8'h21 ? _GEN_2316 : _GEN_1672; // @[executor.scala 473:84]
  wire [7:0] _GEN_2321 = _GEN_8842 == 8'h21 ? _GEN_2317 : _GEN_1673; // @[executor.scala 473:84]
  wire [7:0] _GEN_2322 = mask_1[0] ? byte_512 : _GEN_1674; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2323 = mask_1[1] ? byte_513 : _GEN_1675; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2324 = mask_1[2] ? byte_514 : _GEN_1676; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2325 = mask_1[3] ? byte_515 : _GEN_1677; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2326 = _GEN_8842 == 8'h22 ? _GEN_2322 : _GEN_1674; // @[executor.scala 473:84]
  wire [7:0] _GEN_2327 = _GEN_8842 == 8'h22 ? _GEN_2323 : _GEN_1675; // @[executor.scala 473:84]
  wire [7:0] _GEN_2328 = _GEN_8842 == 8'h22 ? _GEN_2324 : _GEN_1676; // @[executor.scala 473:84]
  wire [7:0] _GEN_2329 = _GEN_8842 == 8'h22 ? _GEN_2325 : _GEN_1677; // @[executor.scala 473:84]
  wire [7:0] _GEN_2330 = mask_1[0] ? byte_512 : _GEN_1678; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2331 = mask_1[1] ? byte_513 : _GEN_1679; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2332 = mask_1[2] ? byte_514 : _GEN_1680; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2333 = mask_1[3] ? byte_515 : _GEN_1681; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2334 = _GEN_8842 == 8'h23 ? _GEN_2330 : _GEN_1678; // @[executor.scala 473:84]
  wire [7:0] _GEN_2335 = _GEN_8842 == 8'h23 ? _GEN_2331 : _GEN_1679; // @[executor.scala 473:84]
  wire [7:0] _GEN_2336 = _GEN_8842 == 8'h23 ? _GEN_2332 : _GEN_1680; // @[executor.scala 473:84]
  wire [7:0] _GEN_2337 = _GEN_8842 == 8'h23 ? _GEN_2333 : _GEN_1681; // @[executor.scala 473:84]
  wire [7:0] _GEN_2338 = mask_1[0] ? byte_512 : _GEN_1682; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2339 = mask_1[1] ? byte_513 : _GEN_1683; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2340 = mask_1[2] ? byte_514 : _GEN_1684; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2341 = mask_1[3] ? byte_515 : _GEN_1685; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2342 = _GEN_8842 == 8'h24 ? _GEN_2338 : _GEN_1682; // @[executor.scala 473:84]
  wire [7:0] _GEN_2343 = _GEN_8842 == 8'h24 ? _GEN_2339 : _GEN_1683; // @[executor.scala 473:84]
  wire [7:0] _GEN_2344 = _GEN_8842 == 8'h24 ? _GEN_2340 : _GEN_1684; // @[executor.scala 473:84]
  wire [7:0] _GEN_2345 = _GEN_8842 == 8'h24 ? _GEN_2341 : _GEN_1685; // @[executor.scala 473:84]
  wire [7:0] _GEN_2346 = mask_1[0] ? byte_512 : _GEN_1686; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2347 = mask_1[1] ? byte_513 : _GEN_1687; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2348 = mask_1[2] ? byte_514 : _GEN_1688; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2349 = mask_1[3] ? byte_515 : _GEN_1689; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2350 = _GEN_8842 == 8'h25 ? _GEN_2346 : _GEN_1686; // @[executor.scala 473:84]
  wire [7:0] _GEN_2351 = _GEN_8842 == 8'h25 ? _GEN_2347 : _GEN_1687; // @[executor.scala 473:84]
  wire [7:0] _GEN_2352 = _GEN_8842 == 8'h25 ? _GEN_2348 : _GEN_1688; // @[executor.scala 473:84]
  wire [7:0] _GEN_2353 = _GEN_8842 == 8'h25 ? _GEN_2349 : _GEN_1689; // @[executor.scala 473:84]
  wire [7:0] _GEN_2354 = mask_1[0] ? byte_512 : _GEN_1690; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2355 = mask_1[1] ? byte_513 : _GEN_1691; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2356 = mask_1[2] ? byte_514 : _GEN_1692; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2357 = mask_1[3] ? byte_515 : _GEN_1693; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2358 = _GEN_8842 == 8'h26 ? _GEN_2354 : _GEN_1690; // @[executor.scala 473:84]
  wire [7:0] _GEN_2359 = _GEN_8842 == 8'h26 ? _GEN_2355 : _GEN_1691; // @[executor.scala 473:84]
  wire [7:0] _GEN_2360 = _GEN_8842 == 8'h26 ? _GEN_2356 : _GEN_1692; // @[executor.scala 473:84]
  wire [7:0] _GEN_2361 = _GEN_8842 == 8'h26 ? _GEN_2357 : _GEN_1693; // @[executor.scala 473:84]
  wire [7:0] _GEN_2362 = mask_1[0] ? byte_512 : _GEN_1694; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2363 = mask_1[1] ? byte_513 : _GEN_1695; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2364 = mask_1[2] ? byte_514 : _GEN_1696; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2365 = mask_1[3] ? byte_515 : _GEN_1697; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2366 = _GEN_8842 == 8'h27 ? _GEN_2362 : _GEN_1694; // @[executor.scala 473:84]
  wire [7:0] _GEN_2367 = _GEN_8842 == 8'h27 ? _GEN_2363 : _GEN_1695; // @[executor.scala 473:84]
  wire [7:0] _GEN_2368 = _GEN_8842 == 8'h27 ? _GEN_2364 : _GEN_1696; // @[executor.scala 473:84]
  wire [7:0] _GEN_2369 = _GEN_8842 == 8'h27 ? _GEN_2365 : _GEN_1697; // @[executor.scala 473:84]
  wire [7:0] _GEN_2370 = mask_1[0] ? byte_512 : _GEN_1698; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2371 = mask_1[1] ? byte_513 : _GEN_1699; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2372 = mask_1[2] ? byte_514 : _GEN_1700; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2373 = mask_1[3] ? byte_515 : _GEN_1701; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2374 = _GEN_8842 == 8'h28 ? _GEN_2370 : _GEN_1698; // @[executor.scala 473:84]
  wire [7:0] _GEN_2375 = _GEN_8842 == 8'h28 ? _GEN_2371 : _GEN_1699; // @[executor.scala 473:84]
  wire [7:0] _GEN_2376 = _GEN_8842 == 8'h28 ? _GEN_2372 : _GEN_1700; // @[executor.scala 473:84]
  wire [7:0] _GEN_2377 = _GEN_8842 == 8'h28 ? _GEN_2373 : _GEN_1701; // @[executor.scala 473:84]
  wire [7:0] _GEN_2378 = mask_1[0] ? byte_512 : _GEN_1702; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2379 = mask_1[1] ? byte_513 : _GEN_1703; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2380 = mask_1[2] ? byte_514 : _GEN_1704; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2381 = mask_1[3] ? byte_515 : _GEN_1705; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2382 = _GEN_8842 == 8'h29 ? _GEN_2378 : _GEN_1702; // @[executor.scala 473:84]
  wire [7:0] _GEN_2383 = _GEN_8842 == 8'h29 ? _GEN_2379 : _GEN_1703; // @[executor.scala 473:84]
  wire [7:0] _GEN_2384 = _GEN_8842 == 8'h29 ? _GEN_2380 : _GEN_1704; // @[executor.scala 473:84]
  wire [7:0] _GEN_2385 = _GEN_8842 == 8'h29 ? _GEN_2381 : _GEN_1705; // @[executor.scala 473:84]
  wire [7:0] _GEN_2386 = mask_1[0] ? byte_512 : _GEN_1706; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2387 = mask_1[1] ? byte_513 : _GEN_1707; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2388 = mask_1[2] ? byte_514 : _GEN_1708; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2389 = mask_1[3] ? byte_515 : _GEN_1709; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2390 = _GEN_8842 == 8'h2a ? _GEN_2386 : _GEN_1706; // @[executor.scala 473:84]
  wire [7:0] _GEN_2391 = _GEN_8842 == 8'h2a ? _GEN_2387 : _GEN_1707; // @[executor.scala 473:84]
  wire [7:0] _GEN_2392 = _GEN_8842 == 8'h2a ? _GEN_2388 : _GEN_1708; // @[executor.scala 473:84]
  wire [7:0] _GEN_2393 = _GEN_8842 == 8'h2a ? _GEN_2389 : _GEN_1709; // @[executor.scala 473:84]
  wire [7:0] _GEN_2394 = mask_1[0] ? byte_512 : _GEN_1710; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2395 = mask_1[1] ? byte_513 : _GEN_1711; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2396 = mask_1[2] ? byte_514 : _GEN_1712; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2397 = mask_1[3] ? byte_515 : _GEN_1713; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2398 = _GEN_8842 == 8'h2b ? _GEN_2394 : _GEN_1710; // @[executor.scala 473:84]
  wire [7:0] _GEN_2399 = _GEN_8842 == 8'h2b ? _GEN_2395 : _GEN_1711; // @[executor.scala 473:84]
  wire [7:0] _GEN_2400 = _GEN_8842 == 8'h2b ? _GEN_2396 : _GEN_1712; // @[executor.scala 473:84]
  wire [7:0] _GEN_2401 = _GEN_8842 == 8'h2b ? _GEN_2397 : _GEN_1713; // @[executor.scala 473:84]
  wire [7:0] _GEN_2402 = mask_1[0] ? byte_512 : _GEN_1714; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2403 = mask_1[1] ? byte_513 : _GEN_1715; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2404 = mask_1[2] ? byte_514 : _GEN_1716; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2405 = mask_1[3] ? byte_515 : _GEN_1717; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2406 = _GEN_8842 == 8'h2c ? _GEN_2402 : _GEN_1714; // @[executor.scala 473:84]
  wire [7:0] _GEN_2407 = _GEN_8842 == 8'h2c ? _GEN_2403 : _GEN_1715; // @[executor.scala 473:84]
  wire [7:0] _GEN_2408 = _GEN_8842 == 8'h2c ? _GEN_2404 : _GEN_1716; // @[executor.scala 473:84]
  wire [7:0] _GEN_2409 = _GEN_8842 == 8'h2c ? _GEN_2405 : _GEN_1717; // @[executor.scala 473:84]
  wire [7:0] _GEN_2410 = mask_1[0] ? byte_512 : _GEN_1718; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2411 = mask_1[1] ? byte_513 : _GEN_1719; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2412 = mask_1[2] ? byte_514 : _GEN_1720; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2413 = mask_1[3] ? byte_515 : _GEN_1721; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2414 = _GEN_8842 == 8'h2d ? _GEN_2410 : _GEN_1718; // @[executor.scala 473:84]
  wire [7:0] _GEN_2415 = _GEN_8842 == 8'h2d ? _GEN_2411 : _GEN_1719; // @[executor.scala 473:84]
  wire [7:0] _GEN_2416 = _GEN_8842 == 8'h2d ? _GEN_2412 : _GEN_1720; // @[executor.scala 473:84]
  wire [7:0] _GEN_2417 = _GEN_8842 == 8'h2d ? _GEN_2413 : _GEN_1721; // @[executor.scala 473:84]
  wire [7:0] _GEN_2418 = mask_1[0] ? byte_512 : _GEN_1722; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2419 = mask_1[1] ? byte_513 : _GEN_1723; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2420 = mask_1[2] ? byte_514 : _GEN_1724; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2421 = mask_1[3] ? byte_515 : _GEN_1725; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2422 = _GEN_8842 == 8'h2e ? _GEN_2418 : _GEN_1722; // @[executor.scala 473:84]
  wire [7:0] _GEN_2423 = _GEN_8842 == 8'h2e ? _GEN_2419 : _GEN_1723; // @[executor.scala 473:84]
  wire [7:0] _GEN_2424 = _GEN_8842 == 8'h2e ? _GEN_2420 : _GEN_1724; // @[executor.scala 473:84]
  wire [7:0] _GEN_2425 = _GEN_8842 == 8'h2e ? _GEN_2421 : _GEN_1725; // @[executor.scala 473:84]
  wire [7:0] _GEN_2426 = mask_1[0] ? byte_512 : _GEN_1726; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2427 = mask_1[1] ? byte_513 : _GEN_1727; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2428 = mask_1[2] ? byte_514 : _GEN_1728; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2429 = mask_1[3] ? byte_515 : _GEN_1729; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2430 = _GEN_8842 == 8'h2f ? _GEN_2426 : _GEN_1726; // @[executor.scala 473:84]
  wire [7:0] _GEN_2431 = _GEN_8842 == 8'h2f ? _GEN_2427 : _GEN_1727; // @[executor.scala 473:84]
  wire [7:0] _GEN_2432 = _GEN_8842 == 8'h2f ? _GEN_2428 : _GEN_1728; // @[executor.scala 473:84]
  wire [7:0] _GEN_2433 = _GEN_8842 == 8'h2f ? _GEN_2429 : _GEN_1729; // @[executor.scala 473:84]
  wire [7:0] _GEN_2434 = mask_1[0] ? byte_512 : _GEN_1730; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2435 = mask_1[1] ? byte_513 : _GEN_1731; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2436 = mask_1[2] ? byte_514 : _GEN_1732; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2437 = mask_1[3] ? byte_515 : _GEN_1733; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2438 = _GEN_8842 == 8'h30 ? _GEN_2434 : _GEN_1730; // @[executor.scala 473:84]
  wire [7:0] _GEN_2439 = _GEN_8842 == 8'h30 ? _GEN_2435 : _GEN_1731; // @[executor.scala 473:84]
  wire [7:0] _GEN_2440 = _GEN_8842 == 8'h30 ? _GEN_2436 : _GEN_1732; // @[executor.scala 473:84]
  wire [7:0] _GEN_2441 = _GEN_8842 == 8'h30 ? _GEN_2437 : _GEN_1733; // @[executor.scala 473:84]
  wire [7:0] _GEN_2442 = mask_1[0] ? byte_512 : _GEN_1734; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2443 = mask_1[1] ? byte_513 : _GEN_1735; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2444 = mask_1[2] ? byte_514 : _GEN_1736; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2445 = mask_1[3] ? byte_515 : _GEN_1737; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2446 = _GEN_8842 == 8'h31 ? _GEN_2442 : _GEN_1734; // @[executor.scala 473:84]
  wire [7:0] _GEN_2447 = _GEN_8842 == 8'h31 ? _GEN_2443 : _GEN_1735; // @[executor.scala 473:84]
  wire [7:0] _GEN_2448 = _GEN_8842 == 8'h31 ? _GEN_2444 : _GEN_1736; // @[executor.scala 473:84]
  wire [7:0] _GEN_2449 = _GEN_8842 == 8'h31 ? _GEN_2445 : _GEN_1737; // @[executor.scala 473:84]
  wire [7:0] _GEN_2450 = mask_1[0] ? byte_512 : _GEN_1738; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2451 = mask_1[1] ? byte_513 : _GEN_1739; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2452 = mask_1[2] ? byte_514 : _GEN_1740; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2453 = mask_1[3] ? byte_515 : _GEN_1741; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2454 = _GEN_8842 == 8'h32 ? _GEN_2450 : _GEN_1738; // @[executor.scala 473:84]
  wire [7:0] _GEN_2455 = _GEN_8842 == 8'h32 ? _GEN_2451 : _GEN_1739; // @[executor.scala 473:84]
  wire [7:0] _GEN_2456 = _GEN_8842 == 8'h32 ? _GEN_2452 : _GEN_1740; // @[executor.scala 473:84]
  wire [7:0] _GEN_2457 = _GEN_8842 == 8'h32 ? _GEN_2453 : _GEN_1741; // @[executor.scala 473:84]
  wire [7:0] _GEN_2458 = mask_1[0] ? byte_512 : _GEN_1742; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2459 = mask_1[1] ? byte_513 : _GEN_1743; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2460 = mask_1[2] ? byte_514 : _GEN_1744; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2461 = mask_1[3] ? byte_515 : _GEN_1745; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2462 = _GEN_8842 == 8'h33 ? _GEN_2458 : _GEN_1742; // @[executor.scala 473:84]
  wire [7:0] _GEN_2463 = _GEN_8842 == 8'h33 ? _GEN_2459 : _GEN_1743; // @[executor.scala 473:84]
  wire [7:0] _GEN_2464 = _GEN_8842 == 8'h33 ? _GEN_2460 : _GEN_1744; // @[executor.scala 473:84]
  wire [7:0] _GEN_2465 = _GEN_8842 == 8'h33 ? _GEN_2461 : _GEN_1745; // @[executor.scala 473:84]
  wire [7:0] _GEN_2466 = mask_1[0] ? byte_512 : _GEN_1746; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2467 = mask_1[1] ? byte_513 : _GEN_1747; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2468 = mask_1[2] ? byte_514 : _GEN_1748; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2469 = mask_1[3] ? byte_515 : _GEN_1749; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2470 = _GEN_8842 == 8'h34 ? _GEN_2466 : _GEN_1746; // @[executor.scala 473:84]
  wire [7:0] _GEN_2471 = _GEN_8842 == 8'h34 ? _GEN_2467 : _GEN_1747; // @[executor.scala 473:84]
  wire [7:0] _GEN_2472 = _GEN_8842 == 8'h34 ? _GEN_2468 : _GEN_1748; // @[executor.scala 473:84]
  wire [7:0] _GEN_2473 = _GEN_8842 == 8'h34 ? _GEN_2469 : _GEN_1749; // @[executor.scala 473:84]
  wire [7:0] _GEN_2474 = mask_1[0] ? byte_512 : _GEN_1750; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2475 = mask_1[1] ? byte_513 : _GEN_1751; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2476 = mask_1[2] ? byte_514 : _GEN_1752; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2477 = mask_1[3] ? byte_515 : _GEN_1753; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2478 = _GEN_8842 == 8'h35 ? _GEN_2474 : _GEN_1750; // @[executor.scala 473:84]
  wire [7:0] _GEN_2479 = _GEN_8842 == 8'h35 ? _GEN_2475 : _GEN_1751; // @[executor.scala 473:84]
  wire [7:0] _GEN_2480 = _GEN_8842 == 8'h35 ? _GEN_2476 : _GEN_1752; // @[executor.scala 473:84]
  wire [7:0] _GEN_2481 = _GEN_8842 == 8'h35 ? _GEN_2477 : _GEN_1753; // @[executor.scala 473:84]
  wire [7:0] _GEN_2482 = mask_1[0] ? byte_512 : _GEN_1754; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2483 = mask_1[1] ? byte_513 : _GEN_1755; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2484 = mask_1[2] ? byte_514 : _GEN_1756; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2485 = mask_1[3] ? byte_515 : _GEN_1757; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2486 = _GEN_8842 == 8'h36 ? _GEN_2482 : _GEN_1754; // @[executor.scala 473:84]
  wire [7:0] _GEN_2487 = _GEN_8842 == 8'h36 ? _GEN_2483 : _GEN_1755; // @[executor.scala 473:84]
  wire [7:0] _GEN_2488 = _GEN_8842 == 8'h36 ? _GEN_2484 : _GEN_1756; // @[executor.scala 473:84]
  wire [7:0] _GEN_2489 = _GEN_8842 == 8'h36 ? _GEN_2485 : _GEN_1757; // @[executor.scala 473:84]
  wire [7:0] _GEN_2490 = mask_1[0] ? byte_512 : _GEN_1758; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2491 = mask_1[1] ? byte_513 : _GEN_1759; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2492 = mask_1[2] ? byte_514 : _GEN_1760; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2493 = mask_1[3] ? byte_515 : _GEN_1761; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2494 = _GEN_8842 == 8'h37 ? _GEN_2490 : _GEN_1758; // @[executor.scala 473:84]
  wire [7:0] _GEN_2495 = _GEN_8842 == 8'h37 ? _GEN_2491 : _GEN_1759; // @[executor.scala 473:84]
  wire [7:0] _GEN_2496 = _GEN_8842 == 8'h37 ? _GEN_2492 : _GEN_1760; // @[executor.scala 473:84]
  wire [7:0] _GEN_2497 = _GEN_8842 == 8'h37 ? _GEN_2493 : _GEN_1761; // @[executor.scala 473:84]
  wire [7:0] _GEN_2498 = mask_1[0] ? byte_512 : _GEN_1762; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2499 = mask_1[1] ? byte_513 : _GEN_1763; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2500 = mask_1[2] ? byte_514 : _GEN_1764; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2501 = mask_1[3] ? byte_515 : _GEN_1765; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2502 = _GEN_8842 == 8'h38 ? _GEN_2498 : _GEN_1762; // @[executor.scala 473:84]
  wire [7:0] _GEN_2503 = _GEN_8842 == 8'h38 ? _GEN_2499 : _GEN_1763; // @[executor.scala 473:84]
  wire [7:0] _GEN_2504 = _GEN_8842 == 8'h38 ? _GEN_2500 : _GEN_1764; // @[executor.scala 473:84]
  wire [7:0] _GEN_2505 = _GEN_8842 == 8'h38 ? _GEN_2501 : _GEN_1765; // @[executor.scala 473:84]
  wire [7:0] _GEN_2506 = mask_1[0] ? byte_512 : _GEN_1766; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2507 = mask_1[1] ? byte_513 : _GEN_1767; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2508 = mask_1[2] ? byte_514 : _GEN_1768; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2509 = mask_1[3] ? byte_515 : _GEN_1769; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2510 = _GEN_8842 == 8'h39 ? _GEN_2506 : _GEN_1766; // @[executor.scala 473:84]
  wire [7:0] _GEN_2511 = _GEN_8842 == 8'h39 ? _GEN_2507 : _GEN_1767; // @[executor.scala 473:84]
  wire [7:0] _GEN_2512 = _GEN_8842 == 8'h39 ? _GEN_2508 : _GEN_1768; // @[executor.scala 473:84]
  wire [7:0] _GEN_2513 = _GEN_8842 == 8'h39 ? _GEN_2509 : _GEN_1769; // @[executor.scala 473:84]
  wire [7:0] _GEN_2514 = mask_1[0] ? byte_512 : _GEN_1770; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2515 = mask_1[1] ? byte_513 : _GEN_1771; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2516 = mask_1[2] ? byte_514 : _GEN_1772; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2517 = mask_1[3] ? byte_515 : _GEN_1773; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2518 = _GEN_8842 == 8'h3a ? _GEN_2514 : _GEN_1770; // @[executor.scala 473:84]
  wire [7:0] _GEN_2519 = _GEN_8842 == 8'h3a ? _GEN_2515 : _GEN_1771; // @[executor.scala 473:84]
  wire [7:0] _GEN_2520 = _GEN_8842 == 8'h3a ? _GEN_2516 : _GEN_1772; // @[executor.scala 473:84]
  wire [7:0] _GEN_2521 = _GEN_8842 == 8'h3a ? _GEN_2517 : _GEN_1773; // @[executor.scala 473:84]
  wire [7:0] _GEN_2522 = mask_1[0] ? byte_512 : _GEN_1774; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2523 = mask_1[1] ? byte_513 : _GEN_1775; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2524 = mask_1[2] ? byte_514 : _GEN_1776; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2525 = mask_1[3] ? byte_515 : _GEN_1777; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2526 = _GEN_8842 == 8'h3b ? _GEN_2522 : _GEN_1774; // @[executor.scala 473:84]
  wire [7:0] _GEN_2527 = _GEN_8842 == 8'h3b ? _GEN_2523 : _GEN_1775; // @[executor.scala 473:84]
  wire [7:0] _GEN_2528 = _GEN_8842 == 8'h3b ? _GEN_2524 : _GEN_1776; // @[executor.scala 473:84]
  wire [7:0] _GEN_2529 = _GEN_8842 == 8'h3b ? _GEN_2525 : _GEN_1777; // @[executor.scala 473:84]
  wire [7:0] _GEN_2530 = mask_1[0] ? byte_512 : _GEN_1778; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2531 = mask_1[1] ? byte_513 : _GEN_1779; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2532 = mask_1[2] ? byte_514 : _GEN_1780; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2533 = mask_1[3] ? byte_515 : _GEN_1781; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2534 = _GEN_8842 == 8'h3c ? _GEN_2530 : _GEN_1778; // @[executor.scala 473:84]
  wire [7:0] _GEN_2535 = _GEN_8842 == 8'h3c ? _GEN_2531 : _GEN_1779; // @[executor.scala 473:84]
  wire [7:0] _GEN_2536 = _GEN_8842 == 8'h3c ? _GEN_2532 : _GEN_1780; // @[executor.scala 473:84]
  wire [7:0] _GEN_2537 = _GEN_8842 == 8'h3c ? _GEN_2533 : _GEN_1781; // @[executor.scala 473:84]
  wire [7:0] _GEN_2538 = mask_1[0] ? byte_512 : _GEN_1782; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2539 = mask_1[1] ? byte_513 : _GEN_1783; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2540 = mask_1[2] ? byte_514 : _GEN_1784; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2541 = mask_1[3] ? byte_515 : _GEN_1785; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2542 = _GEN_8842 == 8'h3d ? _GEN_2538 : _GEN_1782; // @[executor.scala 473:84]
  wire [7:0] _GEN_2543 = _GEN_8842 == 8'h3d ? _GEN_2539 : _GEN_1783; // @[executor.scala 473:84]
  wire [7:0] _GEN_2544 = _GEN_8842 == 8'h3d ? _GEN_2540 : _GEN_1784; // @[executor.scala 473:84]
  wire [7:0] _GEN_2545 = _GEN_8842 == 8'h3d ? _GEN_2541 : _GEN_1785; // @[executor.scala 473:84]
  wire [7:0] _GEN_2546 = mask_1[0] ? byte_512 : _GEN_1786; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2547 = mask_1[1] ? byte_513 : _GEN_1787; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2548 = mask_1[2] ? byte_514 : _GEN_1788; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2549 = mask_1[3] ? byte_515 : _GEN_1789; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2550 = _GEN_8842 == 8'h3e ? _GEN_2546 : _GEN_1786; // @[executor.scala 473:84]
  wire [7:0] _GEN_2551 = _GEN_8842 == 8'h3e ? _GEN_2547 : _GEN_1787; // @[executor.scala 473:84]
  wire [7:0] _GEN_2552 = _GEN_8842 == 8'h3e ? _GEN_2548 : _GEN_1788; // @[executor.scala 473:84]
  wire [7:0] _GEN_2553 = _GEN_8842 == 8'h3e ? _GEN_2549 : _GEN_1789; // @[executor.scala 473:84]
  wire [7:0] _GEN_2554 = mask_1[0] ? byte_512 : _GEN_1790; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2555 = mask_1[1] ? byte_513 : _GEN_1791; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2556 = mask_1[2] ? byte_514 : _GEN_1792; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2557 = mask_1[3] ? byte_515 : _GEN_1793; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2558 = _GEN_8842 == 8'h3f ? _GEN_2554 : _GEN_1790; // @[executor.scala 473:84]
  wire [7:0] _GEN_2559 = _GEN_8842 == 8'h3f ? _GEN_2555 : _GEN_1791; // @[executor.scala 473:84]
  wire [7:0] _GEN_2560 = _GEN_8842 == 8'h3f ? _GEN_2556 : _GEN_1792; // @[executor.scala 473:84]
  wire [7:0] _GEN_2561 = _GEN_8842 == 8'h3f ? _GEN_2557 : _GEN_1793; // @[executor.scala 473:84]
  wire [7:0] _GEN_2562 = mask_1[0] ? byte_512 : _GEN_1794; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2563 = mask_1[1] ? byte_513 : _GEN_1795; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2564 = mask_1[2] ? byte_514 : _GEN_1796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2565 = mask_1[3] ? byte_515 : _GEN_1797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2566 = _GEN_8842 == 8'h40 ? _GEN_2562 : _GEN_1794; // @[executor.scala 473:84]
  wire [7:0] _GEN_2567 = _GEN_8842 == 8'h40 ? _GEN_2563 : _GEN_1795; // @[executor.scala 473:84]
  wire [7:0] _GEN_2568 = _GEN_8842 == 8'h40 ? _GEN_2564 : _GEN_1796; // @[executor.scala 473:84]
  wire [7:0] _GEN_2569 = _GEN_8842 == 8'h40 ? _GEN_2565 : _GEN_1797; // @[executor.scala 473:84]
  wire [7:0] _GEN_2570 = mask_1[0] ? byte_512 : _GEN_1798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2571 = mask_1[1] ? byte_513 : _GEN_1799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2572 = mask_1[2] ? byte_514 : _GEN_1800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2573 = mask_1[3] ? byte_515 : _GEN_1801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2574 = _GEN_8842 == 8'h41 ? _GEN_2570 : _GEN_1798; // @[executor.scala 473:84]
  wire [7:0] _GEN_2575 = _GEN_8842 == 8'h41 ? _GEN_2571 : _GEN_1799; // @[executor.scala 473:84]
  wire [7:0] _GEN_2576 = _GEN_8842 == 8'h41 ? _GEN_2572 : _GEN_1800; // @[executor.scala 473:84]
  wire [7:0] _GEN_2577 = _GEN_8842 == 8'h41 ? _GEN_2573 : _GEN_1801; // @[executor.scala 473:84]
  wire [7:0] _GEN_2578 = mask_1[0] ? byte_512 : _GEN_1802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2579 = mask_1[1] ? byte_513 : _GEN_1803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2580 = mask_1[2] ? byte_514 : _GEN_1804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2581 = mask_1[3] ? byte_515 : _GEN_1805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2582 = _GEN_8842 == 8'h42 ? _GEN_2578 : _GEN_1802; // @[executor.scala 473:84]
  wire [7:0] _GEN_2583 = _GEN_8842 == 8'h42 ? _GEN_2579 : _GEN_1803; // @[executor.scala 473:84]
  wire [7:0] _GEN_2584 = _GEN_8842 == 8'h42 ? _GEN_2580 : _GEN_1804; // @[executor.scala 473:84]
  wire [7:0] _GEN_2585 = _GEN_8842 == 8'h42 ? _GEN_2581 : _GEN_1805; // @[executor.scala 473:84]
  wire [7:0] _GEN_2586 = mask_1[0] ? byte_512 : _GEN_1806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2587 = mask_1[1] ? byte_513 : _GEN_1807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2588 = mask_1[2] ? byte_514 : _GEN_1808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2589 = mask_1[3] ? byte_515 : _GEN_1809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2590 = _GEN_8842 == 8'h43 ? _GEN_2586 : _GEN_1806; // @[executor.scala 473:84]
  wire [7:0] _GEN_2591 = _GEN_8842 == 8'h43 ? _GEN_2587 : _GEN_1807; // @[executor.scala 473:84]
  wire [7:0] _GEN_2592 = _GEN_8842 == 8'h43 ? _GEN_2588 : _GEN_1808; // @[executor.scala 473:84]
  wire [7:0] _GEN_2593 = _GEN_8842 == 8'h43 ? _GEN_2589 : _GEN_1809; // @[executor.scala 473:84]
  wire [7:0] _GEN_2594 = mask_1[0] ? byte_512 : _GEN_1810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2595 = mask_1[1] ? byte_513 : _GEN_1811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2596 = mask_1[2] ? byte_514 : _GEN_1812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2597 = mask_1[3] ? byte_515 : _GEN_1813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2598 = _GEN_8842 == 8'h44 ? _GEN_2594 : _GEN_1810; // @[executor.scala 473:84]
  wire [7:0] _GEN_2599 = _GEN_8842 == 8'h44 ? _GEN_2595 : _GEN_1811; // @[executor.scala 473:84]
  wire [7:0] _GEN_2600 = _GEN_8842 == 8'h44 ? _GEN_2596 : _GEN_1812; // @[executor.scala 473:84]
  wire [7:0] _GEN_2601 = _GEN_8842 == 8'h44 ? _GEN_2597 : _GEN_1813; // @[executor.scala 473:84]
  wire [7:0] _GEN_2602 = mask_1[0] ? byte_512 : _GEN_1814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2603 = mask_1[1] ? byte_513 : _GEN_1815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2604 = mask_1[2] ? byte_514 : _GEN_1816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2605 = mask_1[3] ? byte_515 : _GEN_1817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2606 = _GEN_8842 == 8'h45 ? _GEN_2602 : _GEN_1814; // @[executor.scala 473:84]
  wire [7:0] _GEN_2607 = _GEN_8842 == 8'h45 ? _GEN_2603 : _GEN_1815; // @[executor.scala 473:84]
  wire [7:0] _GEN_2608 = _GEN_8842 == 8'h45 ? _GEN_2604 : _GEN_1816; // @[executor.scala 473:84]
  wire [7:0] _GEN_2609 = _GEN_8842 == 8'h45 ? _GEN_2605 : _GEN_1817; // @[executor.scala 473:84]
  wire [7:0] _GEN_2610 = mask_1[0] ? byte_512 : _GEN_1818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2611 = mask_1[1] ? byte_513 : _GEN_1819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2612 = mask_1[2] ? byte_514 : _GEN_1820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2613 = mask_1[3] ? byte_515 : _GEN_1821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2614 = _GEN_8842 == 8'h46 ? _GEN_2610 : _GEN_1818; // @[executor.scala 473:84]
  wire [7:0] _GEN_2615 = _GEN_8842 == 8'h46 ? _GEN_2611 : _GEN_1819; // @[executor.scala 473:84]
  wire [7:0] _GEN_2616 = _GEN_8842 == 8'h46 ? _GEN_2612 : _GEN_1820; // @[executor.scala 473:84]
  wire [7:0] _GEN_2617 = _GEN_8842 == 8'h46 ? _GEN_2613 : _GEN_1821; // @[executor.scala 473:84]
  wire [7:0] _GEN_2618 = mask_1[0] ? byte_512 : _GEN_1822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2619 = mask_1[1] ? byte_513 : _GEN_1823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2620 = mask_1[2] ? byte_514 : _GEN_1824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2621 = mask_1[3] ? byte_515 : _GEN_1825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2622 = _GEN_8842 == 8'h47 ? _GEN_2618 : _GEN_1822; // @[executor.scala 473:84]
  wire [7:0] _GEN_2623 = _GEN_8842 == 8'h47 ? _GEN_2619 : _GEN_1823; // @[executor.scala 473:84]
  wire [7:0] _GEN_2624 = _GEN_8842 == 8'h47 ? _GEN_2620 : _GEN_1824; // @[executor.scala 473:84]
  wire [7:0] _GEN_2625 = _GEN_8842 == 8'h47 ? _GEN_2621 : _GEN_1825; // @[executor.scala 473:84]
  wire [7:0] _GEN_2626 = mask_1[0] ? byte_512 : _GEN_1826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2627 = mask_1[1] ? byte_513 : _GEN_1827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2628 = mask_1[2] ? byte_514 : _GEN_1828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2629 = mask_1[3] ? byte_515 : _GEN_1829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2630 = _GEN_8842 == 8'h48 ? _GEN_2626 : _GEN_1826; // @[executor.scala 473:84]
  wire [7:0] _GEN_2631 = _GEN_8842 == 8'h48 ? _GEN_2627 : _GEN_1827; // @[executor.scala 473:84]
  wire [7:0] _GEN_2632 = _GEN_8842 == 8'h48 ? _GEN_2628 : _GEN_1828; // @[executor.scala 473:84]
  wire [7:0] _GEN_2633 = _GEN_8842 == 8'h48 ? _GEN_2629 : _GEN_1829; // @[executor.scala 473:84]
  wire [7:0] _GEN_2634 = mask_1[0] ? byte_512 : _GEN_1830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2635 = mask_1[1] ? byte_513 : _GEN_1831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2636 = mask_1[2] ? byte_514 : _GEN_1832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2637 = mask_1[3] ? byte_515 : _GEN_1833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2638 = _GEN_8842 == 8'h49 ? _GEN_2634 : _GEN_1830; // @[executor.scala 473:84]
  wire [7:0] _GEN_2639 = _GEN_8842 == 8'h49 ? _GEN_2635 : _GEN_1831; // @[executor.scala 473:84]
  wire [7:0] _GEN_2640 = _GEN_8842 == 8'h49 ? _GEN_2636 : _GEN_1832; // @[executor.scala 473:84]
  wire [7:0] _GEN_2641 = _GEN_8842 == 8'h49 ? _GEN_2637 : _GEN_1833; // @[executor.scala 473:84]
  wire [7:0] _GEN_2642 = mask_1[0] ? byte_512 : _GEN_1834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2643 = mask_1[1] ? byte_513 : _GEN_1835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2644 = mask_1[2] ? byte_514 : _GEN_1836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2645 = mask_1[3] ? byte_515 : _GEN_1837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2646 = _GEN_8842 == 8'h4a ? _GEN_2642 : _GEN_1834; // @[executor.scala 473:84]
  wire [7:0] _GEN_2647 = _GEN_8842 == 8'h4a ? _GEN_2643 : _GEN_1835; // @[executor.scala 473:84]
  wire [7:0] _GEN_2648 = _GEN_8842 == 8'h4a ? _GEN_2644 : _GEN_1836; // @[executor.scala 473:84]
  wire [7:0] _GEN_2649 = _GEN_8842 == 8'h4a ? _GEN_2645 : _GEN_1837; // @[executor.scala 473:84]
  wire [7:0] _GEN_2650 = mask_1[0] ? byte_512 : _GEN_1838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2651 = mask_1[1] ? byte_513 : _GEN_1839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2652 = mask_1[2] ? byte_514 : _GEN_1840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2653 = mask_1[3] ? byte_515 : _GEN_1841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2654 = _GEN_8842 == 8'h4b ? _GEN_2650 : _GEN_1838; // @[executor.scala 473:84]
  wire [7:0] _GEN_2655 = _GEN_8842 == 8'h4b ? _GEN_2651 : _GEN_1839; // @[executor.scala 473:84]
  wire [7:0] _GEN_2656 = _GEN_8842 == 8'h4b ? _GEN_2652 : _GEN_1840; // @[executor.scala 473:84]
  wire [7:0] _GEN_2657 = _GEN_8842 == 8'h4b ? _GEN_2653 : _GEN_1841; // @[executor.scala 473:84]
  wire [7:0] _GEN_2658 = mask_1[0] ? byte_512 : _GEN_1842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2659 = mask_1[1] ? byte_513 : _GEN_1843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2660 = mask_1[2] ? byte_514 : _GEN_1844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2661 = mask_1[3] ? byte_515 : _GEN_1845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2662 = _GEN_8842 == 8'h4c ? _GEN_2658 : _GEN_1842; // @[executor.scala 473:84]
  wire [7:0] _GEN_2663 = _GEN_8842 == 8'h4c ? _GEN_2659 : _GEN_1843; // @[executor.scala 473:84]
  wire [7:0] _GEN_2664 = _GEN_8842 == 8'h4c ? _GEN_2660 : _GEN_1844; // @[executor.scala 473:84]
  wire [7:0] _GEN_2665 = _GEN_8842 == 8'h4c ? _GEN_2661 : _GEN_1845; // @[executor.scala 473:84]
  wire [7:0] _GEN_2666 = mask_1[0] ? byte_512 : _GEN_1846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2667 = mask_1[1] ? byte_513 : _GEN_1847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2668 = mask_1[2] ? byte_514 : _GEN_1848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2669 = mask_1[3] ? byte_515 : _GEN_1849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2670 = _GEN_8842 == 8'h4d ? _GEN_2666 : _GEN_1846; // @[executor.scala 473:84]
  wire [7:0] _GEN_2671 = _GEN_8842 == 8'h4d ? _GEN_2667 : _GEN_1847; // @[executor.scala 473:84]
  wire [7:0] _GEN_2672 = _GEN_8842 == 8'h4d ? _GEN_2668 : _GEN_1848; // @[executor.scala 473:84]
  wire [7:0] _GEN_2673 = _GEN_8842 == 8'h4d ? _GEN_2669 : _GEN_1849; // @[executor.scala 473:84]
  wire [7:0] _GEN_2674 = mask_1[0] ? byte_512 : _GEN_1850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2675 = mask_1[1] ? byte_513 : _GEN_1851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2676 = mask_1[2] ? byte_514 : _GEN_1852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2677 = mask_1[3] ? byte_515 : _GEN_1853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2678 = _GEN_8842 == 8'h4e ? _GEN_2674 : _GEN_1850; // @[executor.scala 473:84]
  wire [7:0] _GEN_2679 = _GEN_8842 == 8'h4e ? _GEN_2675 : _GEN_1851; // @[executor.scala 473:84]
  wire [7:0] _GEN_2680 = _GEN_8842 == 8'h4e ? _GEN_2676 : _GEN_1852; // @[executor.scala 473:84]
  wire [7:0] _GEN_2681 = _GEN_8842 == 8'h4e ? _GEN_2677 : _GEN_1853; // @[executor.scala 473:84]
  wire [7:0] _GEN_2682 = mask_1[0] ? byte_512 : _GEN_1854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2683 = mask_1[1] ? byte_513 : _GEN_1855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2684 = mask_1[2] ? byte_514 : _GEN_1856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2685 = mask_1[3] ? byte_515 : _GEN_1857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2686 = _GEN_8842 == 8'h4f ? _GEN_2682 : _GEN_1854; // @[executor.scala 473:84]
  wire [7:0] _GEN_2687 = _GEN_8842 == 8'h4f ? _GEN_2683 : _GEN_1855; // @[executor.scala 473:84]
  wire [7:0] _GEN_2688 = _GEN_8842 == 8'h4f ? _GEN_2684 : _GEN_1856; // @[executor.scala 473:84]
  wire [7:0] _GEN_2689 = _GEN_8842 == 8'h4f ? _GEN_2685 : _GEN_1857; // @[executor.scala 473:84]
  wire [7:0] _GEN_2690 = mask_1[0] ? byte_512 : _GEN_1858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2691 = mask_1[1] ? byte_513 : _GEN_1859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2692 = mask_1[2] ? byte_514 : _GEN_1860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2693 = mask_1[3] ? byte_515 : _GEN_1861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2694 = _GEN_8842 == 8'h50 ? _GEN_2690 : _GEN_1858; // @[executor.scala 473:84]
  wire [7:0] _GEN_2695 = _GEN_8842 == 8'h50 ? _GEN_2691 : _GEN_1859; // @[executor.scala 473:84]
  wire [7:0] _GEN_2696 = _GEN_8842 == 8'h50 ? _GEN_2692 : _GEN_1860; // @[executor.scala 473:84]
  wire [7:0] _GEN_2697 = _GEN_8842 == 8'h50 ? _GEN_2693 : _GEN_1861; // @[executor.scala 473:84]
  wire [7:0] _GEN_2698 = mask_1[0] ? byte_512 : _GEN_1862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2699 = mask_1[1] ? byte_513 : _GEN_1863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2700 = mask_1[2] ? byte_514 : _GEN_1864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2701 = mask_1[3] ? byte_515 : _GEN_1865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2702 = _GEN_8842 == 8'h51 ? _GEN_2698 : _GEN_1862; // @[executor.scala 473:84]
  wire [7:0] _GEN_2703 = _GEN_8842 == 8'h51 ? _GEN_2699 : _GEN_1863; // @[executor.scala 473:84]
  wire [7:0] _GEN_2704 = _GEN_8842 == 8'h51 ? _GEN_2700 : _GEN_1864; // @[executor.scala 473:84]
  wire [7:0] _GEN_2705 = _GEN_8842 == 8'h51 ? _GEN_2701 : _GEN_1865; // @[executor.scala 473:84]
  wire [7:0] _GEN_2706 = mask_1[0] ? byte_512 : _GEN_1866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2707 = mask_1[1] ? byte_513 : _GEN_1867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2708 = mask_1[2] ? byte_514 : _GEN_1868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2709 = mask_1[3] ? byte_515 : _GEN_1869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2710 = _GEN_8842 == 8'h52 ? _GEN_2706 : _GEN_1866; // @[executor.scala 473:84]
  wire [7:0] _GEN_2711 = _GEN_8842 == 8'h52 ? _GEN_2707 : _GEN_1867; // @[executor.scala 473:84]
  wire [7:0] _GEN_2712 = _GEN_8842 == 8'h52 ? _GEN_2708 : _GEN_1868; // @[executor.scala 473:84]
  wire [7:0] _GEN_2713 = _GEN_8842 == 8'h52 ? _GEN_2709 : _GEN_1869; // @[executor.scala 473:84]
  wire [7:0] _GEN_2714 = mask_1[0] ? byte_512 : _GEN_1870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2715 = mask_1[1] ? byte_513 : _GEN_1871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2716 = mask_1[2] ? byte_514 : _GEN_1872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2717 = mask_1[3] ? byte_515 : _GEN_1873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2718 = _GEN_8842 == 8'h53 ? _GEN_2714 : _GEN_1870; // @[executor.scala 473:84]
  wire [7:0] _GEN_2719 = _GEN_8842 == 8'h53 ? _GEN_2715 : _GEN_1871; // @[executor.scala 473:84]
  wire [7:0] _GEN_2720 = _GEN_8842 == 8'h53 ? _GEN_2716 : _GEN_1872; // @[executor.scala 473:84]
  wire [7:0] _GEN_2721 = _GEN_8842 == 8'h53 ? _GEN_2717 : _GEN_1873; // @[executor.scala 473:84]
  wire [7:0] _GEN_2722 = mask_1[0] ? byte_512 : _GEN_1874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2723 = mask_1[1] ? byte_513 : _GEN_1875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2724 = mask_1[2] ? byte_514 : _GEN_1876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2725 = mask_1[3] ? byte_515 : _GEN_1877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2726 = _GEN_8842 == 8'h54 ? _GEN_2722 : _GEN_1874; // @[executor.scala 473:84]
  wire [7:0] _GEN_2727 = _GEN_8842 == 8'h54 ? _GEN_2723 : _GEN_1875; // @[executor.scala 473:84]
  wire [7:0] _GEN_2728 = _GEN_8842 == 8'h54 ? _GEN_2724 : _GEN_1876; // @[executor.scala 473:84]
  wire [7:0] _GEN_2729 = _GEN_8842 == 8'h54 ? _GEN_2725 : _GEN_1877; // @[executor.scala 473:84]
  wire [7:0] _GEN_2730 = mask_1[0] ? byte_512 : _GEN_1878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2731 = mask_1[1] ? byte_513 : _GEN_1879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2732 = mask_1[2] ? byte_514 : _GEN_1880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2733 = mask_1[3] ? byte_515 : _GEN_1881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2734 = _GEN_8842 == 8'h55 ? _GEN_2730 : _GEN_1878; // @[executor.scala 473:84]
  wire [7:0] _GEN_2735 = _GEN_8842 == 8'h55 ? _GEN_2731 : _GEN_1879; // @[executor.scala 473:84]
  wire [7:0] _GEN_2736 = _GEN_8842 == 8'h55 ? _GEN_2732 : _GEN_1880; // @[executor.scala 473:84]
  wire [7:0] _GEN_2737 = _GEN_8842 == 8'h55 ? _GEN_2733 : _GEN_1881; // @[executor.scala 473:84]
  wire [7:0] _GEN_2738 = mask_1[0] ? byte_512 : _GEN_1882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2739 = mask_1[1] ? byte_513 : _GEN_1883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2740 = mask_1[2] ? byte_514 : _GEN_1884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2741 = mask_1[3] ? byte_515 : _GEN_1885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2742 = _GEN_8842 == 8'h56 ? _GEN_2738 : _GEN_1882; // @[executor.scala 473:84]
  wire [7:0] _GEN_2743 = _GEN_8842 == 8'h56 ? _GEN_2739 : _GEN_1883; // @[executor.scala 473:84]
  wire [7:0] _GEN_2744 = _GEN_8842 == 8'h56 ? _GEN_2740 : _GEN_1884; // @[executor.scala 473:84]
  wire [7:0] _GEN_2745 = _GEN_8842 == 8'h56 ? _GEN_2741 : _GEN_1885; // @[executor.scala 473:84]
  wire [7:0] _GEN_2746 = mask_1[0] ? byte_512 : _GEN_1886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2747 = mask_1[1] ? byte_513 : _GEN_1887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2748 = mask_1[2] ? byte_514 : _GEN_1888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2749 = mask_1[3] ? byte_515 : _GEN_1889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2750 = _GEN_8842 == 8'h57 ? _GEN_2746 : _GEN_1886; // @[executor.scala 473:84]
  wire [7:0] _GEN_2751 = _GEN_8842 == 8'h57 ? _GEN_2747 : _GEN_1887; // @[executor.scala 473:84]
  wire [7:0] _GEN_2752 = _GEN_8842 == 8'h57 ? _GEN_2748 : _GEN_1888; // @[executor.scala 473:84]
  wire [7:0] _GEN_2753 = _GEN_8842 == 8'h57 ? _GEN_2749 : _GEN_1889; // @[executor.scala 473:84]
  wire [7:0] _GEN_2754 = mask_1[0] ? byte_512 : _GEN_1890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2755 = mask_1[1] ? byte_513 : _GEN_1891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2756 = mask_1[2] ? byte_514 : _GEN_1892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2757 = mask_1[3] ? byte_515 : _GEN_1893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2758 = _GEN_8842 == 8'h58 ? _GEN_2754 : _GEN_1890; // @[executor.scala 473:84]
  wire [7:0] _GEN_2759 = _GEN_8842 == 8'h58 ? _GEN_2755 : _GEN_1891; // @[executor.scala 473:84]
  wire [7:0] _GEN_2760 = _GEN_8842 == 8'h58 ? _GEN_2756 : _GEN_1892; // @[executor.scala 473:84]
  wire [7:0] _GEN_2761 = _GEN_8842 == 8'h58 ? _GEN_2757 : _GEN_1893; // @[executor.scala 473:84]
  wire [7:0] _GEN_2762 = mask_1[0] ? byte_512 : _GEN_1894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2763 = mask_1[1] ? byte_513 : _GEN_1895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2764 = mask_1[2] ? byte_514 : _GEN_1896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2765 = mask_1[3] ? byte_515 : _GEN_1897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2766 = _GEN_8842 == 8'h59 ? _GEN_2762 : _GEN_1894; // @[executor.scala 473:84]
  wire [7:0] _GEN_2767 = _GEN_8842 == 8'h59 ? _GEN_2763 : _GEN_1895; // @[executor.scala 473:84]
  wire [7:0] _GEN_2768 = _GEN_8842 == 8'h59 ? _GEN_2764 : _GEN_1896; // @[executor.scala 473:84]
  wire [7:0] _GEN_2769 = _GEN_8842 == 8'h59 ? _GEN_2765 : _GEN_1897; // @[executor.scala 473:84]
  wire [7:0] _GEN_2770 = mask_1[0] ? byte_512 : _GEN_1898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2771 = mask_1[1] ? byte_513 : _GEN_1899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2772 = mask_1[2] ? byte_514 : _GEN_1900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2773 = mask_1[3] ? byte_515 : _GEN_1901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2774 = _GEN_8842 == 8'h5a ? _GEN_2770 : _GEN_1898; // @[executor.scala 473:84]
  wire [7:0] _GEN_2775 = _GEN_8842 == 8'h5a ? _GEN_2771 : _GEN_1899; // @[executor.scala 473:84]
  wire [7:0] _GEN_2776 = _GEN_8842 == 8'h5a ? _GEN_2772 : _GEN_1900; // @[executor.scala 473:84]
  wire [7:0] _GEN_2777 = _GEN_8842 == 8'h5a ? _GEN_2773 : _GEN_1901; // @[executor.scala 473:84]
  wire [7:0] _GEN_2778 = mask_1[0] ? byte_512 : _GEN_1902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2779 = mask_1[1] ? byte_513 : _GEN_1903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2780 = mask_1[2] ? byte_514 : _GEN_1904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2781 = mask_1[3] ? byte_515 : _GEN_1905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2782 = _GEN_8842 == 8'h5b ? _GEN_2778 : _GEN_1902; // @[executor.scala 473:84]
  wire [7:0] _GEN_2783 = _GEN_8842 == 8'h5b ? _GEN_2779 : _GEN_1903; // @[executor.scala 473:84]
  wire [7:0] _GEN_2784 = _GEN_8842 == 8'h5b ? _GEN_2780 : _GEN_1904; // @[executor.scala 473:84]
  wire [7:0] _GEN_2785 = _GEN_8842 == 8'h5b ? _GEN_2781 : _GEN_1905; // @[executor.scala 473:84]
  wire [7:0] _GEN_2786 = mask_1[0] ? byte_512 : _GEN_1906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2787 = mask_1[1] ? byte_513 : _GEN_1907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2788 = mask_1[2] ? byte_514 : _GEN_1908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2789 = mask_1[3] ? byte_515 : _GEN_1909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2790 = _GEN_8842 == 8'h5c ? _GEN_2786 : _GEN_1906; // @[executor.scala 473:84]
  wire [7:0] _GEN_2791 = _GEN_8842 == 8'h5c ? _GEN_2787 : _GEN_1907; // @[executor.scala 473:84]
  wire [7:0] _GEN_2792 = _GEN_8842 == 8'h5c ? _GEN_2788 : _GEN_1908; // @[executor.scala 473:84]
  wire [7:0] _GEN_2793 = _GEN_8842 == 8'h5c ? _GEN_2789 : _GEN_1909; // @[executor.scala 473:84]
  wire [7:0] _GEN_2794 = mask_1[0] ? byte_512 : _GEN_1910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2795 = mask_1[1] ? byte_513 : _GEN_1911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2796 = mask_1[2] ? byte_514 : _GEN_1912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2797 = mask_1[3] ? byte_515 : _GEN_1913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2798 = _GEN_8842 == 8'h5d ? _GEN_2794 : _GEN_1910; // @[executor.scala 473:84]
  wire [7:0] _GEN_2799 = _GEN_8842 == 8'h5d ? _GEN_2795 : _GEN_1911; // @[executor.scala 473:84]
  wire [7:0] _GEN_2800 = _GEN_8842 == 8'h5d ? _GEN_2796 : _GEN_1912; // @[executor.scala 473:84]
  wire [7:0] _GEN_2801 = _GEN_8842 == 8'h5d ? _GEN_2797 : _GEN_1913; // @[executor.scala 473:84]
  wire [7:0] _GEN_2802 = mask_1[0] ? byte_512 : _GEN_1914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2803 = mask_1[1] ? byte_513 : _GEN_1915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2804 = mask_1[2] ? byte_514 : _GEN_1916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2805 = mask_1[3] ? byte_515 : _GEN_1917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2806 = _GEN_8842 == 8'h5e ? _GEN_2802 : _GEN_1914; // @[executor.scala 473:84]
  wire [7:0] _GEN_2807 = _GEN_8842 == 8'h5e ? _GEN_2803 : _GEN_1915; // @[executor.scala 473:84]
  wire [7:0] _GEN_2808 = _GEN_8842 == 8'h5e ? _GEN_2804 : _GEN_1916; // @[executor.scala 473:84]
  wire [7:0] _GEN_2809 = _GEN_8842 == 8'h5e ? _GEN_2805 : _GEN_1917; // @[executor.scala 473:84]
  wire [7:0] _GEN_2810 = mask_1[0] ? byte_512 : _GEN_1918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2811 = mask_1[1] ? byte_513 : _GEN_1919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2812 = mask_1[2] ? byte_514 : _GEN_1920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2813 = mask_1[3] ? byte_515 : _GEN_1921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2814 = _GEN_8842 == 8'h5f ? _GEN_2810 : _GEN_1918; // @[executor.scala 473:84]
  wire [7:0] _GEN_2815 = _GEN_8842 == 8'h5f ? _GEN_2811 : _GEN_1919; // @[executor.scala 473:84]
  wire [7:0] _GEN_2816 = _GEN_8842 == 8'h5f ? _GEN_2812 : _GEN_1920; // @[executor.scala 473:84]
  wire [7:0] _GEN_2817 = _GEN_8842 == 8'h5f ? _GEN_2813 : _GEN_1921; // @[executor.scala 473:84]
  wire [7:0] _GEN_2818 = mask_1[0] ? byte_512 : _GEN_1922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2819 = mask_1[1] ? byte_513 : _GEN_1923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2820 = mask_1[2] ? byte_514 : _GEN_1924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2821 = mask_1[3] ? byte_515 : _GEN_1925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2822 = _GEN_8842 == 8'h60 ? _GEN_2818 : _GEN_1922; // @[executor.scala 473:84]
  wire [7:0] _GEN_2823 = _GEN_8842 == 8'h60 ? _GEN_2819 : _GEN_1923; // @[executor.scala 473:84]
  wire [7:0] _GEN_2824 = _GEN_8842 == 8'h60 ? _GEN_2820 : _GEN_1924; // @[executor.scala 473:84]
  wire [7:0] _GEN_2825 = _GEN_8842 == 8'h60 ? _GEN_2821 : _GEN_1925; // @[executor.scala 473:84]
  wire [7:0] _GEN_2826 = mask_1[0] ? byte_512 : _GEN_1926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2827 = mask_1[1] ? byte_513 : _GEN_1927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2828 = mask_1[2] ? byte_514 : _GEN_1928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2829 = mask_1[3] ? byte_515 : _GEN_1929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2830 = _GEN_8842 == 8'h61 ? _GEN_2826 : _GEN_1926; // @[executor.scala 473:84]
  wire [7:0] _GEN_2831 = _GEN_8842 == 8'h61 ? _GEN_2827 : _GEN_1927; // @[executor.scala 473:84]
  wire [7:0] _GEN_2832 = _GEN_8842 == 8'h61 ? _GEN_2828 : _GEN_1928; // @[executor.scala 473:84]
  wire [7:0] _GEN_2833 = _GEN_8842 == 8'h61 ? _GEN_2829 : _GEN_1929; // @[executor.scala 473:84]
  wire [7:0] _GEN_2834 = mask_1[0] ? byte_512 : _GEN_1930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2835 = mask_1[1] ? byte_513 : _GEN_1931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2836 = mask_1[2] ? byte_514 : _GEN_1932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2837 = mask_1[3] ? byte_515 : _GEN_1933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2838 = _GEN_8842 == 8'h62 ? _GEN_2834 : _GEN_1930; // @[executor.scala 473:84]
  wire [7:0] _GEN_2839 = _GEN_8842 == 8'h62 ? _GEN_2835 : _GEN_1931; // @[executor.scala 473:84]
  wire [7:0] _GEN_2840 = _GEN_8842 == 8'h62 ? _GEN_2836 : _GEN_1932; // @[executor.scala 473:84]
  wire [7:0] _GEN_2841 = _GEN_8842 == 8'h62 ? _GEN_2837 : _GEN_1933; // @[executor.scala 473:84]
  wire [7:0] _GEN_2842 = mask_1[0] ? byte_512 : _GEN_1934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2843 = mask_1[1] ? byte_513 : _GEN_1935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2844 = mask_1[2] ? byte_514 : _GEN_1936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2845 = mask_1[3] ? byte_515 : _GEN_1937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2846 = _GEN_8842 == 8'h63 ? _GEN_2842 : _GEN_1934; // @[executor.scala 473:84]
  wire [7:0] _GEN_2847 = _GEN_8842 == 8'h63 ? _GEN_2843 : _GEN_1935; // @[executor.scala 473:84]
  wire [7:0] _GEN_2848 = _GEN_8842 == 8'h63 ? _GEN_2844 : _GEN_1936; // @[executor.scala 473:84]
  wire [7:0] _GEN_2849 = _GEN_8842 == 8'h63 ? _GEN_2845 : _GEN_1937; // @[executor.scala 473:84]
  wire [7:0] _GEN_2850 = mask_1[0] ? byte_512 : _GEN_1938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2851 = mask_1[1] ? byte_513 : _GEN_1939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2852 = mask_1[2] ? byte_514 : _GEN_1940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2853 = mask_1[3] ? byte_515 : _GEN_1941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2854 = _GEN_8842 == 8'h64 ? _GEN_2850 : _GEN_1938; // @[executor.scala 473:84]
  wire [7:0] _GEN_2855 = _GEN_8842 == 8'h64 ? _GEN_2851 : _GEN_1939; // @[executor.scala 473:84]
  wire [7:0] _GEN_2856 = _GEN_8842 == 8'h64 ? _GEN_2852 : _GEN_1940; // @[executor.scala 473:84]
  wire [7:0] _GEN_2857 = _GEN_8842 == 8'h64 ? _GEN_2853 : _GEN_1941; // @[executor.scala 473:84]
  wire [7:0] _GEN_2858 = mask_1[0] ? byte_512 : _GEN_1942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2859 = mask_1[1] ? byte_513 : _GEN_1943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2860 = mask_1[2] ? byte_514 : _GEN_1944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2861 = mask_1[3] ? byte_515 : _GEN_1945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2862 = _GEN_8842 == 8'h65 ? _GEN_2858 : _GEN_1942; // @[executor.scala 473:84]
  wire [7:0] _GEN_2863 = _GEN_8842 == 8'h65 ? _GEN_2859 : _GEN_1943; // @[executor.scala 473:84]
  wire [7:0] _GEN_2864 = _GEN_8842 == 8'h65 ? _GEN_2860 : _GEN_1944; // @[executor.scala 473:84]
  wire [7:0] _GEN_2865 = _GEN_8842 == 8'h65 ? _GEN_2861 : _GEN_1945; // @[executor.scala 473:84]
  wire [7:0] _GEN_2866 = mask_1[0] ? byte_512 : _GEN_1946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2867 = mask_1[1] ? byte_513 : _GEN_1947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2868 = mask_1[2] ? byte_514 : _GEN_1948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2869 = mask_1[3] ? byte_515 : _GEN_1949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2870 = _GEN_8842 == 8'h66 ? _GEN_2866 : _GEN_1946; // @[executor.scala 473:84]
  wire [7:0] _GEN_2871 = _GEN_8842 == 8'h66 ? _GEN_2867 : _GEN_1947; // @[executor.scala 473:84]
  wire [7:0] _GEN_2872 = _GEN_8842 == 8'h66 ? _GEN_2868 : _GEN_1948; // @[executor.scala 473:84]
  wire [7:0] _GEN_2873 = _GEN_8842 == 8'h66 ? _GEN_2869 : _GEN_1949; // @[executor.scala 473:84]
  wire [7:0] _GEN_2874 = mask_1[0] ? byte_512 : _GEN_1950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2875 = mask_1[1] ? byte_513 : _GEN_1951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2876 = mask_1[2] ? byte_514 : _GEN_1952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2877 = mask_1[3] ? byte_515 : _GEN_1953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2878 = _GEN_8842 == 8'h67 ? _GEN_2874 : _GEN_1950; // @[executor.scala 473:84]
  wire [7:0] _GEN_2879 = _GEN_8842 == 8'h67 ? _GEN_2875 : _GEN_1951; // @[executor.scala 473:84]
  wire [7:0] _GEN_2880 = _GEN_8842 == 8'h67 ? _GEN_2876 : _GEN_1952; // @[executor.scala 473:84]
  wire [7:0] _GEN_2881 = _GEN_8842 == 8'h67 ? _GEN_2877 : _GEN_1953; // @[executor.scala 473:84]
  wire [7:0] _GEN_2882 = mask_1[0] ? byte_512 : _GEN_1954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2883 = mask_1[1] ? byte_513 : _GEN_1955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2884 = mask_1[2] ? byte_514 : _GEN_1956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2885 = mask_1[3] ? byte_515 : _GEN_1957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2886 = _GEN_8842 == 8'h68 ? _GEN_2882 : _GEN_1954; // @[executor.scala 473:84]
  wire [7:0] _GEN_2887 = _GEN_8842 == 8'h68 ? _GEN_2883 : _GEN_1955; // @[executor.scala 473:84]
  wire [7:0] _GEN_2888 = _GEN_8842 == 8'h68 ? _GEN_2884 : _GEN_1956; // @[executor.scala 473:84]
  wire [7:0] _GEN_2889 = _GEN_8842 == 8'h68 ? _GEN_2885 : _GEN_1957; // @[executor.scala 473:84]
  wire [7:0] _GEN_2890 = mask_1[0] ? byte_512 : _GEN_1958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2891 = mask_1[1] ? byte_513 : _GEN_1959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2892 = mask_1[2] ? byte_514 : _GEN_1960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2893 = mask_1[3] ? byte_515 : _GEN_1961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2894 = _GEN_8842 == 8'h69 ? _GEN_2890 : _GEN_1958; // @[executor.scala 473:84]
  wire [7:0] _GEN_2895 = _GEN_8842 == 8'h69 ? _GEN_2891 : _GEN_1959; // @[executor.scala 473:84]
  wire [7:0] _GEN_2896 = _GEN_8842 == 8'h69 ? _GEN_2892 : _GEN_1960; // @[executor.scala 473:84]
  wire [7:0] _GEN_2897 = _GEN_8842 == 8'h69 ? _GEN_2893 : _GEN_1961; // @[executor.scala 473:84]
  wire [7:0] _GEN_2898 = mask_1[0] ? byte_512 : _GEN_1962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2899 = mask_1[1] ? byte_513 : _GEN_1963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2900 = mask_1[2] ? byte_514 : _GEN_1964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2901 = mask_1[3] ? byte_515 : _GEN_1965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2902 = _GEN_8842 == 8'h6a ? _GEN_2898 : _GEN_1962; // @[executor.scala 473:84]
  wire [7:0] _GEN_2903 = _GEN_8842 == 8'h6a ? _GEN_2899 : _GEN_1963; // @[executor.scala 473:84]
  wire [7:0] _GEN_2904 = _GEN_8842 == 8'h6a ? _GEN_2900 : _GEN_1964; // @[executor.scala 473:84]
  wire [7:0] _GEN_2905 = _GEN_8842 == 8'h6a ? _GEN_2901 : _GEN_1965; // @[executor.scala 473:84]
  wire [7:0] _GEN_2906 = mask_1[0] ? byte_512 : _GEN_1966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2907 = mask_1[1] ? byte_513 : _GEN_1967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2908 = mask_1[2] ? byte_514 : _GEN_1968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2909 = mask_1[3] ? byte_515 : _GEN_1969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2910 = _GEN_8842 == 8'h6b ? _GEN_2906 : _GEN_1966; // @[executor.scala 473:84]
  wire [7:0] _GEN_2911 = _GEN_8842 == 8'h6b ? _GEN_2907 : _GEN_1967; // @[executor.scala 473:84]
  wire [7:0] _GEN_2912 = _GEN_8842 == 8'h6b ? _GEN_2908 : _GEN_1968; // @[executor.scala 473:84]
  wire [7:0] _GEN_2913 = _GEN_8842 == 8'h6b ? _GEN_2909 : _GEN_1969; // @[executor.scala 473:84]
  wire [7:0] _GEN_2914 = mask_1[0] ? byte_512 : _GEN_1970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2915 = mask_1[1] ? byte_513 : _GEN_1971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2916 = mask_1[2] ? byte_514 : _GEN_1972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2917 = mask_1[3] ? byte_515 : _GEN_1973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2918 = _GEN_8842 == 8'h6c ? _GEN_2914 : _GEN_1970; // @[executor.scala 473:84]
  wire [7:0] _GEN_2919 = _GEN_8842 == 8'h6c ? _GEN_2915 : _GEN_1971; // @[executor.scala 473:84]
  wire [7:0] _GEN_2920 = _GEN_8842 == 8'h6c ? _GEN_2916 : _GEN_1972; // @[executor.scala 473:84]
  wire [7:0] _GEN_2921 = _GEN_8842 == 8'h6c ? _GEN_2917 : _GEN_1973; // @[executor.scala 473:84]
  wire [7:0] _GEN_2922 = mask_1[0] ? byte_512 : _GEN_1974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2923 = mask_1[1] ? byte_513 : _GEN_1975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2924 = mask_1[2] ? byte_514 : _GEN_1976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2925 = mask_1[3] ? byte_515 : _GEN_1977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2926 = _GEN_8842 == 8'h6d ? _GEN_2922 : _GEN_1974; // @[executor.scala 473:84]
  wire [7:0] _GEN_2927 = _GEN_8842 == 8'h6d ? _GEN_2923 : _GEN_1975; // @[executor.scala 473:84]
  wire [7:0] _GEN_2928 = _GEN_8842 == 8'h6d ? _GEN_2924 : _GEN_1976; // @[executor.scala 473:84]
  wire [7:0] _GEN_2929 = _GEN_8842 == 8'h6d ? _GEN_2925 : _GEN_1977; // @[executor.scala 473:84]
  wire [7:0] _GEN_2930 = mask_1[0] ? byte_512 : _GEN_1978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2931 = mask_1[1] ? byte_513 : _GEN_1979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2932 = mask_1[2] ? byte_514 : _GEN_1980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2933 = mask_1[3] ? byte_515 : _GEN_1981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2934 = _GEN_8842 == 8'h6e ? _GEN_2930 : _GEN_1978; // @[executor.scala 473:84]
  wire [7:0] _GEN_2935 = _GEN_8842 == 8'h6e ? _GEN_2931 : _GEN_1979; // @[executor.scala 473:84]
  wire [7:0] _GEN_2936 = _GEN_8842 == 8'h6e ? _GEN_2932 : _GEN_1980; // @[executor.scala 473:84]
  wire [7:0] _GEN_2937 = _GEN_8842 == 8'h6e ? _GEN_2933 : _GEN_1981; // @[executor.scala 473:84]
  wire [7:0] _GEN_2938 = mask_1[0] ? byte_512 : _GEN_1982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2939 = mask_1[1] ? byte_513 : _GEN_1983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2940 = mask_1[2] ? byte_514 : _GEN_1984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2941 = mask_1[3] ? byte_515 : _GEN_1985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2942 = _GEN_8842 == 8'h6f ? _GEN_2938 : _GEN_1982; // @[executor.scala 473:84]
  wire [7:0] _GEN_2943 = _GEN_8842 == 8'h6f ? _GEN_2939 : _GEN_1983; // @[executor.scala 473:84]
  wire [7:0] _GEN_2944 = _GEN_8842 == 8'h6f ? _GEN_2940 : _GEN_1984; // @[executor.scala 473:84]
  wire [7:0] _GEN_2945 = _GEN_8842 == 8'h6f ? _GEN_2941 : _GEN_1985; // @[executor.scala 473:84]
  wire [7:0] _GEN_2946 = mask_1[0] ? byte_512 : _GEN_1986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2947 = mask_1[1] ? byte_513 : _GEN_1987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2948 = mask_1[2] ? byte_514 : _GEN_1988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2949 = mask_1[3] ? byte_515 : _GEN_1989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2950 = _GEN_8842 == 8'h70 ? _GEN_2946 : _GEN_1986; // @[executor.scala 473:84]
  wire [7:0] _GEN_2951 = _GEN_8842 == 8'h70 ? _GEN_2947 : _GEN_1987; // @[executor.scala 473:84]
  wire [7:0] _GEN_2952 = _GEN_8842 == 8'h70 ? _GEN_2948 : _GEN_1988; // @[executor.scala 473:84]
  wire [7:0] _GEN_2953 = _GEN_8842 == 8'h70 ? _GEN_2949 : _GEN_1989; // @[executor.scala 473:84]
  wire [7:0] _GEN_2954 = mask_1[0] ? byte_512 : _GEN_1990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2955 = mask_1[1] ? byte_513 : _GEN_1991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2956 = mask_1[2] ? byte_514 : _GEN_1992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2957 = mask_1[3] ? byte_515 : _GEN_1993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2958 = _GEN_8842 == 8'h71 ? _GEN_2954 : _GEN_1990; // @[executor.scala 473:84]
  wire [7:0] _GEN_2959 = _GEN_8842 == 8'h71 ? _GEN_2955 : _GEN_1991; // @[executor.scala 473:84]
  wire [7:0] _GEN_2960 = _GEN_8842 == 8'h71 ? _GEN_2956 : _GEN_1992; // @[executor.scala 473:84]
  wire [7:0] _GEN_2961 = _GEN_8842 == 8'h71 ? _GEN_2957 : _GEN_1993; // @[executor.scala 473:84]
  wire [7:0] _GEN_2962 = mask_1[0] ? byte_512 : _GEN_1994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2963 = mask_1[1] ? byte_513 : _GEN_1995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2964 = mask_1[2] ? byte_514 : _GEN_1996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2965 = mask_1[3] ? byte_515 : _GEN_1997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2966 = _GEN_8842 == 8'h72 ? _GEN_2962 : _GEN_1994; // @[executor.scala 473:84]
  wire [7:0] _GEN_2967 = _GEN_8842 == 8'h72 ? _GEN_2963 : _GEN_1995; // @[executor.scala 473:84]
  wire [7:0] _GEN_2968 = _GEN_8842 == 8'h72 ? _GEN_2964 : _GEN_1996; // @[executor.scala 473:84]
  wire [7:0] _GEN_2969 = _GEN_8842 == 8'h72 ? _GEN_2965 : _GEN_1997; // @[executor.scala 473:84]
  wire [7:0] _GEN_2970 = mask_1[0] ? byte_512 : _GEN_1998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2971 = mask_1[1] ? byte_513 : _GEN_1999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2972 = mask_1[2] ? byte_514 : _GEN_2000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2973 = mask_1[3] ? byte_515 : _GEN_2001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2974 = _GEN_8842 == 8'h73 ? _GEN_2970 : _GEN_1998; // @[executor.scala 473:84]
  wire [7:0] _GEN_2975 = _GEN_8842 == 8'h73 ? _GEN_2971 : _GEN_1999; // @[executor.scala 473:84]
  wire [7:0] _GEN_2976 = _GEN_8842 == 8'h73 ? _GEN_2972 : _GEN_2000; // @[executor.scala 473:84]
  wire [7:0] _GEN_2977 = _GEN_8842 == 8'h73 ? _GEN_2973 : _GEN_2001; // @[executor.scala 473:84]
  wire [7:0] _GEN_2978 = mask_1[0] ? byte_512 : _GEN_2002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2979 = mask_1[1] ? byte_513 : _GEN_2003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2980 = mask_1[2] ? byte_514 : _GEN_2004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2981 = mask_1[3] ? byte_515 : _GEN_2005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2982 = _GEN_8842 == 8'h74 ? _GEN_2978 : _GEN_2002; // @[executor.scala 473:84]
  wire [7:0] _GEN_2983 = _GEN_8842 == 8'h74 ? _GEN_2979 : _GEN_2003; // @[executor.scala 473:84]
  wire [7:0] _GEN_2984 = _GEN_8842 == 8'h74 ? _GEN_2980 : _GEN_2004; // @[executor.scala 473:84]
  wire [7:0] _GEN_2985 = _GEN_8842 == 8'h74 ? _GEN_2981 : _GEN_2005; // @[executor.scala 473:84]
  wire [7:0] _GEN_2986 = mask_1[0] ? byte_512 : _GEN_2006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2987 = mask_1[1] ? byte_513 : _GEN_2007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2988 = mask_1[2] ? byte_514 : _GEN_2008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2989 = mask_1[3] ? byte_515 : _GEN_2009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2990 = _GEN_8842 == 8'h75 ? _GEN_2986 : _GEN_2006; // @[executor.scala 473:84]
  wire [7:0] _GEN_2991 = _GEN_8842 == 8'h75 ? _GEN_2987 : _GEN_2007; // @[executor.scala 473:84]
  wire [7:0] _GEN_2992 = _GEN_8842 == 8'h75 ? _GEN_2988 : _GEN_2008; // @[executor.scala 473:84]
  wire [7:0] _GEN_2993 = _GEN_8842 == 8'h75 ? _GEN_2989 : _GEN_2009; // @[executor.scala 473:84]
  wire [7:0] _GEN_2994 = mask_1[0] ? byte_512 : _GEN_2010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2995 = mask_1[1] ? byte_513 : _GEN_2011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2996 = mask_1[2] ? byte_514 : _GEN_2012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2997 = mask_1[3] ? byte_515 : _GEN_2013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_2998 = _GEN_8842 == 8'h76 ? _GEN_2994 : _GEN_2010; // @[executor.scala 473:84]
  wire [7:0] _GEN_2999 = _GEN_8842 == 8'h76 ? _GEN_2995 : _GEN_2011; // @[executor.scala 473:84]
  wire [7:0] _GEN_3000 = _GEN_8842 == 8'h76 ? _GEN_2996 : _GEN_2012; // @[executor.scala 473:84]
  wire [7:0] _GEN_3001 = _GEN_8842 == 8'h76 ? _GEN_2997 : _GEN_2013; // @[executor.scala 473:84]
  wire [7:0] _GEN_3002 = mask_1[0] ? byte_512 : _GEN_2014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3003 = mask_1[1] ? byte_513 : _GEN_2015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3004 = mask_1[2] ? byte_514 : _GEN_2016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3005 = mask_1[3] ? byte_515 : _GEN_2017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3006 = _GEN_8842 == 8'h77 ? _GEN_3002 : _GEN_2014; // @[executor.scala 473:84]
  wire [7:0] _GEN_3007 = _GEN_8842 == 8'h77 ? _GEN_3003 : _GEN_2015; // @[executor.scala 473:84]
  wire [7:0] _GEN_3008 = _GEN_8842 == 8'h77 ? _GEN_3004 : _GEN_2016; // @[executor.scala 473:84]
  wire [7:0] _GEN_3009 = _GEN_8842 == 8'h77 ? _GEN_3005 : _GEN_2017; // @[executor.scala 473:84]
  wire [7:0] _GEN_3010 = mask_1[0] ? byte_512 : _GEN_2018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3011 = mask_1[1] ? byte_513 : _GEN_2019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3012 = mask_1[2] ? byte_514 : _GEN_2020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3013 = mask_1[3] ? byte_515 : _GEN_2021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3014 = _GEN_8842 == 8'h78 ? _GEN_3010 : _GEN_2018; // @[executor.scala 473:84]
  wire [7:0] _GEN_3015 = _GEN_8842 == 8'h78 ? _GEN_3011 : _GEN_2019; // @[executor.scala 473:84]
  wire [7:0] _GEN_3016 = _GEN_8842 == 8'h78 ? _GEN_3012 : _GEN_2020; // @[executor.scala 473:84]
  wire [7:0] _GEN_3017 = _GEN_8842 == 8'h78 ? _GEN_3013 : _GEN_2021; // @[executor.scala 473:84]
  wire [7:0] _GEN_3018 = mask_1[0] ? byte_512 : _GEN_2022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3019 = mask_1[1] ? byte_513 : _GEN_2023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3020 = mask_1[2] ? byte_514 : _GEN_2024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3021 = mask_1[3] ? byte_515 : _GEN_2025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3022 = _GEN_8842 == 8'h79 ? _GEN_3018 : _GEN_2022; // @[executor.scala 473:84]
  wire [7:0] _GEN_3023 = _GEN_8842 == 8'h79 ? _GEN_3019 : _GEN_2023; // @[executor.scala 473:84]
  wire [7:0] _GEN_3024 = _GEN_8842 == 8'h79 ? _GEN_3020 : _GEN_2024; // @[executor.scala 473:84]
  wire [7:0] _GEN_3025 = _GEN_8842 == 8'h79 ? _GEN_3021 : _GEN_2025; // @[executor.scala 473:84]
  wire [7:0] _GEN_3026 = mask_1[0] ? byte_512 : _GEN_2026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3027 = mask_1[1] ? byte_513 : _GEN_2027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3028 = mask_1[2] ? byte_514 : _GEN_2028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3029 = mask_1[3] ? byte_515 : _GEN_2029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3030 = _GEN_8842 == 8'h7a ? _GEN_3026 : _GEN_2026; // @[executor.scala 473:84]
  wire [7:0] _GEN_3031 = _GEN_8842 == 8'h7a ? _GEN_3027 : _GEN_2027; // @[executor.scala 473:84]
  wire [7:0] _GEN_3032 = _GEN_8842 == 8'h7a ? _GEN_3028 : _GEN_2028; // @[executor.scala 473:84]
  wire [7:0] _GEN_3033 = _GEN_8842 == 8'h7a ? _GEN_3029 : _GEN_2029; // @[executor.scala 473:84]
  wire [7:0] _GEN_3034 = mask_1[0] ? byte_512 : _GEN_2030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3035 = mask_1[1] ? byte_513 : _GEN_2031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3036 = mask_1[2] ? byte_514 : _GEN_2032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3037 = mask_1[3] ? byte_515 : _GEN_2033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3038 = _GEN_8842 == 8'h7b ? _GEN_3034 : _GEN_2030; // @[executor.scala 473:84]
  wire [7:0] _GEN_3039 = _GEN_8842 == 8'h7b ? _GEN_3035 : _GEN_2031; // @[executor.scala 473:84]
  wire [7:0] _GEN_3040 = _GEN_8842 == 8'h7b ? _GEN_3036 : _GEN_2032; // @[executor.scala 473:84]
  wire [7:0] _GEN_3041 = _GEN_8842 == 8'h7b ? _GEN_3037 : _GEN_2033; // @[executor.scala 473:84]
  wire [7:0] _GEN_3042 = mask_1[0] ? byte_512 : _GEN_2034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3043 = mask_1[1] ? byte_513 : _GEN_2035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3044 = mask_1[2] ? byte_514 : _GEN_2036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3045 = mask_1[3] ? byte_515 : _GEN_2037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3046 = _GEN_8842 == 8'h7c ? _GEN_3042 : _GEN_2034; // @[executor.scala 473:84]
  wire [7:0] _GEN_3047 = _GEN_8842 == 8'h7c ? _GEN_3043 : _GEN_2035; // @[executor.scala 473:84]
  wire [7:0] _GEN_3048 = _GEN_8842 == 8'h7c ? _GEN_3044 : _GEN_2036; // @[executor.scala 473:84]
  wire [7:0] _GEN_3049 = _GEN_8842 == 8'h7c ? _GEN_3045 : _GEN_2037; // @[executor.scala 473:84]
  wire [7:0] _GEN_3050 = mask_1[0] ? byte_512 : _GEN_2038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3051 = mask_1[1] ? byte_513 : _GEN_2039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3052 = mask_1[2] ? byte_514 : _GEN_2040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3053 = mask_1[3] ? byte_515 : _GEN_2041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3054 = _GEN_8842 == 8'h7d ? _GEN_3050 : _GEN_2038; // @[executor.scala 473:84]
  wire [7:0] _GEN_3055 = _GEN_8842 == 8'h7d ? _GEN_3051 : _GEN_2039; // @[executor.scala 473:84]
  wire [7:0] _GEN_3056 = _GEN_8842 == 8'h7d ? _GEN_3052 : _GEN_2040; // @[executor.scala 473:84]
  wire [7:0] _GEN_3057 = _GEN_8842 == 8'h7d ? _GEN_3053 : _GEN_2041; // @[executor.scala 473:84]
  wire [7:0] _GEN_3058 = mask_1[0] ? byte_512 : _GEN_2042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3059 = mask_1[1] ? byte_513 : _GEN_2043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3060 = mask_1[2] ? byte_514 : _GEN_2044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3061 = mask_1[3] ? byte_515 : _GEN_2045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3062 = _GEN_8842 == 8'h7e ? _GEN_3058 : _GEN_2042; // @[executor.scala 473:84]
  wire [7:0] _GEN_3063 = _GEN_8842 == 8'h7e ? _GEN_3059 : _GEN_2043; // @[executor.scala 473:84]
  wire [7:0] _GEN_3064 = _GEN_8842 == 8'h7e ? _GEN_3060 : _GEN_2044; // @[executor.scala 473:84]
  wire [7:0] _GEN_3065 = _GEN_8842 == 8'h7e ? _GEN_3061 : _GEN_2045; // @[executor.scala 473:84]
  wire [7:0] _GEN_3066 = mask_1[0] ? byte_512 : _GEN_2046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3067 = mask_1[1] ? byte_513 : _GEN_2047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3068 = mask_1[2] ? byte_514 : _GEN_2048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3069 = mask_1[3] ? byte_515 : _GEN_2049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_3070 = _GEN_8842 == 8'h7f ? _GEN_3066 : _GEN_2046; // @[executor.scala 473:84]
  wire [7:0] _GEN_3071 = _GEN_8842 == 8'h7f ? _GEN_3067 : _GEN_2047; // @[executor.scala 473:84]
  wire [7:0] _GEN_3072 = _GEN_8842 == 8'h7f ? _GEN_3068 : _GEN_2048; // @[executor.scala 473:84]
  wire [7:0] _GEN_3073 = _GEN_8842 == 8'h7f ? _GEN_3069 : _GEN_2049; // @[executor.scala 473:84]
  wire [7:0] _GEN_3074 = opcode_1 != 4'h0 ? _GEN_2054 : _GEN_1538; // @[executor.scala 470:55]
  wire [7:0] _GEN_3075 = opcode_1 != 4'h0 ? _GEN_2055 : _GEN_1539; // @[executor.scala 470:55]
  wire [7:0] _GEN_3076 = opcode_1 != 4'h0 ? _GEN_2056 : _GEN_1540; // @[executor.scala 470:55]
  wire [7:0] _GEN_3077 = opcode_1 != 4'h0 ? _GEN_2057 : _GEN_1541; // @[executor.scala 470:55]
  wire [7:0] _GEN_3078 = opcode_1 != 4'h0 ? _GEN_2062 : _GEN_1542; // @[executor.scala 470:55]
  wire [7:0] _GEN_3079 = opcode_1 != 4'h0 ? _GEN_2063 : _GEN_1543; // @[executor.scala 470:55]
  wire [7:0] _GEN_3080 = opcode_1 != 4'h0 ? _GEN_2064 : _GEN_1544; // @[executor.scala 470:55]
  wire [7:0] _GEN_3081 = opcode_1 != 4'h0 ? _GEN_2065 : _GEN_1545; // @[executor.scala 470:55]
  wire [7:0] _GEN_3082 = opcode_1 != 4'h0 ? _GEN_2070 : _GEN_1546; // @[executor.scala 470:55]
  wire [7:0] _GEN_3083 = opcode_1 != 4'h0 ? _GEN_2071 : _GEN_1547; // @[executor.scala 470:55]
  wire [7:0] _GEN_3084 = opcode_1 != 4'h0 ? _GEN_2072 : _GEN_1548; // @[executor.scala 470:55]
  wire [7:0] _GEN_3085 = opcode_1 != 4'h0 ? _GEN_2073 : _GEN_1549; // @[executor.scala 470:55]
  wire [7:0] _GEN_3086 = opcode_1 != 4'h0 ? _GEN_2078 : _GEN_1550; // @[executor.scala 470:55]
  wire [7:0] _GEN_3087 = opcode_1 != 4'h0 ? _GEN_2079 : _GEN_1551; // @[executor.scala 470:55]
  wire [7:0] _GEN_3088 = opcode_1 != 4'h0 ? _GEN_2080 : _GEN_1552; // @[executor.scala 470:55]
  wire [7:0] _GEN_3089 = opcode_1 != 4'h0 ? _GEN_2081 : _GEN_1553; // @[executor.scala 470:55]
  wire [7:0] _GEN_3090 = opcode_1 != 4'h0 ? _GEN_2086 : _GEN_1554; // @[executor.scala 470:55]
  wire [7:0] _GEN_3091 = opcode_1 != 4'h0 ? _GEN_2087 : _GEN_1555; // @[executor.scala 470:55]
  wire [7:0] _GEN_3092 = opcode_1 != 4'h0 ? _GEN_2088 : _GEN_1556; // @[executor.scala 470:55]
  wire [7:0] _GEN_3093 = opcode_1 != 4'h0 ? _GEN_2089 : _GEN_1557; // @[executor.scala 470:55]
  wire [7:0] _GEN_3094 = opcode_1 != 4'h0 ? _GEN_2094 : _GEN_1558; // @[executor.scala 470:55]
  wire [7:0] _GEN_3095 = opcode_1 != 4'h0 ? _GEN_2095 : _GEN_1559; // @[executor.scala 470:55]
  wire [7:0] _GEN_3096 = opcode_1 != 4'h0 ? _GEN_2096 : _GEN_1560; // @[executor.scala 470:55]
  wire [7:0] _GEN_3097 = opcode_1 != 4'h0 ? _GEN_2097 : _GEN_1561; // @[executor.scala 470:55]
  wire [7:0] _GEN_3098 = opcode_1 != 4'h0 ? _GEN_2102 : _GEN_1562; // @[executor.scala 470:55]
  wire [7:0] _GEN_3099 = opcode_1 != 4'h0 ? _GEN_2103 : _GEN_1563; // @[executor.scala 470:55]
  wire [7:0] _GEN_3100 = opcode_1 != 4'h0 ? _GEN_2104 : _GEN_1564; // @[executor.scala 470:55]
  wire [7:0] _GEN_3101 = opcode_1 != 4'h0 ? _GEN_2105 : _GEN_1565; // @[executor.scala 470:55]
  wire [7:0] _GEN_3102 = opcode_1 != 4'h0 ? _GEN_2110 : _GEN_1566; // @[executor.scala 470:55]
  wire [7:0] _GEN_3103 = opcode_1 != 4'h0 ? _GEN_2111 : _GEN_1567; // @[executor.scala 470:55]
  wire [7:0] _GEN_3104 = opcode_1 != 4'h0 ? _GEN_2112 : _GEN_1568; // @[executor.scala 470:55]
  wire [7:0] _GEN_3105 = opcode_1 != 4'h0 ? _GEN_2113 : _GEN_1569; // @[executor.scala 470:55]
  wire [7:0] _GEN_3106 = opcode_1 != 4'h0 ? _GEN_2118 : _GEN_1570; // @[executor.scala 470:55]
  wire [7:0] _GEN_3107 = opcode_1 != 4'h0 ? _GEN_2119 : _GEN_1571; // @[executor.scala 470:55]
  wire [7:0] _GEN_3108 = opcode_1 != 4'h0 ? _GEN_2120 : _GEN_1572; // @[executor.scala 470:55]
  wire [7:0] _GEN_3109 = opcode_1 != 4'h0 ? _GEN_2121 : _GEN_1573; // @[executor.scala 470:55]
  wire [7:0] _GEN_3110 = opcode_1 != 4'h0 ? _GEN_2126 : _GEN_1574; // @[executor.scala 470:55]
  wire [7:0] _GEN_3111 = opcode_1 != 4'h0 ? _GEN_2127 : _GEN_1575; // @[executor.scala 470:55]
  wire [7:0] _GEN_3112 = opcode_1 != 4'h0 ? _GEN_2128 : _GEN_1576; // @[executor.scala 470:55]
  wire [7:0] _GEN_3113 = opcode_1 != 4'h0 ? _GEN_2129 : _GEN_1577; // @[executor.scala 470:55]
  wire [7:0] _GEN_3114 = opcode_1 != 4'h0 ? _GEN_2134 : _GEN_1578; // @[executor.scala 470:55]
  wire [7:0] _GEN_3115 = opcode_1 != 4'h0 ? _GEN_2135 : _GEN_1579; // @[executor.scala 470:55]
  wire [7:0] _GEN_3116 = opcode_1 != 4'h0 ? _GEN_2136 : _GEN_1580; // @[executor.scala 470:55]
  wire [7:0] _GEN_3117 = opcode_1 != 4'h0 ? _GEN_2137 : _GEN_1581; // @[executor.scala 470:55]
  wire [7:0] _GEN_3118 = opcode_1 != 4'h0 ? _GEN_2142 : _GEN_1582; // @[executor.scala 470:55]
  wire [7:0] _GEN_3119 = opcode_1 != 4'h0 ? _GEN_2143 : _GEN_1583; // @[executor.scala 470:55]
  wire [7:0] _GEN_3120 = opcode_1 != 4'h0 ? _GEN_2144 : _GEN_1584; // @[executor.scala 470:55]
  wire [7:0] _GEN_3121 = opcode_1 != 4'h0 ? _GEN_2145 : _GEN_1585; // @[executor.scala 470:55]
  wire [7:0] _GEN_3122 = opcode_1 != 4'h0 ? _GEN_2150 : _GEN_1586; // @[executor.scala 470:55]
  wire [7:0] _GEN_3123 = opcode_1 != 4'h0 ? _GEN_2151 : _GEN_1587; // @[executor.scala 470:55]
  wire [7:0] _GEN_3124 = opcode_1 != 4'h0 ? _GEN_2152 : _GEN_1588; // @[executor.scala 470:55]
  wire [7:0] _GEN_3125 = opcode_1 != 4'h0 ? _GEN_2153 : _GEN_1589; // @[executor.scala 470:55]
  wire [7:0] _GEN_3126 = opcode_1 != 4'h0 ? _GEN_2158 : _GEN_1590; // @[executor.scala 470:55]
  wire [7:0] _GEN_3127 = opcode_1 != 4'h0 ? _GEN_2159 : _GEN_1591; // @[executor.scala 470:55]
  wire [7:0] _GEN_3128 = opcode_1 != 4'h0 ? _GEN_2160 : _GEN_1592; // @[executor.scala 470:55]
  wire [7:0] _GEN_3129 = opcode_1 != 4'h0 ? _GEN_2161 : _GEN_1593; // @[executor.scala 470:55]
  wire [7:0] _GEN_3130 = opcode_1 != 4'h0 ? _GEN_2166 : _GEN_1594; // @[executor.scala 470:55]
  wire [7:0] _GEN_3131 = opcode_1 != 4'h0 ? _GEN_2167 : _GEN_1595; // @[executor.scala 470:55]
  wire [7:0] _GEN_3132 = opcode_1 != 4'h0 ? _GEN_2168 : _GEN_1596; // @[executor.scala 470:55]
  wire [7:0] _GEN_3133 = opcode_1 != 4'h0 ? _GEN_2169 : _GEN_1597; // @[executor.scala 470:55]
  wire [7:0] _GEN_3134 = opcode_1 != 4'h0 ? _GEN_2174 : _GEN_1598; // @[executor.scala 470:55]
  wire [7:0] _GEN_3135 = opcode_1 != 4'h0 ? _GEN_2175 : _GEN_1599; // @[executor.scala 470:55]
  wire [7:0] _GEN_3136 = opcode_1 != 4'h0 ? _GEN_2176 : _GEN_1600; // @[executor.scala 470:55]
  wire [7:0] _GEN_3137 = opcode_1 != 4'h0 ? _GEN_2177 : _GEN_1601; // @[executor.scala 470:55]
  wire [7:0] _GEN_3138 = opcode_1 != 4'h0 ? _GEN_2182 : _GEN_1602; // @[executor.scala 470:55]
  wire [7:0] _GEN_3139 = opcode_1 != 4'h0 ? _GEN_2183 : _GEN_1603; // @[executor.scala 470:55]
  wire [7:0] _GEN_3140 = opcode_1 != 4'h0 ? _GEN_2184 : _GEN_1604; // @[executor.scala 470:55]
  wire [7:0] _GEN_3141 = opcode_1 != 4'h0 ? _GEN_2185 : _GEN_1605; // @[executor.scala 470:55]
  wire [7:0] _GEN_3142 = opcode_1 != 4'h0 ? _GEN_2190 : _GEN_1606; // @[executor.scala 470:55]
  wire [7:0] _GEN_3143 = opcode_1 != 4'h0 ? _GEN_2191 : _GEN_1607; // @[executor.scala 470:55]
  wire [7:0] _GEN_3144 = opcode_1 != 4'h0 ? _GEN_2192 : _GEN_1608; // @[executor.scala 470:55]
  wire [7:0] _GEN_3145 = opcode_1 != 4'h0 ? _GEN_2193 : _GEN_1609; // @[executor.scala 470:55]
  wire [7:0] _GEN_3146 = opcode_1 != 4'h0 ? _GEN_2198 : _GEN_1610; // @[executor.scala 470:55]
  wire [7:0] _GEN_3147 = opcode_1 != 4'h0 ? _GEN_2199 : _GEN_1611; // @[executor.scala 470:55]
  wire [7:0] _GEN_3148 = opcode_1 != 4'h0 ? _GEN_2200 : _GEN_1612; // @[executor.scala 470:55]
  wire [7:0] _GEN_3149 = opcode_1 != 4'h0 ? _GEN_2201 : _GEN_1613; // @[executor.scala 470:55]
  wire [7:0] _GEN_3150 = opcode_1 != 4'h0 ? _GEN_2206 : _GEN_1614; // @[executor.scala 470:55]
  wire [7:0] _GEN_3151 = opcode_1 != 4'h0 ? _GEN_2207 : _GEN_1615; // @[executor.scala 470:55]
  wire [7:0] _GEN_3152 = opcode_1 != 4'h0 ? _GEN_2208 : _GEN_1616; // @[executor.scala 470:55]
  wire [7:0] _GEN_3153 = opcode_1 != 4'h0 ? _GEN_2209 : _GEN_1617; // @[executor.scala 470:55]
  wire [7:0] _GEN_3154 = opcode_1 != 4'h0 ? _GEN_2214 : _GEN_1618; // @[executor.scala 470:55]
  wire [7:0] _GEN_3155 = opcode_1 != 4'h0 ? _GEN_2215 : _GEN_1619; // @[executor.scala 470:55]
  wire [7:0] _GEN_3156 = opcode_1 != 4'h0 ? _GEN_2216 : _GEN_1620; // @[executor.scala 470:55]
  wire [7:0] _GEN_3157 = opcode_1 != 4'h0 ? _GEN_2217 : _GEN_1621; // @[executor.scala 470:55]
  wire [7:0] _GEN_3158 = opcode_1 != 4'h0 ? _GEN_2222 : _GEN_1622; // @[executor.scala 470:55]
  wire [7:0] _GEN_3159 = opcode_1 != 4'h0 ? _GEN_2223 : _GEN_1623; // @[executor.scala 470:55]
  wire [7:0] _GEN_3160 = opcode_1 != 4'h0 ? _GEN_2224 : _GEN_1624; // @[executor.scala 470:55]
  wire [7:0] _GEN_3161 = opcode_1 != 4'h0 ? _GEN_2225 : _GEN_1625; // @[executor.scala 470:55]
  wire [7:0] _GEN_3162 = opcode_1 != 4'h0 ? _GEN_2230 : _GEN_1626; // @[executor.scala 470:55]
  wire [7:0] _GEN_3163 = opcode_1 != 4'h0 ? _GEN_2231 : _GEN_1627; // @[executor.scala 470:55]
  wire [7:0] _GEN_3164 = opcode_1 != 4'h0 ? _GEN_2232 : _GEN_1628; // @[executor.scala 470:55]
  wire [7:0] _GEN_3165 = opcode_1 != 4'h0 ? _GEN_2233 : _GEN_1629; // @[executor.scala 470:55]
  wire [7:0] _GEN_3166 = opcode_1 != 4'h0 ? _GEN_2238 : _GEN_1630; // @[executor.scala 470:55]
  wire [7:0] _GEN_3167 = opcode_1 != 4'h0 ? _GEN_2239 : _GEN_1631; // @[executor.scala 470:55]
  wire [7:0] _GEN_3168 = opcode_1 != 4'h0 ? _GEN_2240 : _GEN_1632; // @[executor.scala 470:55]
  wire [7:0] _GEN_3169 = opcode_1 != 4'h0 ? _GEN_2241 : _GEN_1633; // @[executor.scala 470:55]
  wire [7:0] _GEN_3170 = opcode_1 != 4'h0 ? _GEN_2246 : _GEN_1634; // @[executor.scala 470:55]
  wire [7:0] _GEN_3171 = opcode_1 != 4'h0 ? _GEN_2247 : _GEN_1635; // @[executor.scala 470:55]
  wire [7:0] _GEN_3172 = opcode_1 != 4'h0 ? _GEN_2248 : _GEN_1636; // @[executor.scala 470:55]
  wire [7:0] _GEN_3173 = opcode_1 != 4'h0 ? _GEN_2249 : _GEN_1637; // @[executor.scala 470:55]
  wire [7:0] _GEN_3174 = opcode_1 != 4'h0 ? _GEN_2254 : _GEN_1638; // @[executor.scala 470:55]
  wire [7:0] _GEN_3175 = opcode_1 != 4'h0 ? _GEN_2255 : _GEN_1639; // @[executor.scala 470:55]
  wire [7:0] _GEN_3176 = opcode_1 != 4'h0 ? _GEN_2256 : _GEN_1640; // @[executor.scala 470:55]
  wire [7:0] _GEN_3177 = opcode_1 != 4'h0 ? _GEN_2257 : _GEN_1641; // @[executor.scala 470:55]
  wire [7:0] _GEN_3178 = opcode_1 != 4'h0 ? _GEN_2262 : _GEN_1642; // @[executor.scala 470:55]
  wire [7:0] _GEN_3179 = opcode_1 != 4'h0 ? _GEN_2263 : _GEN_1643; // @[executor.scala 470:55]
  wire [7:0] _GEN_3180 = opcode_1 != 4'h0 ? _GEN_2264 : _GEN_1644; // @[executor.scala 470:55]
  wire [7:0] _GEN_3181 = opcode_1 != 4'h0 ? _GEN_2265 : _GEN_1645; // @[executor.scala 470:55]
  wire [7:0] _GEN_3182 = opcode_1 != 4'h0 ? _GEN_2270 : _GEN_1646; // @[executor.scala 470:55]
  wire [7:0] _GEN_3183 = opcode_1 != 4'h0 ? _GEN_2271 : _GEN_1647; // @[executor.scala 470:55]
  wire [7:0] _GEN_3184 = opcode_1 != 4'h0 ? _GEN_2272 : _GEN_1648; // @[executor.scala 470:55]
  wire [7:0] _GEN_3185 = opcode_1 != 4'h0 ? _GEN_2273 : _GEN_1649; // @[executor.scala 470:55]
  wire [7:0] _GEN_3186 = opcode_1 != 4'h0 ? _GEN_2278 : _GEN_1650; // @[executor.scala 470:55]
  wire [7:0] _GEN_3187 = opcode_1 != 4'h0 ? _GEN_2279 : _GEN_1651; // @[executor.scala 470:55]
  wire [7:0] _GEN_3188 = opcode_1 != 4'h0 ? _GEN_2280 : _GEN_1652; // @[executor.scala 470:55]
  wire [7:0] _GEN_3189 = opcode_1 != 4'h0 ? _GEN_2281 : _GEN_1653; // @[executor.scala 470:55]
  wire [7:0] _GEN_3190 = opcode_1 != 4'h0 ? _GEN_2286 : _GEN_1654; // @[executor.scala 470:55]
  wire [7:0] _GEN_3191 = opcode_1 != 4'h0 ? _GEN_2287 : _GEN_1655; // @[executor.scala 470:55]
  wire [7:0] _GEN_3192 = opcode_1 != 4'h0 ? _GEN_2288 : _GEN_1656; // @[executor.scala 470:55]
  wire [7:0] _GEN_3193 = opcode_1 != 4'h0 ? _GEN_2289 : _GEN_1657; // @[executor.scala 470:55]
  wire [7:0] _GEN_3194 = opcode_1 != 4'h0 ? _GEN_2294 : _GEN_1658; // @[executor.scala 470:55]
  wire [7:0] _GEN_3195 = opcode_1 != 4'h0 ? _GEN_2295 : _GEN_1659; // @[executor.scala 470:55]
  wire [7:0] _GEN_3196 = opcode_1 != 4'h0 ? _GEN_2296 : _GEN_1660; // @[executor.scala 470:55]
  wire [7:0] _GEN_3197 = opcode_1 != 4'h0 ? _GEN_2297 : _GEN_1661; // @[executor.scala 470:55]
  wire [7:0] _GEN_3198 = opcode_1 != 4'h0 ? _GEN_2302 : _GEN_1662; // @[executor.scala 470:55]
  wire [7:0] _GEN_3199 = opcode_1 != 4'h0 ? _GEN_2303 : _GEN_1663; // @[executor.scala 470:55]
  wire [7:0] _GEN_3200 = opcode_1 != 4'h0 ? _GEN_2304 : _GEN_1664; // @[executor.scala 470:55]
  wire [7:0] _GEN_3201 = opcode_1 != 4'h0 ? _GEN_2305 : _GEN_1665; // @[executor.scala 470:55]
  wire [7:0] _GEN_3202 = opcode_1 != 4'h0 ? _GEN_2310 : _GEN_1666; // @[executor.scala 470:55]
  wire [7:0] _GEN_3203 = opcode_1 != 4'h0 ? _GEN_2311 : _GEN_1667; // @[executor.scala 470:55]
  wire [7:0] _GEN_3204 = opcode_1 != 4'h0 ? _GEN_2312 : _GEN_1668; // @[executor.scala 470:55]
  wire [7:0] _GEN_3205 = opcode_1 != 4'h0 ? _GEN_2313 : _GEN_1669; // @[executor.scala 470:55]
  wire [7:0] _GEN_3206 = opcode_1 != 4'h0 ? _GEN_2318 : _GEN_1670; // @[executor.scala 470:55]
  wire [7:0] _GEN_3207 = opcode_1 != 4'h0 ? _GEN_2319 : _GEN_1671; // @[executor.scala 470:55]
  wire [7:0] _GEN_3208 = opcode_1 != 4'h0 ? _GEN_2320 : _GEN_1672; // @[executor.scala 470:55]
  wire [7:0] _GEN_3209 = opcode_1 != 4'h0 ? _GEN_2321 : _GEN_1673; // @[executor.scala 470:55]
  wire [7:0] _GEN_3210 = opcode_1 != 4'h0 ? _GEN_2326 : _GEN_1674; // @[executor.scala 470:55]
  wire [7:0] _GEN_3211 = opcode_1 != 4'h0 ? _GEN_2327 : _GEN_1675; // @[executor.scala 470:55]
  wire [7:0] _GEN_3212 = opcode_1 != 4'h0 ? _GEN_2328 : _GEN_1676; // @[executor.scala 470:55]
  wire [7:0] _GEN_3213 = opcode_1 != 4'h0 ? _GEN_2329 : _GEN_1677; // @[executor.scala 470:55]
  wire [7:0] _GEN_3214 = opcode_1 != 4'h0 ? _GEN_2334 : _GEN_1678; // @[executor.scala 470:55]
  wire [7:0] _GEN_3215 = opcode_1 != 4'h0 ? _GEN_2335 : _GEN_1679; // @[executor.scala 470:55]
  wire [7:0] _GEN_3216 = opcode_1 != 4'h0 ? _GEN_2336 : _GEN_1680; // @[executor.scala 470:55]
  wire [7:0] _GEN_3217 = opcode_1 != 4'h0 ? _GEN_2337 : _GEN_1681; // @[executor.scala 470:55]
  wire [7:0] _GEN_3218 = opcode_1 != 4'h0 ? _GEN_2342 : _GEN_1682; // @[executor.scala 470:55]
  wire [7:0] _GEN_3219 = opcode_1 != 4'h0 ? _GEN_2343 : _GEN_1683; // @[executor.scala 470:55]
  wire [7:0] _GEN_3220 = opcode_1 != 4'h0 ? _GEN_2344 : _GEN_1684; // @[executor.scala 470:55]
  wire [7:0] _GEN_3221 = opcode_1 != 4'h0 ? _GEN_2345 : _GEN_1685; // @[executor.scala 470:55]
  wire [7:0] _GEN_3222 = opcode_1 != 4'h0 ? _GEN_2350 : _GEN_1686; // @[executor.scala 470:55]
  wire [7:0] _GEN_3223 = opcode_1 != 4'h0 ? _GEN_2351 : _GEN_1687; // @[executor.scala 470:55]
  wire [7:0] _GEN_3224 = opcode_1 != 4'h0 ? _GEN_2352 : _GEN_1688; // @[executor.scala 470:55]
  wire [7:0] _GEN_3225 = opcode_1 != 4'h0 ? _GEN_2353 : _GEN_1689; // @[executor.scala 470:55]
  wire [7:0] _GEN_3226 = opcode_1 != 4'h0 ? _GEN_2358 : _GEN_1690; // @[executor.scala 470:55]
  wire [7:0] _GEN_3227 = opcode_1 != 4'h0 ? _GEN_2359 : _GEN_1691; // @[executor.scala 470:55]
  wire [7:0] _GEN_3228 = opcode_1 != 4'h0 ? _GEN_2360 : _GEN_1692; // @[executor.scala 470:55]
  wire [7:0] _GEN_3229 = opcode_1 != 4'h0 ? _GEN_2361 : _GEN_1693; // @[executor.scala 470:55]
  wire [7:0] _GEN_3230 = opcode_1 != 4'h0 ? _GEN_2366 : _GEN_1694; // @[executor.scala 470:55]
  wire [7:0] _GEN_3231 = opcode_1 != 4'h0 ? _GEN_2367 : _GEN_1695; // @[executor.scala 470:55]
  wire [7:0] _GEN_3232 = opcode_1 != 4'h0 ? _GEN_2368 : _GEN_1696; // @[executor.scala 470:55]
  wire [7:0] _GEN_3233 = opcode_1 != 4'h0 ? _GEN_2369 : _GEN_1697; // @[executor.scala 470:55]
  wire [7:0] _GEN_3234 = opcode_1 != 4'h0 ? _GEN_2374 : _GEN_1698; // @[executor.scala 470:55]
  wire [7:0] _GEN_3235 = opcode_1 != 4'h0 ? _GEN_2375 : _GEN_1699; // @[executor.scala 470:55]
  wire [7:0] _GEN_3236 = opcode_1 != 4'h0 ? _GEN_2376 : _GEN_1700; // @[executor.scala 470:55]
  wire [7:0] _GEN_3237 = opcode_1 != 4'h0 ? _GEN_2377 : _GEN_1701; // @[executor.scala 470:55]
  wire [7:0] _GEN_3238 = opcode_1 != 4'h0 ? _GEN_2382 : _GEN_1702; // @[executor.scala 470:55]
  wire [7:0] _GEN_3239 = opcode_1 != 4'h0 ? _GEN_2383 : _GEN_1703; // @[executor.scala 470:55]
  wire [7:0] _GEN_3240 = opcode_1 != 4'h0 ? _GEN_2384 : _GEN_1704; // @[executor.scala 470:55]
  wire [7:0] _GEN_3241 = opcode_1 != 4'h0 ? _GEN_2385 : _GEN_1705; // @[executor.scala 470:55]
  wire [7:0] _GEN_3242 = opcode_1 != 4'h0 ? _GEN_2390 : _GEN_1706; // @[executor.scala 470:55]
  wire [7:0] _GEN_3243 = opcode_1 != 4'h0 ? _GEN_2391 : _GEN_1707; // @[executor.scala 470:55]
  wire [7:0] _GEN_3244 = opcode_1 != 4'h0 ? _GEN_2392 : _GEN_1708; // @[executor.scala 470:55]
  wire [7:0] _GEN_3245 = opcode_1 != 4'h0 ? _GEN_2393 : _GEN_1709; // @[executor.scala 470:55]
  wire [7:0] _GEN_3246 = opcode_1 != 4'h0 ? _GEN_2398 : _GEN_1710; // @[executor.scala 470:55]
  wire [7:0] _GEN_3247 = opcode_1 != 4'h0 ? _GEN_2399 : _GEN_1711; // @[executor.scala 470:55]
  wire [7:0] _GEN_3248 = opcode_1 != 4'h0 ? _GEN_2400 : _GEN_1712; // @[executor.scala 470:55]
  wire [7:0] _GEN_3249 = opcode_1 != 4'h0 ? _GEN_2401 : _GEN_1713; // @[executor.scala 470:55]
  wire [7:0] _GEN_3250 = opcode_1 != 4'h0 ? _GEN_2406 : _GEN_1714; // @[executor.scala 470:55]
  wire [7:0] _GEN_3251 = opcode_1 != 4'h0 ? _GEN_2407 : _GEN_1715; // @[executor.scala 470:55]
  wire [7:0] _GEN_3252 = opcode_1 != 4'h0 ? _GEN_2408 : _GEN_1716; // @[executor.scala 470:55]
  wire [7:0] _GEN_3253 = opcode_1 != 4'h0 ? _GEN_2409 : _GEN_1717; // @[executor.scala 470:55]
  wire [7:0] _GEN_3254 = opcode_1 != 4'h0 ? _GEN_2414 : _GEN_1718; // @[executor.scala 470:55]
  wire [7:0] _GEN_3255 = opcode_1 != 4'h0 ? _GEN_2415 : _GEN_1719; // @[executor.scala 470:55]
  wire [7:0] _GEN_3256 = opcode_1 != 4'h0 ? _GEN_2416 : _GEN_1720; // @[executor.scala 470:55]
  wire [7:0] _GEN_3257 = opcode_1 != 4'h0 ? _GEN_2417 : _GEN_1721; // @[executor.scala 470:55]
  wire [7:0] _GEN_3258 = opcode_1 != 4'h0 ? _GEN_2422 : _GEN_1722; // @[executor.scala 470:55]
  wire [7:0] _GEN_3259 = opcode_1 != 4'h0 ? _GEN_2423 : _GEN_1723; // @[executor.scala 470:55]
  wire [7:0] _GEN_3260 = opcode_1 != 4'h0 ? _GEN_2424 : _GEN_1724; // @[executor.scala 470:55]
  wire [7:0] _GEN_3261 = opcode_1 != 4'h0 ? _GEN_2425 : _GEN_1725; // @[executor.scala 470:55]
  wire [7:0] _GEN_3262 = opcode_1 != 4'h0 ? _GEN_2430 : _GEN_1726; // @[executor.scala 470:55]
  wire [7:0] _GEN_3263 = opcode_1 != 4'h0 ? _GEN_2431 : _GEN_1727; // @[executor.scala 470:55]
  wire [7:0] _GEN_3264 = opcode_1 != 4'h0 ? _GEN_2432 : _GEN_1728; // @[executor.scala 470:55]
  wire [7:0] _GEN_3265 = opcode_1 != 4'h0 ? _GEN_2433 : _GEN_1729; // @[executor.scala 470:55]
  wire [7:0] _GEN_3266 = opcode_1 != 4'h0 ? _GEN_2438 : _GEN_1730; // @[executor.scala 470:55]
  wire [7:0] _GEN_3267 = opcode_1 != 4'h0 ? _GEN_2439 : _GEN_1731; // @[executor.scala 470:55]
  wire [7:0] _GEN_3268 = opcode_1 != 4'h0 ? _GEN_2440 : _GEN_1732; // @[executor.scala 470:55]
  wire [7:0] _GEN_3269 = opcode_1 != 4'h0 ? _GEN_2441 : _GEN_1733; // @[executor.scala 470:55]
  wire [7:0] _GEN_3270 = opcode_1 != 4'h0 ? _GEN_2446 : _GEN_1734; // @[executor.scala 470:55]
  wire [7:0] _GEN_3271 = opcode_1 != 4'h0 ? _GEN_2447 : _GEN_1735; // @[executor.scala 470:55]
  wire [7:0] _GEN_3272 = opcode_1 != 4'h0 ? _GEN_2448 : _GEN_1736; // @[executor.scala 470:55]
  wire [7:0] _GEN_3273 = opcode_1 != 4'h0 ? _GEN_2449 : _GEN_1737; // @[executor.scala 470:55]
  wire [7:0] _GEN_3274 = opcode_1 != 4'h0 ? _GEN_2454 : _GEN_1738; // @[executor.scala 470:55]
  wire [7:0] _GEN_3275 = opcode_1 != 4'h0 ? _GEN_2455 : _GEN_1739; // @[executor.scala 470:55]
  wire [7:0] _GEN_3276 = opcode_1 != 4'h0 ? _GEN_2456 : _GEN_1740; // @[executor.scala 470:55]
  wire [7:0] _GEN_3277 = opcode_1 != 4'h0 ? _GEN_2457 : _GEN_1741; // @[executor.scala 470:55]
  wire [7:0] _GEN_3278 = opcode_1 != 4'h0 ? _GEN_2462 : _GEN_1742; // @[executor.scala 470:55]
  wire [7:0] _GEN_3279 = opcode_1 != 4'h0 ? _GEN_2463 : _GEN_1743; // @[executor.scala 470:55]
  wire [7:0] _GEN_3280 = opcode_1 != 4'h0 ? _GEN_2464 : _GEN_1744; // @[executor.scala 470:55]
  wire [7:0] _GEN_3281 = opcode_1 != 4'h0 ? _GEN_2465 : _GEN_1745; // @[executor.scala 470:55]
  wire [7:0] _GEN_3282 = opcode_1 != 4'h0 ? _GEN_2470 : _GEN_1746; // @[executor.scala 470:55]
  wire [7:0] _GEN_3283 = opcode_1 != 4'h0 ? _GEN_2471 : _GEN_1747; // @[executor.scala 470:55]
  wire [7:0] _GEN_3284 = opcode_1 != 4'h0 ? _GEN_2472 : _GEN_1748; // @[executor.scala 470:55]
  wire [7:0] _GEN_3285 = opcode_1 != 4'h0 ? _GEN_2473 : _GEN_1749; // @[executor.scala 470:55]
  wire [7:0] _GEN_3286 = opcode_1 != 4'h0 ? _GEN_2478 : _GEN_1750; // @[executor.scala 470:55]
  wire [7:0] _GEN_3287 = opcode_1 != 4'h0 ? _GEN_2479 : _GEN_1751; // @[executor.scala 470:55]
  wire [7:0] _GEN_3288 = opcode_1 != 4'h0 ? _GEN_2480 : _GEN_1752; // @[executor.scala 470:55]
  wire [7:0] _GEN_3289 = opcode_1 != 4'h0 ? _GEN_2481 : _GEN_1753; // @[executor.scala 470:55]
  wire [7:0] _GEN_3290 = opcode_1 != 4'h0 ? _GEN_2486 : _GEN_1754; // @[executor.scala 470:55]
  wire [7:0] _GEN_3291 = opcode_1 != 4'h0 ? _GEN_2487 : _GEN_1755; // @[executor.scala 470:55]
  wire [7:0] _GEN_3292 = opcode_1 != 4'h0 ? _GEN_2488 : _GEN_1756; // @[executor.scala 470:55]
  wire [7:0] _GEN_3293 = opcode_1 != 4'h0 ? _GEN_2489 : _GEN_1757; // @[executor.scala 470:55]
  wire [7:0] _GEN_3294 = opcode_1 != 4'h0 ? _GEN_2494 : _GEN_1758; // @[executor.scala 470:55]
  wire [7:0] _GEN_3295 = opcode_1 != 4'h0 ? _GEN_2495 : _GEN_1759; // @[executor.scala 470:55]
  wire [7:0] _GEN_3296 = opcode_1 != 4'h0 ? _GEN_2496 : _GEN_1760; // @[executor.scala 470:55]
  wire [7:0] _GEN_3297 = opcode_1 != 4'h0 ? _GEN_2497 : _GEN_1761; // @[executor.scala 470:55]
  wire [7:0] _GEN_3298 = opcode_1 != 4'h0 ? _GEN_2502 : _GEN_1762; // @[executor.scala 470:55]
  wire [7:0] _GEN_3299 = opcode_1 != 4'h0 ? _GEN_2503 : _GEN_1763; // @[executor.scala 470:55]
  wire [7:0] _GEN_3300 = opcode_1 != 4'h0 ? _GEN_2504 : _GEN_1764; // @[executor.scala 470:55]
  wire [7:0] _GEN_3301 = opcode_1 != 4'h0 ? _GEN_2505 : _GEN_1765; // @[executor.scala 470:55]
  wire [7:0] _GEN_3302 = opcode_1 != 4'h0 ? _GEN_2510 : _GEN_1766; // @[executor.scala 470:55]
  wire [7:0] _GEN_3303 = opcode_1 != 4'h0 ? _GEN_2511 : _GEN_1767; // @[executor.scala 470:55]
  wire [7:0] _GEN_3304 = opcode_1 != 4'h0 ? _GEN_2512 : _GEN_1768; // @[executor.scala 470:55]
  wire [7:0] _GEN_3305 = opcode_1 != 4'h0 ? _GEN_2513 : _GEN_1769; // @[executor.scala 470:55]
  wire [7:0] _GEN_3306 = opcode_1 != 4'h0 ? _GEN_2518 : _GEN_1770; // @[executor.scala 470:55]
  wire [7:0] _GEN_3307 = opcode_1 != 4'h0 ? _GEN_2519 : _GEN_1771; // @[executor.scala 470:55]
  wire [7:0] _GEN_3308 = opcode_1 != 4'h0 ? _GEN_2520 : _GEN_1772; // @[executor.scala 470:55]
  wire [7:0] _GEN_3309 = opcode_1 != 4'h0 ? _GEN_2521 : _GEN_1773; // @[executor.scala 470:55]
  wire [7:0] _GEN_3310 = opcode_1 != 4'h0 ? _GEN_2526 : _GEN_1774; // @[executor.scala 470:55]
  wire [7:0] _GEN_3311 = opcode_1 != 4'h0 ? _GEN_2527 : _GEN_1775; // @[executor.scala 470:55]
  wire [7:0] _GEN_3312 = opcode_1 != 4'h0 ? _GEN_2528 : _GEN_1776; // @[executor.scala 470:55]
  wire [7:0] _GEN_3313 = opcode_1 != 4'h0 ? _GEN_2529 : _GEN_1777; // @[executor.scala 470:55]
  wire [7:0] _GEN_3314 = opcode_1 != 4'h0 ? _GEN_2534 : _GEN_1778; // @[executor.scala 470:55]
  wire [7:0] _GEN_3315 = opcode_1 != 4'h0 ? _GEN_2535 : _GEN_1779; // @[executor.scala 470:55]
  wire [7:0] _GEN_3316 = opcode_1 != 4'h0 ? _GEN_2536 : _GEN_1780; // @[executor.scala 470:55]
  wire [7:0] _GEN_3317 = opcode_1 != 4'h0 ? _GEN_2537 : _GEN_1781; // @[executor.scala 470:55]
  wire [7:0] _GEN_3318 = opcode_1 != 4'h0 ? _GEN_2542 : _GEN_1782; // @[executor.scala 470:55]
  wire [7:0] _GEN_3319 = opcode_1 != 4'h0 ? _GEN_2543 : _GEN_1783; // @[executor.scala 470:55]
  wire [7:0] _GEN_3320 = opcode_1 != 4'h0 ? _GEN_2544 : _GEN_1784; // @[executor.scala 470:55]
  wire [7:0] _GEN_3321 = opcode_1 != 4'h0 ? _GEN_2545 : _GEN_1785; // @[executor.scala 470:55]
  wire [7:0] _GEN_3322 = opcode_1 != 4'h0 ? _GEN_2550 : _GEN_1786; // @[executor.scala 470:55]
  wire [7:0] _GEN_3323 = opcode_1 != 4'h0 ? _GEN_2551 : _GEN_1787; // @[executor.scala 470:55]
  wire [7:0] _GEN_3324 = opcode_1 != 4'h0 ? _GEN_2552 : _GEN_1788; // @[executor.scala 470:55]
  wire [7:0] _GEN_3325 = opcode_1 != 4'h0 ? _GEN_2553 : _GEN_1789; // @[executor.scala 470:55]
  wire [7:0] _GEN_3326 = opcode_1 != 4'h0 ? _GEN_2558 : _GEN_1790; // @[executor.scala 470:55]
  wire [7:0] _GEN_3327 = opcode_1 != 4'h0 ? _GEN_2559 : _GEN_1791; // @[executor.scala 470:55]
  wire [7:0] _GEN_3328 = opcode_1 != 4'h0 ? _GEN_2560 : _GEN_1792; // @[executor.scala 470:55]
  wire [7:0] _GEN_3329 = opcode_1 != 4'h0 ? _GEN_2561 : _GEN_1793; // @[executor.scala 470:55]
  wire [7:0] _GEN_3330 = opcode_1 != 4'h0 ? _GEN_2566 : _GEN_1794; // @[executor.scala 470:55]
  wire [7:0] _GEN_3331 = opcode_1 != 4'h0 ? _GEN_2567 : _GEN_1795; // @[executor.scala 470:55]
  wire [7:0] _GEN_3332 = opcode_1 != 4'h0 ? _GEN_2568 : _GEN_1796; // @[executor.scala 470:55]
  wire [7:0] _GEN_3333 = opcode_1 != 4'h0 ? _GEN_2569 : _GEN_1797; // @[executor.scala 470:55]
  wire [7:0] _GEN_3334 = opcode_1 != 4'h0 ? _GEN_2574 : _GEN_1798; // @[executor.scala 470:55]
  wire [7:0] _GEN_3335 = opcode_1 != 4'h0 ? _GEN_2575 : _GEN_1799; // @[executor.scala 470:55]
  wire [7:0] _GEN_3336 = opcode_1 != 4'h0 ? _GEN_2576 : _GEN_1800; // @[executor.scala 470:55]
  wire [7:0] _GEN_3337 = opcode_1 != 4'h0 ? _GEN_2577 : _GEN_1801; // @[executor.scala 470:55]
  wire [7:0] _GEN_3338 = opcode_1 != 4'h0 ? _GEN_2582 : _GEN_1802; // @[executor.scala 470:55]
  wire [7:0] _GEN_3339 = opcode_1 != 4'h0 ? _GEN_2583 : _GEN_1803; // @[executor.scala 470:55]
  wire [7:0] _GEN_3340 = opcode_1 != 4'h0 ? _GEN_2584 : _GEN_1804; // @[executor.scala 470:55]
  wire [7:0] _GEN_3341 = opcode_1 != 4'h0 ? _GEN_2585 : _GEN_1805; // @[executor.scala 470:55]
  wire [7:0] _GEN_3342 = opcode_1 != 4'h0 ? _GEN_2590 : _GEN_1806; // @[executor.scala 470:55]
  wire [7:0] _GEN_3343 = opcode_1 != 4'h0 ? _GEN_2591 : _GEN_1807; // @[executor.scala 470:55]
  wire [7:0] _GEN_3344 = opcode_1 != 4'h0 ? _GEN_2592 : _GEN_1808; // @[executor.scala 470:55]
  wire [7:0] _GEN_3345 = opcode_1 != 4'h0 ? _GEN_2593 : _GEN_1809; // @[executor.scala 470:55]
  wire [7:0] _GEN_3346 = opcode_1 != 4'h0 ? _GEN_2598 : _GEN_1810; // @[executor.scala 470:55]
  wire [7:0] _GEN_3347 = opcode_1 != 4'h0 ? _GEN_2599 : _GEN_1811; // @[executor.scala 470:55]
  wire [7:0] _GEN_3348 = opcode_1 != 4'h0 ? _GEN_2600 : _GEN_1812; // @[executor.scala 470:55]
  wire [7:0] _GEN_3349 = opcode_1 != 4'h0 ? _GEN_2601 : _GEN_1813; // @[executor.scala 470:55]
  wire [7:0] _GEN_3350 = opcode_1 != 4'h0 ? _GEN_2606 : _GEN_1814; // @[executor.scala 470:55]
  wire [7:0] _GEN_3351 = opcode_1 != 4'h0 ? _GEN_2607 : _GEN_1815; // @[executor.scala 470:55]
  wire [7:0] _GEN_3352 = opcode_1 != 4'h0 ? _GEN_2608 : _GEN_1816; // @[executor.scala 470:55]
  wire [7:0] _GEN_3353 = opcode_1 != 4'h0 ? _GEN_2609 : _GEN_1817; // @[executor.scala 470:55]
  wire [7:0] _GEN_3354 = opcode_1 != 4'h0 ? _GEN_2614 : _GEN_1818; // @[executor.scala 470:55]
  wire [7:0] _GEN_3355 = opcode_1 != 4'h0 ? _GEN_2615 : _GEN_1819; // @[executor.scala 470:55]
  wire [7:0] _GEN_3356 = opcode_1 != 4'h0 ? _GEN_2616 : _GEN_1820; // @[executor.scala 470:55]
  wire [7:0] _GEN_3357 = opcode_1 != 4'h0 ? _GEN_2617 : _GEN_1821; // @[executor.scala 470:55]
  wire [7:0] _GEN_3358 = opcode_1 != 4'h0 ? _GEN_2622 : _GEN_1822; // @[executor.scala 470:55]
  wire [7:0] _GEN_3359 = opcode_1 != 4'h0 ? _GEN_2623 : _GEN_1823; // @[executor.scala 470:55]
  wire [7:0] _GEN_3360 = opcode_1 != 4'h0 ? _GEN_2624 : _GEN_1824; // @[executor.scala 470:55]
  wire [7:0] _GEN_3361 = opcode_1 != 4'h0 ? _GEN_2625 : _GEN_1825; // @[executor.scala 470:55]
  wire [7:0] _GEN_3362 = opcode_1 != 4'h0 ? _GEN_2630 : _GEN_1826; // @[executor.scala 470:55]
  wire [7:0] _GEN_3363 = opcode_1 != 4'h0 ? _GEN_2631 : _GEN_1827; // @[executor.scala 470:55]
  wire [7:0] _GEN_3364 = opcode_1 != 4'h0 ? _GEN_2632 : _GEN_1828; // @[executor.scala 470:55]
  wire [7:0] _GEN_3365 = opcode_1 != 4'h0 ? _GEN_2633 : _GEN_1829; // @[executor.scala 470:55]
  wire [7:0] _GEN_3366 = opcode_1 != 4'h0 ? _GEN_2638 : _GEN_1830; // @[executor.scala 470:55]
  wire [7:0] _GEN_3367 = opcode_1 != 4'h0 ? _GEN_2639 : _GEN_1831; // @[executor.scala 470:55]
  wire [7:0] _GEN_3368 = opcode_1 != 4'h0 ? _GEN_2640 : _GEN_1832; // @[executor.scala 470:55]
  wire [7:0] _GEN_3369 = opcode_1 != 4'h0 ? _GEN_2641 : _GEN_1833; // @[executor.scala 470:55]
  wire [7:0] _GEN_3370 = opcode_1 != 4'h0 ? _GEN_2646 : _GEN_1834; // @[executor.scala 470:55]
  wire [7:0] _GEN_3371 = opcode_1 != 4'h0 ? _GEN_2647 : _GEN_1835; // @[executor.scala 470:55]
  wire [7:0] _GEN_3372 = opcode_1 != 4'h0 ? _GEN_2648 : _GEN_1836; // @[executor.scala 470:55]
  wire [7:0] _GEN_3373 = opcode_1 != 4'h0 ? _GEN_2649 : _GEN_1837; // @[executor.scala 470:55]
  wire [7:0] _GEN_3374 = opcode_1 != 4'h0 ? _GEN_2654 : _GEN_1838; // @[executor.scala 470:55]
  wire [7:0] _GEN_3375 = opcode_1 != 4'h0 ? _GEN_2655 : _GEN_1839; // @[executor.scala 470:55]
  wire [7:0] _GEN_3376 = opcode_1 != 4'h0 ? _GEN_2656 : _GEN_1840; // @[executor.scala 470:55]
  wire [7:0] _GEN_3377 = opcode_1 != 4'h0 ? _GEN_2657 : _GEN_1841; // @[executor.scala 470:55]
  wire [7:0] _GEN_3378 = opcode_1 != 4'h0 ? _GEN_2662 : _GEN_1842; // @[executor.scala 470:55]
  wire [7:0] _GEN_3379 = opcode_1 != 4'h0 ? _GEN_2663 : _GEN_1843; // @[executor.scala 470:55]
  wire [7:0] _GEN_3380 = opcode_1 != 4'h0 ? _GEN_2664 : _GEN_1844; // @[executor.scala 470:55]
  wire [7:0] _GEN_3381 = opcode_1 != 4'h0 ? _GEN_2665 : _GEN_1845; // @[executor.scala 470:55]
  wire [7:0] _GEN_3382 = opcode_1 != 4'h0 ? _GEN_2670 : _GEN_1846; // @[executor.scala 470:55]
  wire [7:0] _GEN_3383 = opcode_1 != 4'h0 ? _GEN_2671 : _GEN_1847; // @[executor.scala 470:55]
  wire [7:0] _GEN_3384 = opcode_1 != 4'h0 ? _GEN_2672 : _GEN_1848; // @[executor.scala 470:55]
  wire [7:0] _GEN_3385 = opcode_1 != 4'h0 ? _GEN_2673 : _GEN_1849; // @[executor.scala 470:55]
  wire [7:0] _GEN_3386 = opcode_1 != 4'h0 ? _GEN_2678 : _GEN_1850; // @[executor.scala 470:55]
  wire [7:0] _GEN_3387 = opcode_1 != 4'h0 ? _GEN_2679 : _GEN_1851; // @[executor.scala 470:55]
  wire [7:0] _GEN_3388 = opcode_1 != 4'h0 ? _GEN_2680 : _GEN_1852; // @[executor.scala 470:55]
  wire [7:0] _GEN_3389 = opcode_1 != 4'h0 ? _GEN_2681 : _GEN_1853; // @[executor.scala 470:55]
  wire [7:0] _GEN_3390 = opcode_1 != 4'h0 ? _GEN_2686 : _GEN_1854; // @[executor.scala 470:55]
  wire [7:0] _GEN_3391 = opcode_1 != 4'h0 ? _GEN_2687 : _GEN_1855; // @[executor.scala 470:55]
  wire [7:0] _GEN_3392 = opcode_1 != 4'h0 ? _GEN_2688 : _GEN_1856; // @[executor.scala 470:55]
  wire [7:0] _GEN_3393 = opcode_1 != 4'h0 ? _GEN_2689 : _GEN_1857; // @[executor.scala 470:55]
  wire [7:0] _GEN_3394 = opcode_1 != 4'h0 ? _GEN_2694 : _GEN_1858; // @[executor.scala 470:55]
  wire [7:0] _GEN_3395 = opcode_1 != 4'h0 ? _GEN_2695 : _GEN_1859; // @[executor.scala 470:55]
  wire [7:0] _GEN_3396 = opcode_1 != 4'h0 ? _GEN_2696 : _GEN_1860; // @[executor.scala 470:55]
  wire [7:0] _GEN_3397 = opcode_1 != 4'h0 ? _GEN_2697 : _GEN_1861; // @[executor.scala 470:55]
  wire [7:0] _GEN_3398 = opcode_1 != 4'h0 ? _GEN_2702 : _GEN_1862; // @[executor.scala 470:55]
  wire [7:0] _GEN_3399 = opcode_1 != 4'h0 ? _GEN_2703 : _GEN_1863; // @[executor.scala 470:55]
  wire [7:0] _GEN_3400 = opcode_1 != 4'h0 ? _GEN_2704 : _GEN_1864; // @[executor.scala 470:55]
  wire [7:0] _GEN_3401 = opcode_1 != 4'h0 ? _GEN_2705 : _GEN_1865; // @[executor.scala 470:55]
  wire [7:0] _GEN_3402 = opcode_1 != 4'h0 ? _GEN_2710 : _GEN_1866; // @[executor.scala 470:55]
  wire [7:0] _GEN_3403 = opcode_1 != 4'h0 ? _GEN_2711 : _GEN_1867; // @[executor.scala 470:55]
  wire [7:0] _GEN_3404 = opcode_1 != 4'h0 ? _GEN_2712 : _GEN_1868; // @[executor.scala 470:55]
  wire [7:0] _GEN_3405 = opcode_1 != 4'h0 ? _GEN_2713 : _GEN_1869; // @[executor.scala 470:55]
  wire [7:0] _GEN_3406 = opcode_1 != 4'h0 ? _GEN_2718 : _GEN_1870; // @[executor.scala 470:55]
  wire [7:0] _GEN_3407 = opcode_1 != 4'h0 ? _GEN_2719 : _GEN_1871; // @[executor.scala 470:55]
  wire [7:0] _GEN_3408 = opcode_1 != 4'h0 ? _GEN_2720 : _GEN_1872; // @[executor.scala 470:55]
  wire [7:0] _GEN_3409 = opcode_1 != 4'h0 ? _GEN_2721 : _GEN_1873; // @[executor.scala 470:55]
  wire [7:0] _GEN_3410 = opcode_1 != 4'h0 ? _GEN_2726 : _GEN_1874; // @[executor.scala 470:55]
  wire [7:0] _GEN_3411 = opcode_1 != 4'h0 ? _GEN_2727 : _GEN_1875; // @[executor.scala 470:55]
  wire [7:0] _GEN_3412 = opcode_1 != 4'h0 ? _GEN_2728 : _GEN_1876; // @[executor.scala 470:55]
  wire [7:0] _GEN_3413 = opcode_1 != 4'h0 ? _GEN_2729 : _GEN_1877; // @[executor.scala 470:55]
  wire [7:0] _GEN_3414 = opcode_1 != 4'h0 ? _GEN_2734 : _GEN_1878; // @[executor.scala 470:55]
  wire [7:0] _GEN_3415 = opcode_1 != 4'h0 ? _GEN_2735 : _GEN_1879; // @[executor.scala 470:55]
  wire [7:0] _GEN_3416 = opcode_1 != 4'h0 ? _GEN_2736 : _GEN_1880; // @[executor.scala 470:55]
  wire [7:0] _GEN_3417 = opcode_1 != 4'h0 ? _GEN_2737 : _GEN_1881; // @[executor.scala 470:55]
  wire [7:0] _GEN_3418 = opcode_1 != 4'h0 ? _GEN_2742 : _GEN_1882; // @[executor.scala 470:55]
  wire [7:0] _GEN_3419 = opcode_1 != 4'h0 ? _GEN_2743 : _GEN_1883; // @[executor.scala 470:55]
  wire [7:0] _GEN_3420 = opcode_1 != 4'h0 ? _GEN_2744 : _GEN_1884; // @[executor.scala 470:55]
  wire [7:0] _GEN_3421 = opcode_1 != 4'h0 ? _GEN_2745 : _GEN_1885; // @[executor.scala 470:55]
  wire [7:0] _GEN_3422 = opcode_1 != 4'h0 ? _GEN_2750 : _GEN_1886; // @[executor.scala 470:55]
  wire [7:0] _GEN_3423 = opcode_1 != 4'h0 ? _GEN_2751 : _GEN_1887; // @[executor.scala 470:55]
  wire [7:0] _GEN_3424 = opcode_1 != 4'h0 ? _GEN_2752 : _GEN_1888; // @[executor.scala 470:55]
  wire [7:0] _GEN_3425 = opcode_1 != 4'h0 ? _GEN_2753 : _GEN_1889; // @[executor.scala 470:55]
  wire [7:0] _GEN_3426 = opcode_1 != 4'h0 ? _GEN_2758 : _GEN_1890; // @[executor.scala 470:55]
  wire [7:0] _GEN_3427 = opcode_1 != 4'h0 ? _GEN_2759 : _GEN_1891; // @[executor.scala 470:55]
  wire [7:0] _GEN_3428 = opcode_1 != 4'h0 ? _GEN_2760 : _GEN_1892; // @[executor.scala 470:55]
  wire [7:0] _GEN_3429 = opcode_1 != 4'h0 ? _GEN_2761 : _GEN_1893; // @[executor.scala 470:55]
  wire [7:0] _GEN_3430 = opcode_1 != 4'h0 ? _GEN_2766 : _GEN_1894; // @[executor.scala 470:55]
  wire [7:0] _GEN_3431 = opcode_1 != 4'h0 ? _GEN_2767 : _GEN_1895; // @[executor.scala 470:55]
  wire [7:0] _GEN_3432 = opcode_1 != 4'h0 ? _GEN_2768 : _GEN_1896; // @[executor.scala 470:55]
  wire [7:0] _GEN_3433 = opcode_1 != 4'h0 ? _GEN_2769 : _GEN_1897; // @[executor.scala 470:55]
  wire [7:0] _GEN_3434 = opcode_1 != 4'h0 ? _GEN_2774 : _GEN_1898; // @[executor.scala 470:55]
  wire [7:0] _GEN_3435 = opcode_1 != 4'h0 ? _GEN_2775 : _GEN_1899; // @[executor.scala 470:55]
  wire [7:0] _GEN_3436 = opcode_1 != 4'h0 ? _GEN_2776 : _GEN_1900; // @[executor.scala 470:55]
  wire [7:0] _GEN_3437 = opcode_1 != 4'h0 ? _GEN_2777 : _GEN_1901; // @[executor.scala 470:55]
  wire [7:0] _GEN_3438 = opcode_1 != 4'h0 ? _GEN_2782 : _GEN_1902; // @[executor.scala 470:55]
  wire [7:0] _GEN_3439 = opcode_1 != 4'h0 ? _GEN_2783 : _GEN_1903; // @[executor.scala 470:55]
  wire [7:0] _GEN_3440 = opcode_1 != 4'h0 ? _GEN_2784 : _GEN_1904; // @[executor.scala 470:55]
  wire [7:0] _GEN_3441 = opcode_1 != 4'h0 ? _GEN_2785 : _GEN_1905; // @[executor.scala 470:55]
  wire [7:0] _GEN_3442 = opcode_1 != 4'h0 ? _GEN_2790 : _GEN_1906; // @[executor.scala 470:55]
  wire [7:0] _GEN_3443 = opcode_1 != 4'h0 ? _GEN_2791 : _GEN_1907; // @[executor.scala 470:55]
  wire [7:0] _GEN_3444 = opcode_1 != 4'h0 ? _GEN_2792 : _GEN_1908; // @[executor.scala 470:55]
  wire [7:0] _GEN_3445 = opcode_1 != 4'h0 ? _GEN_2793 : _GEN_1909; // @[executor.scala 470:55]
  wire [7:0] _GEN_3446 = opcode_1 != 4'h0 ? _GEN_2798 : _GEN_1910; // @[executor.scala 470:55]
  wire [7:0] _GEN_3447 = opcode_1 != 4'h0 ? _GEN_2799 : _GEN_1911; // @[executor.scala 470:55]
  wire [7:0] _GEN_3448 = opcode_1 != 4'h0 ? _GEN_2800 : _GEN_1912; // @[executor.scala 470:55]
  wire [7:0] _GEN_3449 = opcode_1 != 4'h0 ? _GEN_2801 : _GEN_1913; // @[executor.scala 470:55]
  wire [7:0] _GEN_3450 = opcode_1 != 4'h0 ? _GEN_2806 : _GEN_1914; // @[executor.scala 470:55]
  wire [7:0] _GEN_3451 = opcode_1 != 4'h0 ? _GEN_2807 : _GEN_1915; // @[executor.scala 470:55]
  wire [7:0] _GEN_3452 = opcode_1 != 4'h0 ? _GEN_2808 : _GEN_1916; // @[executor.scala 470:55]
  wire [7:0] _GEN_3453 = opcode_1 != 4'h0 ? _GEN_2809 : _GEN_1917; // @[executor.scala 470:55]
  wire [7:0] _GEN_3454 = opcode_1 != 4'h0 ? _GEN_2814 : _GEN_1918; // @[executor.scala 470:55]
  wire [7:0] _GEN_3455 = opcode_1 != 4'h0 ? _GEN_2815 : _GEN_1919; // @[executor.scala 470:55]
  wire [7:0] _GEN_3456 = opcode_1 != 4'h0 ? _GEN_2816 : _GEN_1920; // @[executor.scala 470:55]
  wire [7:0] _GEN_3457 = opcode_1 != 4'h0 ? _GEN_2817 : _GEN_1921; // @[executor.scala 470:55]
  wire [7:0] _GEN_3458 = opcode_1 != 4'h0 ? _GEN_2822 : _GEN_1922; // @[executor.scala 470:55]
  wire [7:0] _GEN_3459 = opcode_1 != 4'h0 ? _GEN_2823 : _GEN_1923; // @[executor.scala 470:55]
  wire [7:0] _GEN_3460 = opcode_1 != 4'h0 ? _GEN_2824 : _GEN_1924; // @[executor.scala 470:55]
  wire [7:0] _GEN_3461 = opcode_1 != 4'h0 ? _GEN_2825 : _GEN_1925; // @[executor.scala 470:55]
  wire [7:0] _GEN_3462 = opcode_1 != 4'h0 ? _GEN_2830 : _GEN_1926; // @[executor.scala 470:55]
  wire [7:0] _GEN_3463 = opcode_1 != 4'h0 ? _GEN_2831 : _GEN_1927; // @[executor.scala 470:55]
  wire [7:0] _GEN_3464 = opcode_1 != 4'h0 ? _GEN_2832 : _GEN_1928; // @[executor.scala 470:55]
  wire [7:0] _GEN_3465 = opcode_1 != 4'h0 ? _GEN_2833 : _GEN_1929; // @[executor.scala 470:55]
  wire [7:0] _GEN_3466 = opcode_1 != 4'h0 ? _GEN_2838 : _GEN_1930; // @[executor.scala 470:55]
  wire [7:0] _GEN_3467 = opcode_1 != 4'h0 ? _GEN_2839 : _GEN_1931; // @[executor.scala 470:55]
  wire [7:0] _GEN_3468 = opcode_1 != 4'h0 ? _GEN_2840 : _GEN_1932; // @[executor.scala 470:55]
  wire [7:0] _GEN_3469 = opcode_1 != 4'h0 ? _GEN_2841 : _GEN_1933; // @[executor.scala 470:55]
  wire [7:0] _GEN_3470 = opcode_1 != 4'h0 ? _GEN_2846 : _GEN_1934; // @[executor.scala 470:55]
  wire [7:0] _GEN_3471 = opcode_1 != 4'h0 ? _GEN_2847 : _GEN_1935; // @[executor.scala 470:55]
  wire [7:0] _GEN_3472 = opcode_1 != 4'h0 ? _GEN_2848 : _GEN_1936; // @[executor.scala 470:55]
  wire [7:0] _GEN_3473 = opcode_1 != 4'h0 ? _GEN_2849 : _GEN_1937; // @[executor.scala 470:55]
  wire [7:0] _GEN_3474 = opcode_1 != 4'h0 ? _GEN_2854 : _GEN_1938; // @[executor.scala 470:55]
  wire [7:0] _GEN_3475 = opcode_1 != 4'h0 ? _GEN_2855 : _GEN_1939; // @[executor.scala 470:55]
  wire [7:0] _GEN_3476 = opcode_1 != 4'h0 ? _GEN_2856 : _GEN_1940; // @[executor.scala 470:55]
  wire [7:0] _GEN_3477 = opcode_1 != 4'h0 ? _GEN_2857 : _GEN_1941; // @[executor.scala 470:55]
  wire [7:0] _GEN_3478 = opcode_1 != 4'h0 ? _GEN_2862 : _GEN_1942; // @[executor.scala 470:55]
  wire [7:0] _GEN_3479 = opcode_1 != 4'h0 ? _GEN_2863 : _GEN_1943; // @[executor.scala 470:55]
  wire [7:0] _GEN_3480 = opcode_1 != 4'h0 ? _GEN_2864 : _GEN_1944; // @[executor.scala 470:55]
  wire [7:0] _GEN_3481 = opcode_1 != 4'h0 ? _GEN_2865 : _GEN_1945; // @[executor.scala 470:55]
  wire [7:0] _GEN_3482 = opcode_1 != 4'h0 ? _GEN_2870 : _GEN_1946; // @[executor.scala 470:55]
  wire [7:0] _GEN_3483 = opcode_1 != 4'h0 ? _GEN_2871 : _GEN_1947; // @[executor.scala 470:55]
  wire [7:0] _GEN_3484 = opcode_1 != 4'h0 ? _GEN_2872 : _GEN_1948; // @[executor.scala 470:55]
  wire [7:0] _GEN_3485 = opcode_1 != 4'h0 ? _GEN_2873 : _GEN_1949; // @[executor.scala 470:55]
  wire [7:0] _GEN_3486 = opcode_1 != 4'h0 ? _GEN_2878 : _GEN_1950; // @[executor.scala 470:55]
  wire [7:0] _GEN_3487 = opcode_1 != 4'h0 ? _GEN_2879 : _GEN_1951; // @[executor.scala 470:55]
  wire [7:0] _GEN_3488 = opcode_1 != 4'h0 ? _GEN_2880 : _GEN_1952; // @[executor.scala 470:55]
  wire [7:0] _GEN_3489 = opcode_1 != 4'h0 ? _GEN_2881 : _GEN_1953; // @[executor.scala 470:55]
  wire [7:0] _GEN_3490 = opcode_1 != 4'h0 ? _GEN_2886 : _GEN_1954; // @[executor.scala 470:55]
  wire [7:0] _GEN_3491 = opcode_1 != 4'h0 ? _GEN_2887 : _GEN_1955; // @[executor.scala 470:55]
  wire [7:0] _GEN_3492 = opcode_1 != 4'h0 ? _GEN_2888 : _GEN_1956; // @[executor.scala 470:55]
  wire [7:0] _GEN_3493 = opcode_1 != 4'h0 ? _GEN_2889 : _GEN_1957; // @[executor.scala 470:55]
  wire [7:0] _GEN_3494 = opcode_1 != 4'h0 ? _GEN_2894 : _GEN_1958; // @[executor.scala 470:55]
  wire [7:0] _GEN_3495 = opcode_1 != 4'h0 ? _GEN_2895 : _GEN_1959; // @[executor.scala 470:55]
  wire [7:0] _GEN_3496 = opcode_1 != 4'h0 ? _GEN_2896 : _GEN_1960; // @[executor.scala 470:55]
  wire [7:0] _GEN_3497 = opcode_1 != 4'h0 ? _GEN_2897 : _GEN_1961; // @[executor.scala 470:55]
  wire [7:0] _GEN_3498 = opcode_1 != 4'h0 ? _GEN_2902 : _GEN_1962; // @[executor.scala 470:55]
  wire [7:0] _GEN_3499 = opcode_1 != 4'h0 ? _GEN_2903 : _GEN_1963; // @[executor.scala 470:55]
  wire [7:0] _GEN_3500 = opcode_1 != 4'h0 ? _GEN_2904 : _GEN_1964; // @[executor.scala 470:55]
  wire [7:0] _GEN_3501 = opcode_1 != 4'h0 ? _GEN_2905 : _GEN_1965; // @[executor.scala 470:55]
  wire [7:0] _GEN_3502 = opcode_1 != 4'h0 ? _GEN_2910 : _GEN_1966; // @[executor.scala 470:55]
  wire [7:0] _GEN_3503 = opcode_1 != 4'h0 ? _GEN_2911 : _GEN_1967; // @[executor.scala 470:55]
  wire [7:0] _GEN_3504 = opcode_1 != 4'h0 ? _GEN_2912 : _GEN_1968; // @[executor.scala 470:55]
  wire [7:0] _GEN_3505 = opcode_1 != 4'h0 ? _GEN_2913 : _GEN_1969; // @[executor.scala 470:55]
  wire [7:0] _GEN_3506 = opcode_1 != 4'h0 ? _GEN_2918 : _GEN_1970; // @[executor.scala 470:55]
  wire [7:0] _GEN_3507 = opcode_1 != 4'h0 ? _GEN_2919 : _GEN_1971; // @[executor.scala 470:55]
  wire [7:0] _GEN_3508 = opcode_1 != 4'h0 ? _GEN_2920 : _GEN_1972; // @[executor.scala 470:55]
  wire [7:0] _GEN_3509 = opcode_1 != 4'h0 ? _GEN_2921 : _GEN_1973; // @[executor.scala 470:55]
  wire [7:0] _GEN_3510 = opcode_1 != 4'h0 ? _GEN_2926 : _GEN_1974; // @[executor.scala 470:55]
  wire [7:0] _GEN_3511 = opcode_1 != 4'h0 ? _GEN_2927 : _GEN_1975; // @[executor.scala 470:55]
  wire [7:0] _GEN_3512 = opcode_1 != 4'h0 ? _GEN_2928 : _GEN_1976; // @[executor.scala 470:55]
  wire [7:0] _GEN_3513 = opcode_1 != 4'h0 ? _GEN_2929 : _GEN_1977; // @[executor.scala 470:55]
  wire [7:0] _GEN_3514 = opcode_1 != 4'h0 ? _GEN_2934 : _GEN_1978; // @[executor.scala 470:55]
  wire [7:0] _GEN_3515 = opcode_1 != 4'h0 ? _GEN_2935 : _GEN_1979; // @[executor.scala 470:55]
  wire [7:0] _GEN_3516 = opcode_1 != 4'h0 ? _GEN_2936 : _GEN_1980; // @[executor.scala 470:55]
  wire [7:0] _GEN_3517 = opcode_1 != 4'h0 ? _GEN_2937 : _GEN_1981; // @[executor.scala 470:55]
  wire [7:0] _GEN_3518 = opcode_1 != 4'h0 ? _GEN_2942 : _GEN_1982; // @[executor.scala 470:55]
  wire [7:0] _GEN_3519 = opcode_1 != 4'h0 ? _GEN_2943 : _GEN_1983; // @[executor.scala 470:55]
  wire [7:0] _GEN_3520 = opcode_1 != 4'h0 ? _GEN_2944 : _GEN_1984; // @[executor.scala 470:55]
  wire [7:0] _GEN_3521 = opcode_1 != 4'h0 ? _GEN_2945 : _GEN_1985; // @[executor.scala 470:55]
  wire [7:0] _GEN_3522 = opcode_1 != 4'h0 ? _GEN_2950 : _GEN_1986; // @[executor.scala 470:55]
  wire [7:0] _GEN_3523 = opcode_1 != 4'h0 ? _GEN_2951 : _GEN_1987; // @[executor.scala 470:55]
  wire [7:0] _GEN_3524 = opcode_1 != 4'h0 ? _GEN_2952 : _GEN_1988; // @[executor.scala 470:55]
  wire [7:0] _GEN_3525 = opcode_1 != 4'h0 ? _GEN_2953 : _GEN_1989; // @[executor.scala 470:55]
  wire [7:0] _GEN_3526 = opcode_1 != 4'h0 ? _GEN_2958 : _GEN_1990; // @[executor.scala 470:55]
  wire [7:0] _GEN_3527 = opcode_1 != 4'h0 ? _GEN_2959 : _GEN_1991; // @[executor.scala 470:55]
  wire [7:0] _GEN_3528 = opcode_1 != 4'h0 ? _GEN_2960 : _GEN_1992; // @[executor.scala 470:55]
  wire [7:0] _GEN_3529 = opcode_1 != 4'h0 ? _GEN_2961 : _GEN_1993; // @[executor.scala 470:55]
  wire [7:0] _GEN_3530 = opcode_1 != 4'h0 ? _GEN_2966 : _GEN_1994; // @[executor.scala 470:55]
  wire [7:0] _GEN_3531 = opcode_1 != 4'h0 ? _GEN_2967 : _GEN_1995; // @[executor.scala 470:55]
  wire [7:0] _GEN_3532 = opcode_1 != 4'h0 ? _GEN_2968 : _GEN_1996; // @[executor.scala 470:55]
  wire [7:0] _GEN_3533 = opcode_1 != 4'h0 ? _GEN_2969 : _GEN_1997; // @[executor.scala 470:55]
  wire [7:0] _GEN_3534 = opcode_1 != 4'h0 ? _GEN_2974 : _GEN_1998; // @[executor.scala 470:55]
  wire [7:0] _GEN_3535 = opcode_1 != 4'h0 ? _GEN_2975 : _GEN_1999; // @[executor.scala 470:55]
  wire [7:0] _GEN_3536 = opcode_1 != 4'h0 ? _GEN_2976 : _GEN_2000; // @[executor.scala 470:55]
  wire [7:0] _GEN_3537 = opcode_1 != 4'h0 ? _GEN_2977 : _GEN_2001; // @[executor.scala 470:55]
  wire [7:0] _GEN_3538 = opcode_1 != 4'h0 ? _GEN_2982 : _GEN_2002; // @[executor.scala 470:55]
  wire [7:0] _GEN_3539 = opcode_1 != 4'h0 ? _GEN_2983 : _GEN_2003; // @[executor.scala 470:55]
  wire [7:0] _GEN_3540 = opcode_1 != 4'h0 ? _GEN_2984 : _GEN_2004; // @[executor.scala 470:55]
  wire [7:0] _GEN_3541 = opcode_1 != 4'h0 ? _GEN_2985 : _GEN_2005; // @[executor.scala 470:55]
  wire [7:0] _GEN_3542 = opcode_1 != 4'h0 ? _GEN_2990 : _GEN_2006; // @[executor.scala 470:55]
  wire [7:0] _GEN_3543 = opcode_1 != 4'h0 ? _GEN_2991 : _GEN_2007; // @[executor.scala 470:55]
  wire [7:0] _GEN_3544 = opcode_1 != 4'h0 ? _GEN_2992 : _GEN_2008; // @[executor.scala 470:55]
  wire [7:0] _GEN_3545 = opcode_1 != 4'h0 ? _GEN_2993 : _GEN_2009; // @[executor.scala 470:55]
  wire [7:0] _GEN_3546 = opcode_1 != 4'h0 ? _GEN_2998 : _GEN_2010; // @[executor.scala 470:55]
  wire [7:0] _GEN_3547 = opcode_1 != 4'h0 ? _GEN_2999 : _GEN_2011; // @[executor.scala 470:55]
  wire [7:0] _GEN_3548 = opcode_1 != 4'h0 ? _GEN_3000 : _GEN_2012; // @[executor.scala 470:55]
  wire [7:0] _GEN_3549 = opcode_1 != 4'h0 ? _GEN_3001 : _GEN_2013; // @[executor.scala 470:55]
  wire [7:0] _GEN_3550 = opcode_1 != 4'h0 ? _GEN_3006 : _GEN_2014; // @[executor.scala 470:55]
  wire [7:0] _GEN_3551 = opcode_1 != 4'h0 ? _GEN_3007 : _GEN_2015; // @[executor.scala 470:55]
  wire [7:0] _GEN_3552 = opcode_1 != 4'h0 ? _GEN_3008 : _GEN_2016; // @[executor.scala 470:55]
  wire [7:0] _GEN_3553 = opcode_1 != 4'h0 ? _GEN_3009 : _GEN_2017; // @[executor.scala 470:55]
  wire [7:0] _GEN_3554 = opcode_1 != 4'h0 ? _GEN_3014 : _GEN_2018; // @[executor.scala 470:55]
  wire [7:0] _GEN_3555 = opcode_1 != 4'h0 ? _GEN_3015 : _GEN_2019; // @[executor.scala 470:55]
  wire [7:0] _GEN_3556 = opcode_1 != 4'h0 ? _GEN_3016 : _GEN_2020; // @[executor.scala 470:55]
  wire [7:0] _GEN_3557 = opcode_1 != 4'h0 ? _GEN_3017 : _GEN_2021; // @[executor.scala 470:55]
  wire [7:0] _GEN_3558 = opcode_1 != 4'h0 ? _GEN_3022 : _GEN_2022; // @[executor.scala 470:55]
  wire [7:0] _GEN_3559 = opcode_1 != 4'h0 ? _GEN_3023 : _GEN_2023; // @[executor.scala 470:55]
  wire [7:0] _GEN_3560 = opcode_1 != 4'h0 ? _GEN_3024 : _GEN_2024; // @[executor.scala 470:55]
  wire [7:0] _GEN_3561 = opcode_1 != 4'h0 ? _GEN_3025 : _GEN_2025; // @[executor.scala 470:55]
  wire [7:0] _GEN_3562 = opcode_1 != 4'h0 ? _GEN_3030 : _GEN_2026; // @[executor.scala 470:55]
  wire [7:0] _GEN_3563 = opcode_1 != 4'h0 ? _GEN_3031 : _GEN_2027; // @[executor.scala 470:55]
  wire [7:0] _GEN_3564 = opcode_1 != 4'h0 ? _GEN_3032 : _GEN_2028; // @[executor.scala 470:55]
  wire [7:0] _GEN_3565 = opcode_1 != 4'h0 ? _GEN_3033 : _GEN_2029; // @[executor.scala 470:55]
  wire [7:0] _GEN_3566 = opcode_1 != 4'h0 ? _GEN_3038 : _GEN_2030; // @[executor.scala 470:55]
  wire [7:0] _GEN_3567 = opcode_1 != 4'h0 ? _GEN_3039 : _GEN_2031; // @[executor.scala 470:55]
  wire [7:0] _GEN_3568 = opcode_1 != 4'h0 ? _GEN_3040 : _GEN_2032; // @[executor.scala 470:55]
  wire [7:0] _GEN_3569 = opcode_1 != 4'h0 ? _GEN_3041 : _GEN_2033; // @[executor.scala 470:55]
  wire [7:0] _GEN_3570 = opcode_1 != 4'h0 ? _GEN_3046 : _GEN_2034; // @[executor.scala 470:55]
  wire [7:0] _GEN_3571 = opcode_1 != 4'h0 ? _GEN_3047 : _GEN_2035; // @[executor.scala 470:55]
  wire [7:0] _GEN_3572 = opcode_1 != 4'h0 ? _GEN_3048 : _GEN_2036; // @[executor.scala 470:55]
  wire [7:0] _GEN_3573 = opcode_1 != 4'h0 ? _GEN_3049 : _GEN_2037; // @[executor.scala 470:55]
  wire [7:0] _GEN_3574 = opcode_1 != 4'h0 ? _GEN_3054 : _GEN_2038; // @[executor.scala 470:55]
  wire [7:0] _GEN_3575 = opcode_1 != 4'h0 ? _GEN_3055 : _GEN_2039; // @[executor.scala 470:55]
  wire [7:0] _GEN_3576 = opcode_1 != 4'h0 ? _GEN_3056 : _GEN_2040; // @[executor.scala 470:55]
  wire [7:0] _GEN_3577 = opcode_1 != 4'h0 ? _GEN_3057 : _GEN_2041; // @[executor.scala 470:55]
  wire [7:0] _GEN_3578 = opcode_1 != 4'h0 ? _GEN_3062 : _GEN_2042; // @[executor.scala 470:55]
  wire [7:0] _GEN_3579 = opcode_1 != 4'h0 ? _GEN_3063 : _GEN_2043; // @[executor.scala 470:55]
  wire [7:0] _GEN_3580 = opcode_1 != 4'h0 ? _GEN_3064 : _GEN_2044; // @[executor.scala 470:55]
  wire [7:0] _GEN_3581 = opcode_1 != 4'h0 ? _GEN_3065 : _GEN_2045; // @[executor.scala 470:55]
  wire [7:0] _GEN_3582 = opcode_1 != 4'h0 ? _GEN_3070 : _GEN_2046; // @[executor.scala 470:55]
  wire [7:0] _GEN_3583 = opcode_1 != 4'h0 ? _GEN_3071 : _GEN_2047; // @[executor.scala 470:55]
  wire [7:0] _GEN_3584 = opcode_1 != 4'h0 ? _GEN_3072 : _GEN_2048; // @[executor.scala 470:55]
  wire [7:0] _GEN_3585 = opcode_1 != 4'h0 ? _GEN_3073 : _GEN_2049; // @[executor.scala 470:55]
  wire [3:0] _GEN_3586 = opcode_1 == 4'hf ? parameter_2_1[13:10] : _GEN_1536; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_3587 = opcode_1 == 4'hf ? parameter_2_1[0] : _GEN_1537; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_3588 = opcode_1 == 4'hf ? _GEN_1538 : _GEN_3074; // @[executor.scala 466:52]
  wire [7:0] _GEN_3589 = opcode_1 == 4'hf ? _GEN_1539 : _GEN_3075; // @[executor.scala 466:52]
  wire [7:0] _GEN_3590 = opcode_1 == 4'hf ? _GEN_1540 : _GEN_3076; // @[executor.scala 466:52]
  wire [7:0] _GEN_3591 = opcode_1 == 4'hf ? _GEN_1541 : _GEN_3077; // @[executor.scala 466:52]
  wire [7:0] _GEN_3592 = opcode_1 == 4'hf ? _GEN_1542 : _GEN_3078; // @[executor.scala 466:52]
  wire [7:0] _GEN_3593 = opcode_1 == 4'hf ? _GEN_1543 : _GEN_3079; // @[executor.scala 466:52]
  wire [7:0] _GEN_3594 = opcode_1 == 4'hf ? _GEN_1544 : _GEN_3080; // @[executor.scala 466:52]
  wire [7:0] _GEN_3595 = opcode_1 == 4'hf ? _GEN_1545 : _GEN_3081; // @[executor.scala 466:52]
  wire [7:0] _GEN_3596 = opcode_1 == 4'hf ? _GEN_1546 : _GEN_3082; // @[executor.scala 466:52]
  wire [7:0] _GEN_3597 = opcode_1 == 4'hf ? _GEN_1547 : _GEN_3083; // @[executor.scala 466:52]
  wire [7:0] _GEN_3598 = opcode_1 == 4'hf ? _GEN_1548 : _GEN_3084; // @[executor.scala 466:52]
  wire [7:0] _GEN_3599 = opcode_1 == 4'hf ? _GEN_1549 : _GEN_3085; // @[executor.scala 466:52]
  wire [7:0] _GEN_3600 = opcode_1 == 4'hf ? _GEN_1550 : _GEN_3086; // @[executor.scala 466:52]
  wire [7:0] _GEN_3601 = opcode_1 == 4'hf ? _GEN_1551 : _GEN_3087; // @[executor.scala 466:52]
  wire [7:0] _GEN_3602 = opcode_1 == 4'hf ? _GEN_1552 : _GEN_3088; // @[executor.scala 466:52]
  wire [7:0] _GEN_3603 = opcode_1 == 4'hf ? _GEN_1553 : _GEN_3089; // @[executor.scala 466:52]
  wire [7:0] _GEN_3604 = opcode_1 == 4'hf ? _GEN_1554 : _GEN_3090; // @[executor.scala 466:52]
  wire [7:0] _GEN_3605 = opcode_1 == 4'hf ? _GEN_1555 : _GEN_3091; // @[executor.scala 466:52]
  wire [7:0] _GEN_3606 = opcode_1 == 4'hf ? _GEN_1556 : _GEN_3092; // @[executor.scala 466:52]
  wire [7:0] _GEN_3607 = opcode_1 == 4'hf ? _GEN_1557 : _GEN_3093; // @[executor.scala 466:52]
  wire [7:0] _GEN_3608 = opcode_1 == 4'hf ? _GEN_1558 : _GEN_3094; // @[executor.scala 466:52]
  wire [7:0] _GEN_3609 = opcode_1 == 4'hf ? _GEN_1559 : _GEN_3095; // @[executor.scala 466:52]
  wire [7:0] _GEN_3610 = opcode_1 == 4'hf ? _GEN_1560 : _GEN_3096; // @[executor.scala 466:52]
  wire [7:0] _GEN_3611 = opcode_1 == 4'hf ? _GEN_1561 : _GEN_3097; // @[executor.scala 466:52]
  wire [7:0] _GEN_3612 = opcode_1 == 4'hf ? _GEN_1562 : _GEN_3098; // @[executor.scala 466:52]
  wire [7:0] _GEN_3613 = opcode_1 == 4'hf ? _GEN_1563 : _GEN_3099; // @[executor.scala 466:52]
  wire [7:0] _GEN_3614 = opcode_1 == 4'hf ? _GEN_1564 : _GEN_3100; // @[executor.scala 466:52]
  wire [7:0] _GEN_3615 = opcode_1 == 4'hf ? _GEN_1565 : _GEN_3101; // @[executor.scala 466:52]
  wire [7:0] _GEN_3616 = opcode_1 == 4'hf ? _GEN_1566 : _GEN_3102; // @[executor.scala 466:52]
  wire [7:0] _GEN_3617 = opcode_1 == 4'hf ? _GEN_1567 : _GEN_3103; // @[executor.scala 466:52]
  wire [7:0] _GEN_3618 = opcode_1 == 4'hf ? _GEN_1568 : _GEN_3104; // @[executor.scala 466:52]
  wire [7:0] _GEN_3619 = opcode_1 == 4'hf ? _GEN_1569 : _GEN_3105; // @[executor.scala 466:52]
  wire [7:0] _GEN_3620 = opcode_1 == 4'hf ? _GEN_1570 : _GEN_3106; // @[executor.scala 466:52]
  wire [7:0] _GEN_3621 = opcode_1 == 4'hf ? _GEN_1571 : _GEN_3107; // @[executor.scala 466:52]
  wire [7:0] _GEN_3622 = opcode_1 == 4'hf ? _GEN_1572 : _GEN_3108; // @[executor.scala 466:52]
  wire [7:0] _GEN_3623 = opcode_1 == 4'hf ? _GEN_1573 : _GEN_3109; // @[executor.scala 466:52]
  wire [7:0] _GEN_3624 = opcode_1 == 4'hf ? _GEN_1574 : _GEN_3110; // @[executor.scala 466:52]
  wire [7:0] _GEN_3625 = opcode_1 == 4'hf ? _GEN_1575 : _GEN_3111; // @[executor.scala 466:52]
  wire [7:0] _GEN_3626 = opcode_1 == 4'hf ? _GEN_1576 : _GEN_3112; // @[executor.scala 466:52]
  wire [7:0] _GEN_3627 = opcode_1 == 4'hf ? _GEN_1577 : _GEN_3113; // @[executor.scala 466:52]
  wire [7:0] _GEN_3628 = opcode_1 == 4'hf ? _GEN_1578 : _GEN_3114; // @[executor.scala 466:52]
  wire [7:0] _GEN_3629 = opcode_1 == 4'hf ? _GEN_1579 : _GEN_3115; // @[executor.scala 466:52]
  wire [7:0] _GEN_3630 = opcode_1 == 4'hf ? _GEN_1580 : _GEN_3116; // @[executor.scala 466:52]
  wire [7:0] _GEN_3631 = opcode_1 == 4'hf ? _GEN_1581 : _GEN_3117; // @[executor.scala 466:52]
  wire [7:0] _GEN_3632 = opcode_1 == 4'hf ? _GEN_1582 : _GEN_3118; // @[executor.scala 466:52]
  wire [7:0] _GEN_3633 = opcode_1 == 4'hf ? _GEN_1583 : _GEN_3119; // @[executor.scala 466:52]
  wire [7:0] _GEN_3634 = opcode_1 == 4'hf ? _GEN_1584 : _GEN_3120; // @[executor.scala 466:52]
  wire [7:0] _GEN_3635 = opcode_1 == 4'hf ? _GEN_1585 : _GEN_3121; // @[executor.scala 466:52]
  wire [7:0] _GEN_3636 = opcode_1 == 4'hf ? _GEN_1586 : _GEN_3122; // @[executor.scala 466:52]
  wire [7:0] _GEN_3637 = opcode_1 == 4'hf ? _GEN_1587 : _GEN_3123; // @[executor.scala 466:52]
  wire [7:0] _GEN_3638 = opcode_1 == 4'hf ? _GEN_1588 : _GEN_3124; // @[executor.scala 466:52]
  wire [7:0] _GEN_3639 = opcode_1 == 4'hf ? _GEN_1589 : _GEN_3125; // @[executor.scala 466:52]
  wire [7:0] _GEN_3640 = opcode_1 == 4'hf ? _GEN_1590 : _GEN_3126; // @[executor.scala 466:52]
  wire [7:0] _GEN_3641 = opcode_1 == 4'hf ? _GEN_1591 : _GEN_3127; // @[executor.scala 466:52]
  wire [7:0] _GEN_3642 = opcode_1 == 4'hf ? _GEN_1592 : _GEN_3128; // @[executor.scala 466:52]
  wire [7:0] _GEN_3643 = opcode_1 == 4'hf ? _GEN_1593 : _GEN_3129; // @[executor.scala 466:52]
  wire [7:0] _GEN_3644 = opcode_1 == 4'hf ? _GEN_1594 : _GEN_3130; // @[executor.scala 466:52]
  wire [7:0] _GEN_3645 = opcode_1 == 4'hf ? _GEN_1595 : _GEN_3131; // @[executor.scala 466:52]
  wire [7:0] _GEN_3646 = opcode_1 == 4'hf ? _GEN_1596 : _GEN_3132; // @[executor.scala 466:52]
  wire [7:0] _GEN_3647 = opcode_1 == 4'hf ? _GEN_1597 : _GEN_3133; // @[executor.scala 466:52]
  wire [7:0] _GEN_3648 = opcode_1 == 4'hf ? _GEN_1598 : _GEN_3134; // @[executor.scala 466:52]
  wire [7:0] _GEN_3649 = opcode_1 == 4'hf ? _GEN_1599 : _GEN_3135; // @[executor.scala 466:52]
  wire [7:0] _GEN_3650 = opcode_1 == 4'hf ? _GEN_1600 : _GEN_3136; // @[executor.scala 466:52]
  wire [7:0] _GEN_3651 = opcode_1 == 4'hf ? _GEN_1601 : _GEN_3137; // @[executor.scala 466:52]
  wire [7:0] _GEN_3652 = opcode_1 == 4'hf ? _GEN_1602 : _GEN_3138; // @[executor.scala 466:52]
  wire [7:0] _GEN_3653 = opcode_1 == 4'hf ? _GEN_1603 : _GEN_3139; // @[executor.scala 466:52]
  wire [7:0] _GEN_3654 = opcode_1 == 4'hf ? _GEN_1604 : _GEN_3140; // @[executor.scala 466:52]
  wire [7:0] _GEN_3655 = opcode_1 == 4'hf ? _GEN_1605 : _GEN_3141; // @[executor.scala 466:52]
  wire [7:0] _GEN_3656 = opcode_1 == 4'hf ? _GEN_1606 : _GEN_3142; // @[executor.scala 466:52]
  wire [7:0] _GEN_3657 = opcode_1 == 4'hf ? _GEN_1607 : _GEN_3143; // @[executor.scala 466:52]
  wire [7:0] _GEN_3658 = opcode_1 == 4'hf ? _GEN_1608 : _GEN_3144; // @[executor.scala 466:52]
  wire [7:0] _GEN_3659 = opcode_1 == 4'hf ? _GEN_1609 : _GEN_3145; // @[executor.scala 466:52]
  wire [7:0] _GEN_3660 = opcode_1 == 4'hf ? _GEN_1610 : _GEN_3146; // @[executor.scala 466:52]
  wire [7:0] _GEN_3661 = opcode_1 == 4'hf ? _GEN_1611 : _GEN_3147; // @[executor.scala 466:52]
  wire [7:0] _GEN_3662 = opcode_1 == 4'hf ? _GEN_1612 : _GEN_3148; // @[executor.scala 466:52]
  wire [7:0] _GEN_3663 = opcode_1 == 4'hf ? _GEN_1613 : _GEN_3149; // @[executor.scala 466:52]
  wire [7:0] _GEN_3664 = opcode_1 == 4'hf ? _GEN_1614 : _GEN_3150; // @[executor.scala 466:52]
  wire [7:0] _GEN_3665 = opcode_1 == 4'hf ? _GEN_1615 : _GEN_3151; // @[executor.scala 466:52]
  wire [7:0] _GEN_3666 = opcode_1 == 4'hf ? _GEN_1616 : _GEN_3152; // @[executor.scala 466:52]
  wire [7:0] _GEN_3667 = opcode_1 == 4'hf ? _GEN_1617 : _GEN_3153; // @[executor.scala 466:52]
  wire [7:0] _GEN_3668 = opcode_1 == 4'hf ? _GEN_1618 : _GEN_3154; // @[executor.scala 466:52]
  wire [7:0] _GEN_3669 = opcode_1 == 4'hf ? _GEN_1619 : _GEN_3155; // @[executor.scala 466:52]
  wire [7:0] _GEN_3670 = opcode_1 == 4'hf ? _GEN_1620 : _GEN_3156; // @[executor.scala 466:52]
  wire [7:0] _GEN_3671 = opcode_1 == 4'hf ? _GEN_1621 : _GEN_3157; // @[executor.scala 466:52]
  wire [7:0] _GEN_3672 = opcode_1 == 4'hf ? _GEN_1622 : _GEN_3158; // @[executor.scala 466:52]
  wire [7:0] _GEN_3673 = opcode_1 == 4'hf ? _GEN_1623 : _GEN_3159; // @[executor.scala 466:52]
  wire [7:0] _GEN_3674 = opcode_1 == 4'hf ? _GEN_1624 : _GEN_3160; // @[executor.scala 466:52]
  wire [7:0] _GEN_3675 = opcode_1 == 4'hf ? _GEN_1625 : _GEN_3161; // @[executor.scala 466:52]
  wire [7:0] _GEN_3676 = opcode_1 == 4'hf ? _GEN_1626 : _GEN_3162; // @[executor.scala 466:52]
  wire [7:0] _GEN_3677 = opcode_1 == 4'hf ? _GEN_1627 : _GEN_3163; // @[executor.scala 466:52]
  wire [7:0] _GEN_3678 = opcode_1 == 4'hf ? _GEN_1628 : _GEN_3164; // @[executor.scala 466:52]
  wire [7:0] _GEN_3679 = opcode_1 == 4'hf ? _GEN_1629 : _GEN_3165; // @[executor.scala 466:52]
  wire [7:0] _GEN_3680 = opcode_1 == 4'hf ? _GEN_1630 : _GEN_3166; // @[executor.scala 466:52]
  wire [7:0] _GEN_3681 = opcode_1 == 4'hf ? _GEN_1631 : _GEN_3167; // @[executor.scala 466:52]
  wire [7:0] _GEN_3682 = opcode_1 == 4'hf ? _GEN_1632 : _GEN_3168; // @[executor.scala 466:52]
  wire [7:0] _GEN_3683 = opcode_1 == 4'hf ? _GEN_1633 : _GEN_3169; // @[executor.scala 466:52]
  wire [7:0] _GEN_3684 = opcode_1 == 4'hf ? _GEN_1634 : _GEN_3170; // @[executor.scala 466:52]
  wire [7:0] _GEN_3685 = opcode_1 == 4'hf ? _GEN_1635 : _GEN_3171; // @[executor.scala 466:52]
  wire [7:0] _GEN_3686 = opcode_1 == 4'hf ? _GEN_1636 : _GEN_3172; // @[executor.scala 466:52]
  wire [7:0] _GEN_3687 = opcode_1 == 4'hf ? _GEN_1637 : _GEN_3173; // @[executor.scala 466:52]
  wire [7:0] _GEN_3688 = opcode_1 == 4'hf ? _GEN_1638 : _GEN_3174; // @[executor.scala 466:52]
  wire [7:0] _GEN_3689 = opcode_1 == 4'hf ? _GEN_1639 : _GEN_3175; // @[executor.scala 466:52]
  wire [7:0] _GEN_3690 = opcode_1 == 4'hf ? _GEN_1640 : _GEN_3176; // @[executor.scala 466:52]
  wire [7:0] _GEN_3691 = opcode_1 == 4'hf ? _GEN_1641 : _GEN_3177; // @[executor.scala 466:52]
  wire [7:0] _GEN_3692 = opcode_1 == 4'hf ? _GEN_1642 : _GEN_3178; // @[executor.scala 466:52]
  wire [7:0] _GEN_3693 = opcode_1 == 4'hf ? _GEN_1643 : _GEN_3179; // @[executor.scala 466:52]
  wire [7:0] _GEN_3694 = opcode_1 == 4'hf ? _GEN_1644 : _GEN_3180; // @[executor.scala 466:52]
  wire [7:0] _GEN_3695 = opcode_1 == 4'hf ? _GEN_1645 : _GEN_3181; // @[executor.scala 466:52]
  wire [7:0] _GEN_3696 = opcode_1 == 4'hf ? _GEN_1646 : _GEN_3182; // @[executor.scala 466:52]
  wire [7:0] _GEN_3697 = opcode_1 == 4'hf ? _GEN_1647 : _GEN_3183; // @[executor.scala 466:52]
  wire [7:0] _GEN_3698 = opcode_1 == 4'hf ? _GEN_1648 : _GEN_3184; // @[executor.scala 466:52]
  wire [7:0] _GEN_3699 = opcode_1 == 4'hf ? _GEN_1649 : _GEN_3185; // @[executor.scala 466:52]
  wire [7:0] _GEN_3700 = opcode_1 == 4'hf ? _GEN_1650 : _GEN_3186; // @[executor.scala 466:52]
  wire [7:0] _GEN_3701 = opcode_1 == 4'hf ? _GEN_1651 : _GEN_3187; // @[executor.scala 466:52]
  wire [7:0] _GEN_3702 = opcode_1 == 4'hf ? _GEN_1652 : _GEN_3188; // @[executor.scala 466:52]
  wire [7:0] _GEN_3703 = opcode_1 == 4'hf ? _GEN_1653 : _GEN_3189; // @[executor.scala 466:52]
  wire [7:0] _GEN_3704 = opcode_1 == 4'hf ? _GEN_1654 : _GEN_3190; // @[executor.scala 466:52]
  wire [7:0] _GEN_3705 = opcode_1 == 4'hf ? _GEN_1655 : _GEN_3191; // @[executor.scala 466:52]
  wire [7:0] _GEN_3706 = opcode_1 == 4'hf ? _GEN_1656 : _GEN_3192; // @[executor.scala 466:52]
  wire [7:0] _GEN_3707 = opcode_1 == 4'hf ? _GEN_1657 : _GEN_3193; // @[executor.scala 466:52]
  wire [7:0] _GEN_3708 = opcode_1 == 4'hf ? _GEN_1658 : _GEN_3194; // @[executor.scala 466:52]
  wire [7:0] _GEN_3709 = opcode_1 == 4'hf ? _GEN_1659 : _GEN_3195; // @[executor.scala 466:52]
  wire [7:0] _GEN_3710 = opcode_1 == 4'hf ? _GEN_1660 : _GEN_3196; // @[executor.scala 466:52]
  wire [7:0] _GEN_3711 = opcode_1 == 4'hf ? _GEN_1661 : _GEN_3197; // @[executor.scala 466:52]
  wire [7:0] _GEN_3712 = opcode_1 == 4'hf ? _GEN_1662 : _GEN_3198; // @[executor.scala 466:52]
  wire [7:0] _GEN_3713 = opcode_1 == 4'hf ? _GEN_1663 : _GEN_3199; // @[executor.scala 466:52]
  wire [7:0] _GEN_3714 = opcode_1 == 4'hf ? _GEN_1664 : _GEN_3200; // @[executor.scala 466:52]
  wire [7:0] _GEN_3715 = opcode_1 == 4'hf ? _GEN_1665 : _GEN_3201; // @[executor.scala 466:52]
  wire [7:0] _GEN_3716 = opcode_1 == 4'hf ? _GEN_1666 : _GEN_3202; // @[executor.scala 466:52]
  wire [7:0] _GEN_3717 = opcode_1 == 4'hf ? _GEN_1667 : _GEN_3203; // @[executor.scala 466:52]
  wire [7:0] _GEN_3718 = opcode_1 == 4'hf ? _GEN_1668 : _GEN_3204; // @[executor.scala 466:52]
  wire [7:0] _GEN_3719 = opcode_1 == 4'hf ? _GEN_1669 : _GEN_3205; // @[executor.scala 466:52]
  wire [7:0] _GEN_3720 = opcode_1 == 4'hf ? _GEN_1670 : _GEN_3206; // @[executor.scala 466:52]
  wire [7:0] _GEN_3721 = opcode_1 == 4'hf ? _GEN_1671 : _GEN_3207; // @[executor.scala 466:52]
  wire [7:0] _GEN_3722 = opcode_1 == 4'hf ? _GEN_1672 : _GEN_3208; // @[executor.scala 466:52]
  wire [7:0] _GEN_3723 = opcode_1 == 4'hf ? _GEN_1673 : _GEN_3209; // @[executor.scala 466:52]
  wire [7:0] _GEN_3724 = opcode_1 == 4'hf ? _GEN_1674 : _GEN_3210; // @[executor.scala 466:52]
  wire [7:0] _GEN_3725 = opcode_1 == 4'hf ? _GEN_1675 : _GEN_3211; // @[executor.scala 466:52]
  wire [7:0] _GEN_3726 = opcode_1 == 4'hf ? _GEN_1676 : _GEN_3212; // @[executor.scala 466:52]
  wire [7:0] _GEN_3727 = opcode_1 == 4'hf ? _GEN_1677 : _GEN_3213; // @[executor.scala 466:52]
  wire [7:0] _GEN_3728 = opcode_1 == 4'hf ? _GEN_1678 : _GEN_3214; // @[executor.scala 466:52]
  wire [7:0] _GEN_3729 = opcode_1 == 4'hf ? _GEN_1679 : _GEN_3215; // @[executor.scala 466:52]
  wire [7:0] _GEN_3730 = opcode_1 == 4'hf ? _GEN_1680 : _GEN_3216; // @[executor.scala 466:52]
  wire [7:0] _GEN_3731 = opcode_1 == 4'hf ? _GEN_1681 : _GEN_3217; // @[executor.scala 466:52]
  wire [7:0] _GEN_3732 = opcode_1 == 4'hf ? _GEN_1682 : _GEN_3218; // @[executor.scala 466:52]
  wire [7:0] _GEN_3733 = opcode_1 == 4'hf ? _GEN_1683 : _GEN_3219; // @[executor.scala 466:52]
  wire [7:0] _GEN_3734 = opcode_1 == 4'hf ? _GEN_1684 : _GEN_3220; // @[executor.scala 466:52]
  wire [7:0] _GEN_3735 = opcode_1 == 4'hf ? _GEN_1685 : _GEN_3221; // @[executor.scala 466:52]
  wire [7:0] _GEN_3736 = opcode_1 == 4'hf ? _GEN_1686 : _GEN_3222; // @[executor.scala 466:52]
  wire [7:0] _GEN_3737 = opcode_1 == 4'hf ? _GEN_1687 : _GEN_3223; // @[executor.scala 466:52]
  wire [7:0] _GEN_3738 = opcode_1 == 4'hf ? _GEN_1688 : _GEN_3224; // @[executor.scala 466:52]
  wire [7:0] _GEN_3739 = opcode_1 == 4'hf ? _GEN_1689 : _GEN_3225; // @[executor.scala 466:52]
  wire [7:0] _GEN_3740 = opcode_1 == 4'hf ? _GEN_1690 : _GEN_3226; // @[executor.scala 466:52]
  wire [7:0] _GEN_3741 = opcode_1 == 4'hf ? _GEN_1691 : _GEN_3227; // @[executor.scala 466:52]
  wire [7:0] _GEN_3742 = opcode_1 == 4'hf ? _GEN_1692 : _GEN_3228; // @[executor.scala 466:52]
  wire [7:0] _GEN_3743 = opcode_1 == 4'hf ? _GEN_1693 : _GEN_3229; // @[executor.scala 466:52]
  wire [7:0] _GEN_3744 = opcode_1 == 4'hf ? _GEN_1694 : _GEN_3230; // @[executor.scala 466:52]
  wire [7:0] _GEN_3745 = opcode_1 == 4'hf ? _GEN_1695 : _GEN_3231; // @[executor.scala 466:52]
  wire [7:0] _GEN_3746 = opcode_1 == 4'hf ? _GEN_1696 : _GEN_3232; // @[executor.scala 466:52]
  wire [7:0] _GEN_3747 = opcode_1 == 4'hf ? _GEN_1697 : _GEN_3233; // @[executor.scala 466:52]
  wire [7:0] _GEN_3748 = opcode_1 == 4'hf ? _GEN_1698 : _GEN_3234; // @[executor.scala 466:52]
  wire [7:0] _GEN_3749 = opcode_1 == 4'hf ? _GEN_1699 : _GEN_3235; // @[executor.scala 466:52]
  wire [7:0] _GEN_3750 = opcode_1 == 4'hf ? _GEN_1700 : _GEN_3236; // @[executor.scala 466:52]
  wire [7:0] _GEN_3751 = opcode_1 == 4'hf ? _GEN_1701 : _GEN_3237; // @[executor.scala 466:52]
  wire [7:0] _GEN_3752 = opcode_1 == 4'hf ? _GEN_1702 : _GEN_3238; // @[executor.scala 466:52]
  wire [7:0] _GEN_3753 = opcode_1 == 4'hf ? _GEN_1703 : _GEN_3239; // @[executor.scala 466:52]
  wire [7:0] _GEN_3754 = opcode_1 == 4'hf ? _GEN_1704 : _GEN_3240; // @[executor.scala 466:52]
  wire [7:0] _GEN_3755 = opcode_1 == 4'hf ? _GEN_1705 : _GEN_3241; // @[executor.scala 466:52]
  wire [7:0] _GEN_3756 = opcode_1 == 4'hf ? _GEN_1706 : _GEN_3242; // @[executor.scala 466:52]
  wire [7:0] _GEN_3757 = opcode_1 == 4'hf ? _GEN_1707 : _GEN_3243; // @[executor.scala 466:52]
  wire [7:0] _GEN_3758 = opcode_1 == 4'hf ? _GEN_1708 : _GEN_3244; // @[executor.scala 466:52]
  wire [7:0] _GEN_3759 = opcode_1 == 4'hf ? _GEN_1709 : _GEN_3245; // @[executor.scala 466:52]
  wire [7:0] _GEN_3760 = opcode_1 == 4'hf ? _GEN_1710 : _GEN_3246; // @[executor.scala 466:52]
  wire [7:0] _GEN_3761 = opcode_1 == 4'hf ? _GEN_1711 : _GEN_3247; // @[executor.scala 466:52]
  wire [7:0] _GEN_3762 = opcode_1 == 4'hf ? _GEN_1712 : _GEN_3248; // @[executor.scala 466:52]
  wire [7:0] _GEN_3763 = opcode_1 == 4'hf ? _GEN_1713 : _GEN_3249; // @[executor.scala 466:52]
  wire [7:0] _GEN_3764 = opcode_1 == 4'hf ? _GEN_1714 : _GEN_3250; // @[executor.scala 466:52]
  wire [7:0] _GEN_3765 = opcode_1 == 4'hf ? _GEN_1715 : _GEN_3251; // @[executor.scala 466:52]
  wire [7:0] _GEN_3766 = opcode_1 == 4'hf ? _GEN_1716 : _GEN_3252; // @[executor.scala 466:52]
  wire [7:0] _GEN_3767 = opcode_1 == 4'hf ? _GEN_1717 : _GEN_3253; // @[executor.scala 466:52]
  wire [7:0] _GEN_3768 = opcode_1 == 4'hf ? _GEN_1718 : _GEN_3254; // @[executor.scala 466:52]
  wire [7:0] _GEN_3769 = opcode_1 == 4'hf ? _GEN_1719 : _GEN_3255; // @[executor.scala 466:52]
  wire [7:0] _GEN_3770 = opcode_1 == 4'hf ? _GEN_1720 : _GEN_3256; // @[executor.scala 466:52]
  wire [7:0] _GEN_3771 = opcode_1 == 4'hf ? _GEN_1721 : _GEN_3257; // @[executor.scala 466:52]
  wire [7:0] _GEN_3772 = opcode_1 == 4'hf ? _GEN_1722 : _GEN_3258; // @[executor.scala 466:52]
  wire [7:0] _GEN_3773 = opcode_1 == 4'hf ? _GEN_1723 : _GEN_3259; // @[executor.scala 466:52]
  wire [7:0] _GEN_3774 = opcode_1 == 4'hf ? _GEN_1724 : _GEN_3260; // @[executor.scala 466:52]
  wire [7:0] _GEN_3775 = opcode_1 == 4'hf ? _GEN_1725 : _GEN_3261; // @[executor.scala 466:52]
  wire [7:0] _GEN_3776 = opcode_1 == 4'hf ? _GEN_1726 : _GEN_3262; // @[executor.scala 466:52]
  wire [7:0] _GEN_3777 = opcode_1 == 4'hf ? _GEN_1727 : _GEN_3263; // @[executor.scala 466:52]
  wire [7:0] _GEN_3778 = opcode_1 == 4'hf ? _GEN_1728 : _GEN_3264; // @[executor.scala 466:52]
  wire [7:0] _GEN_3779 = opcode_1 == 4'hf ? _GEN_1729 : _GEN_3265; // @[executor.scala 466:52]
  wire [7:0] _GEN_3780 = opcode_1 == 4'hf ? _GEN_1730 : _GEN_3266; // @[executor.scala 466:52]
  wire [7:0] _GEN_3781 = opcode_1 == 4'hf ? _GEN_1731 : _GEN_3267; // @[executor.scala 466:52]
  wire [7:0] _GEN_3782 = opcode_1 == 4'hf ? _GEN_1732 : _GEN_3268; // @[executor.scala 466:52]
  wire [7:0] _GEN_3783 = opcode_1 == 4'hf ? _GEN_1733 : _GEN_3269; // @[executor.scala 466:52]
  wire [7:0] _GEN_3784 = opcode_1 == 4'hf ? _GEN_1734 : _GEN_3270; // @[executor.scala 466:52]
  wire [7:0] _GEN_3785 = opcode_1 == 4'hf ? _GEN_1735 : _GEN_3271; // @[executor.scala 466:52]
  wire [7:0] _GEN_3786 = opcode_1 == 4'hf ? _GEN_1736 : _GEN_3272; // @[executor.scala 466:52]
  wire [7:0] _GEN_3787 = opcode_1 == 4'hf ? _GEN_1737 : _GEN_3273; // @[executor.scala 466:52]
  wire [7:0] _GEN_3788 = opcode_1 == 4'hf ? _GEN_1738 : _GEN_3274; // @[executor.scala 466:52]
  wire [7:0] _GEN_3789 = opcode_1 == 4'hf ? _GEN_1739 : _GEN_3275; // @[executor.scala 466:52]
  wire [7:0] _GEN_3790 = opcode_1 == 4'hf ? _GEN_1740 : _GEN_3276; // @[executor.scala 466:52]
  wire [7:0] _GEN_3791 = opcode_1 == 4'hf ? _GEN_1741 : _GEN_3277; // @[executor.scala 466:52]
  wire [7:0] _GEN_3792 = opcode_1 == 4'hf ? _GEN_1742 : _GEN_3278; // @[executor.scala 466:52]
  wire [7:0] _GEN_3793 = opcode_1 == 4'hf ? _GEN_1743 : _GEN_3279; // @[executor.scala 466:52]
  wire [7:0] _GEN_3794 = opcode_1 == 4'hf ? _GEN_1744 : _GEN_3280; // @[executor.scala 466:52]
  wire [7:0] _GEN_3795 = opcode_1 == 4'hf ? _GEN_1745 : _GEN_3281; // @[executor.scala 466:52]
  wire [7:0] _GEN_3796 = opcode_1 == 4'hf ? _GEN_1746 : _GEN_3282; // @[executor.scala 466:52]
  wire [7:0] _GEN_3797 = opcode_1 == 4'hf ? _GEN_1747 : _GEN_3283; // @[executor.scala 466:52]
  wire [7:0] _GEN_3798 = opcode_1 == 4'hf ? _GEN_1748 : _GEN_3284; // @[executor.scala 466:52]
  wire [7:0] _GEN_3799 = opcode_1 == 4'hf ? _GEN_1749 : _GEN_3285; // @[executor.scala 466:52]
  wire [7:0] _GEN_3800 = opcode_1 == 4'hf ? _GEN_1750 : _GEN_3286; // @[executor.scala 466:52]
  wire [7:0] _GEN_3801 = opcode_1 == 4'hf ? _GEN_1751 : _GEN_3287; // @[executor.scala 466:52]
  wire [7:0] _GEN_3802 = opcode_1 == 4'hf ? _GEN_1752 : _GEN_3288; // @[executor.scala 466:52]
  wire [7:0] _GEN_3803 = opcode_1 == 4'hf ? _GEN_1753 : _GEN_3289; // @[executor.scala 466:52]
  wire [7:0] _GEN_3804 = opcode_1 == 4'hf ? _GEN_1754 : _GEN_3290; // @[executor.scala 466:52]
  wire [7:0] _GEN_3805 = opcode_1 == 4'hf ? _GEN_1755 : _GEN_3291; // @[executor.scala 466:52]
  wire [7:0] _GEN_3806 = opcode_1 == 4'hf ? _GEN_1756 : _GEN_3292; // @[executor.scala 466:52]
  wire [7:0] _GEN_3807 = opcode_1 == 4'hf ? _GEN_1757 : _GEN_3293; // @[executor.scala 466:52]
  wire [7:0] _GEN_3808 = opcode_1 == 4'hf ? _GEN_1758 : _GEN_3294; // @[executor.scala 466:52]
  wire [7:0] _GEN_3809 = opcode_1 == 4'hf ? _GEN_1759 : _GEN_3295; // @[executor.scala 466:52]
  wire [7:0] _GEN_3810 = opcode_1 == 4'hf ? _GEN_1760 : _GEN_3296; // @[executor.scala 466:52]
  wire [7:0] _GEN_3811 = opcode_1 == 4'hf ? _GEN_1761 : _GEN_3297; // @[executor.scala 466:52]
  wire [7:0] _GEN_3812 = opcode_1 == 4'hf ? _GEN_1762 : _GEN_3298; // @[executor.scala 466:52]
  wire [7:0] _GEN_3813 = opcode_1 == 4'hf ? _GEN_1763 : _GEN_3299; // @[executor.scala 466:52]
  wire [7:0] _GEN_3814 = opcode_1 == 4'hf ? _GEN_1764 : _GEN_3300; // @[executor.scala 466:52]
  wire [7:0] _GEN_3815 = opcode_1 == 4'hf ? _GEN_1765 : _GEN_3301; // @[executor.scala 466:52]
  wire [7:0] _GEN_3816 = opcode_1 == 4'hf ? _GEN_1766 : _GEN_3302; // @[executor.scala 466:52]
  wire [7:0] _GEN_3817 = opcode_1 == 4'hf ? _GEN_1767 : _GEN_3303; // @[executor.scala 466:52]
  wire [7:0] _GEN_3818 = opcode_1 == 4'hf ? _GEN_1768 : _GEN_3304; // @[executor.scala 466:52]
  wire [7:0] _GEN_3819 = opcode_1 == 4'hf ? _GEN_1769 : _GEN_3305; // @[executor.scala 466:52]
  wire [7:0] _GEN_3820 = opcode_1 == 4'hf ? _GEN_1770 : _GEN_3306; // @[executor.scala 466:52]
  wire [7:0] _GEN_3821 = opcode_1 == 4'hf ? _GEN_1771 : _GEN_3307; // @[executor.scala 466:52]
  wire [7:0] _GEN_3822 = opcode_1 == 4'hf ? _GEN_1772 : _GEN_3308; // @[executor.scala 466:52]
  wire [7:0] _GEN_3823 = opcode_1 == 4'hf ? _GEN_1773 : _GEN_3309; // @[executor.scala 466:52]
  wire [7:0] _GEN_3824 = opcode_1 == 4'hf ? _GEN_1774 : _GEN_3310; // @[executor.scala 466:52]
  wire [7:0] _GEN_3825 = opcode_1 == 4'hf ? _GEN_1775 : _GEN_3311; // @[executor.scala 466:52]
  wire [7:0] _GEN_3826 = opcode_1 == 4'hf ? _GEN_1776 : _GEN_3312; // @[executor.scala 466:52]
  wire [7:0] _GEN_3827 = opcode_1 == 4'hf ? _GEN_1777 : _GEN_3313; // @[executor.scala 466:52]
  wire [7:0] _GEN_3828 = opcode_1 == 4'hf ? _GEN_1778 : _GEN_3314; // @[executor.scala 466:52]
  wire [7:0] _GEN_3829 = opcode_1 == 4'hf ? _GEN_1779 : _GEN_3315; // @[executor.scala 466:52]
  wire [7:0] _GEN_3830 = opcode_1 == 4'hf ? _GEN_1780 : _GEN_3316; // @[executor.scala 466:52]
  wire [7:0] _GEN_3831 = opcode_1 == 4'hf ? _GEN_1781 : _GEN_3317; // @[executor.scala 466:52]
  wire [7:0] _GEN_3832 = opcode_1 == 4'hf ? _GEN_1782 : _GEN_3318; // @[executor.scala 466:52]
  wire [7:0] _GEN_3833 = opcode_1 == 4'hf ? _GEN_1783 : _GEN_3319; // @[executor.scala 466:52]
  wire [7:0] _GEN_3834 = opcode_1 == 4'hf ? _GEN_1784 : _GEN_3320; // @[executor.scala 466:52]
  wire [7:0] _GEN_3835 = opcode_1 == 4'hf ? _GEN_1785 : _GEN_3321; // @[executor.scala 466:52]
  wire [7:0] _GEN_3836 = opcode_1 == 4'hf ? _GEN_1786 : _GEN_3322; // @[executor.scala 466:52]
  wire [7:0] _GEN_3837 = opcode_1 == 4'hf ? _GEN_1787 : _GEN_3323; // @[executor.scala 466:52]
  wire [7:0] _GEN_3838 = opcode_1 == 4'hf ? _GEN_1788 : _GEN_3324; // @[executor.scala 466:52]
  wire [7:0] _GEN_3839 = opcode_1 == 4'hf ? _GEN_1789 : _GEN_3325; // @[executor.scala 466:52]
  wire [7:0] _GEN_3840 = opcode_1 == 4'hf ? _GEN_1790 : _GEN_3326; // @[executor.scala 466:52]
  wire [7:0] _GEN_3841 = opcode_1 == 4'hf ? _GEN_1791 : _GEN_3327; // @[executor.scala 466:52]
  wire [7:0] _GEN_3842 = opcode_1 == 4'hf ? _GEN_1792 : _GEN_3328; // @[executor.scala 466:52]
  wire [7:0] _GEN_3843 = opcode_1 == 4'hf ? _GEN_1793 : _GEN_3329; // @[executor.scala 466:52]
  wire [7:0] _GEN_3844 = opcode_1 == 4'hf ? _GEN_1794 : _GEN_3330; // @[executor.scala 466:52]
  wire [7:0] _GEN_3845 = opcode_1 == 4'hf ? _GEN_1795 : _GEN_3331; // @[executor.scala 466:52]
  wire [7:0] _GEN_3846 = opcode_1 == 4'hf ? _GEN_1796 : _GEN_3332; // @[executor.scala 466:52]
  wire [7:0] _GEN_3847 = opcode_1 == 4'hf ? _GEN_1797 : _GEN_3333; // @[executor.scala 466:52]
  wire [7:0] _GEN_3848 = opcode_1 == 4'hf ? _GEN_1798 : _GEN_3334; // @[executor.scala 466:52]
  wire [7:0] _GEN_3849 = opcode_1 == 4'hf ? _GEN_1799 : _GEN_3335; // @[executor.scala 466:52]
  wire [7:0] _GEN_3850 = opcode_1 == 4'hf ? _GEN_1800 : _GEN_3336; // @[executor.scala 466:52]
  wire [7:0] _GEN_3851 = opcode_1 == 4'hf ? _GEN_1801 : _GEN_3337; // @[executor.scala 466:52]
  wire [7:0] _GEN_3852 = opcode_1 == 4'hf ? _GEN_1802 : _GEN_3338; // @[executor.scala 466:52]
  wire [7:0] _GEN_3853 = opcode_1 == 4'hf ? _GEN_1803 : _GEN_3339; // @[executor.scala 466:52]
  wire [7:0] _GEN_3854 = opcode_1 == 4'hf ? _GEN_1804 : _GEN_3340; // @[executor.scala 466:52]
  wire [7:0] _GEN_3855 = opcode_1 == 4'hf ? _GEN_1805 : _GEN_3341; // @[executor.scala 466:52]
  wire [7:0] _GEN_3856 = opcode_1 == 4'hf ? _GEN_1806 : _GEN_3342; // @[executor.scala 466:52]
  wire [7:0] _GEN_3857 = opcode_1 == 4'hf ? _GEN_1807 : _GEN_3343; // @[executor.scala 466:52]
  wire [7:0] _GEN_3858 = opcode_1 == 4'hf ? _GEN_1808 : _GEN_3344; // @[executor.scala 466:52]
  wire [7:0] _GEN_3859 = opcode_1 == 4'hf ? _GEN_1809 : _GEN_3345; // @[executor.scala 466:52]
  wire [7:0] _GEN_3860 = opcode_1 == 4'hf ? _GEN_1810 : _GEN_3346; // @[executor.scala 466:52]
  wire [7:0] _GEN_3861 = opcode_1 == 4'hf ? _GEN_1811 : _GEN_3347; // @[executor.scala 466:52]
  wire [7:0] _GEN_3862 = opcode_1 == 4'hf ? _GEN_1812 : _GEN_3348; // @[executor.scala 466:52]
  wire [7:0] _GEN_3863 = opcode_1 == 4'hf ? _GEN_1813 : _GEN_3349; // @[executor.scala 466:52]
  wire [7:0] _GEN_3864 = opcode_1 == 4'hf ? _GEN_1814 : _GEN_3350; // @[executor.scala 466:52]
  wire [7:0] _GEN_3865 = opcode_1 == 4'hf ? _GEN_1815 : _GEN_3351; // @[executor.scala 466:52]
  wire [7:0] _GEN_3866 = opcode_1 == 4'hf ? _GEN_1816 : _GEN_3352; // @[executor.scala 466:52]
  wire [7:0] _GEN_3867 = opcode_1 == 4'hf ? _GEN_1817 : _GEN_3353; // @[executor.scala 466:52]
  wire [7:0] _GEN_3868 = opcode_1 == 4'hf ? _GEN_1818 : _GEN_3354; // @[executor.scala 466:52]
  wire [7:0] _GEN_3869 = opcode_1 == 4'hf ? _GEN_1819 : _GEN_3355; // @[executor.scala 466:52]
  wire [7:0] _GEN_3870 = opcode_1 == 4'hf ? _GEN_1820 : _GEN_3356; // @[executor.scala 466:52]
  wire [7:0] _GEN_3871 = opcode_1 == 4'hf ? _GEN_1821 : _GEN_3357; // @[executor.scala 466:52]
  wire [7:0] _GEN_3872 = opcode_1 == 4'hf ? _GEN_1822 : _GEN_3358; // @[executor.scala 466:52]
  wire [7:0] _GEN_3873 = opcode_1 == 4'hf ? _GEN_1823 : _GEN_3359; // @[executor.scala 466:52]
  wire [7:0] _GEN_3874 = opcode_1 == 4'hf ? _GEN_1824 : _GEN_3360; // @[executor.scala 466:52]
  wire [7:0] _GEN_3875 = opcode_1 == 4'hf ? _GEN_1825 : _GEN_3361; // @[executor.scala 466:52]
  wire [7:0] _GEN_3876 = opcode_1 == 4'hf ? _GEN_1826 : _GEN_3362; // @[executor.scala 466:52]
  wire [7:0] _GEN_3877 = opcode_1 == 4'hf ? _GEN_1827 : _GEN_3363; // @[executor.scala 466:52]
  wire [7:0] _GEN_3878 = opcode_1 == 4'hf ? _GEN_1828 : _GEN_3364; // @[executor.scala 466:52]
  wire [7:0] _GEN_3879 = opcode_1 == 4'hf ? _GEN_1829 : _GEN_3365; // @[executor.scala 466:52]
  wire [7:0] _GEN_3880 = opcode_1 == 4'hf ? _GEN_1830 : _GEN_3366; // @[executor.scala 466:52]
  wire [7:0] _GEN_3881 = opcode_1 == 4'hf ? _GEN_1831 : _GEN_3367; // @[executor.scala 466:52]
  wire [7:0] _GEN_3882 = opcode_1 == 4'hf ? _GEN_1832 : _GEN_3368; // @[executor.scala 466:52]
  wire [7:0] _GEN_3883 = opcode_1 == 4'hf ? _GEN_1833 : _GEN_3369; // @[executor.scala 466:52]
  wire [7:0] _GEN_3884 = opcode_1 == 4'hf ? _GEN_1834 : _GEN_3370; // @[executor.scala 466:52]
  wire [7:0] _GEN_3885 = opcode_1 == 4'hf ? _GEN_1835 : _GEN_3371; // @[executor.scala 466:52]
  wire [7:0] _GEN_3886 = opcode_1 == 4'hf ? _GEN_1836 : _GEN_3372; // @[executor.scala 466:52]
  wire [7:0] _GEN_3887 = opcode_1 == 4'hf ? _GEN_1837 : _GEN_3373; // @[executor.scala 466:52]
  wire [7:0] _GEN_3888 = opcode_1 == 4'hf ? _GEN_1838 : _GEN_3374; // @[executor.scala 466:52]
  wire [7:0] _GEN_3889 = opcode_1 == 4'hf ? _GEN_1839 : _GEN_3375; // @[executor.scala 466:52]
  wire [7:0] _GEN_3890 = opcode_1 == 4'hf ? _GEN_1840 : _GEN_3376; // @[executor.scala 466:52]
  wire [7:0] _GEN_3891 = opcode_1 == 4'hf ? _GEN_1841 : _GEN_3377; // @[executor.scala 466:52]
  wire [7:0] _GEN_3892 = opcode_1 == 4'hf ? _GEN_1842 : _GEN_3378; // @[executor.scala 466:52]
  wire [7:0] _GEN_3893 = opcode_1 == 4'hf ? _GEN_1843 : _GEN_3379; // @[executor.scala 466:52]
  wire [7:0] _GEN_3894 = opcode_1 == 4'hf ? _GEN_1844 : _GEN_3380; // @[executor.scala 466:52]
  wire [7:0] _GEN_3895 = opcode_1 == 4'hf ? _GEN_1845 : _GEN_3381; // @[executor.scala 466:52]
  wire [7:0] _GEN_3896 = opcode_1 == 4'hf ? _GEN_1846 : _GEN_3382; // @[executor.scala 466:52]
  wire [7:0] _GEN_3897 = opcode_1 == 4'hf ? _GEN_1847 : _GEN_3383; // @[executor.scala 466:52]
  wire [7:0] _GEN_3898 = opcode_1 == 4'hf ? _GEN_1848 : _GEN_3384; // @[executor.scala 466:52]
  wire [7:0] _GEN_3899 = opcode_1 == 4'hf ? _GEN_1849 : _GEN_3385; // @[executor.scala 466:52]
  wire [7:0] _GEN_3900 = opcode_1 == 4'hf ? _GEN_1850 : _GEN_3386; // @[executor.scala 466:52]
  wire [7:0] _GEN_3901 = opcode_1 == 4'hf ? _GEN_1851 : _GEN_3387; // @[executor.scala 466:52]
  wire [7:0] _GEN_3902 = opcode_1 == 4'hf ? _GEN_1852 : _GEN_3388; // @[executor.scala 466:52]
  wire [7:0] _GEN_3903 = opcode_1 == 4'hf ? _GEN_1853 : _GEN_3389; // @[executor.scala 466:52]
  wire [7:0] _GEN_3904 = opcode_1 == 4'hf ? _GEN_1854 : _GEN_3390; // @[executor.scala 466:52]
  wire [7:0] _GEN_3905 = opcode_1 == 4'hf ? _GEN_1855 : _GEN_3391; // @[executor.scala 466:52]
  wire [7:0] _GEN_3906 = opcode_1 == 4'hf ? _GEN_1856 : _GEN_3392; // @[executor.scala 466:52]
  wire [7:0] _GEN_3907 = opcode_1 == 4'hf ? _GEN_1857 : _GEN_3393; // @[executor.scala 466:52]
  wire [7:0] _GEN_3908 = opcode_1 == 4'hf ? _GEN_1858 : _GEN_3394; // @[executor.scala 466:52]
  wire [7:0] _GEN_3909 = opcode_1 == 4'hf ? _GEN_1859 : _GEN_3395; // @[executor.scala 466:52]
  wire [7:0] _GEN_3910 = opcode_1 == 4'hf ? _GEN_1860 : _GEN_3396; // @[executor.scala 466:52]
  wire [7:0] _GEN_3911 = opcode_1 == 4'hf ? _GEN_1861 : _GEN_3397; // @[executor.scala 466:52]
  wire [7:0] _GEN_3912 = opcode_1 == 4'hf ? _GEN_1862 : _GEN_3398; // @[executor.scala 466:52]
  wire [7:0] _GEN_3913 = opcode_1 == 4'hf ? _GEN_1863 : _GEN_3399; // @[executor.scala 466:52]
  wire [7:0] _GEN_3914 = opcode_1 == 4'hf ? _GEN_1864 : _GEN_3400; // @[executor.scala 466:52]
  wire [7:0] _GEN_3915 = opcode_1 == 4'hf ? _GEN_1865 : _GEN_3401; // @[executor.scala 466:52]
  wire [7:0] _GEN_3916 = opcode_1 == 4'hf ? _GEN_1866 : _GEN_3402; // @[executor.scala 466:52]
  wire [7:0] _GEN_3917 = opcode_1 == 4'hf ? _GEN_1867 : _GEN_3403; // @[executor.scala 466:52]
  wire [7:0] _GEN_3918 = opcode_1 == 4'hf ? _GEN_1868 : _GEN_3404; // @[executor.scala 466:52]
  wire [7:0] _GEN_3919 = opcode_1 == 4'hf ? _GEN_1869 : _GEN_3405; // @[executor.scala 466:52]
  wire [7:0] _GEN_3920 = opcode_1 == 4'hf ? _GEN_1870 : _GEN_3406; // @[executor.scala 466:52]
  wire [7:0] _GEN_3921 = opcode_1 == 4'hf ? _GEN_1871 : _GEN_3407; // @[executor.scala 466:52]
  wire [7:0] _GEN_3922 = opcode_1 == 4'hf ? _GEN_1872 : _GEN_3408; // @[executor.scala 466:52]
  wire [7:0] _GEN_3923 = opcode_1 == 4'hf ? _GEN_1873 : _GEN_3409; // @[executor.scala 466:52]
  wire [7:0] _GEN_3924 = opcode_1 == 4'hf ? _GEN_1874 : _GEN_3410; // @[executor.scala 466:52]
  wire [7:0] _GEN_3925 = opcode_1 == 4'hf ? _GEN_1875 : _GEN_3411; // @[executor.scala 466:52]
  wire [7:0] _GEN_3926 = opcode_1 == 4'hf ? _GEN_1876 : _GEN_3412; // @[executor.scala 466:52]
  wire [7:0] _GEN_3927 = opcode_1 == 4'hf ? _GEN_1877 : _GEN_3413; // @[executor.scala 466:52]
  wire [7:0] _GEN_3928 = opcode_1 == 4'hf ? _GEN_1878 : _GEN_3414; // @[executor.scala 466:52]
  wire [7:0] _GEN_3929 = opcode_1 == 4'hf ? _GEN_1879 : _GEN_3415; // @[executor.scala 466:52]
  wire [7:0] _GEN_3930 = opcode_1 == 4'hf ? _GEN_1880 : _GEN_3416; // @[executor.scala 466:52]
  wire [7:0] _GEN_3931 = opcode_1 == 4'hf ? _GEN_1881 : _GEN_3417; // @[executor.scala 466:52]
  wire [7:0] _GEN_3932 = opcode_1 == 4'hf ? _GEN_1882 : _GEN_3418; // @[executor.scala 466:52]
  wire [7:0] _GEN_3933 = opcode_1 == 4'hf ? _GEN_1883 : _GEN_3419; // @[executor.scala 466:52]
  wire [7:0] _GEN_3934 = opcode_1 == 4'hf ? _GEN_1884 : _GEN_3420; // @[executor.scala 466:52]
  wire [7:0] _GEN_3935 = opcode_1 == 4'hf ? _GEN_1885 : _GEN_3421; // @[executor.scala 466:52]
  wire [7:0] _GEN_3936 = opcode_1 == 4'hf ? _GEN_1886 : _GEN_3422; // @[executor.scala 466:52]
  wire [7:0] _GEN_3937 = opcode_1 == 4'hf ? _GEN_1887 : _GEN_3423; // @[executor.scala 466:52]
  wire [7:0] _GEN_3938 = opcode_1 == 4'hf ? _GEN_1888 : _GEN_3424; // @[executor.scala 466:52]
  wire [7:0] _GEN_3939 = opcode_1 == 4'hf ? _GEN_1889 : _GEN_3425; // @[executor.scala 466:52]
  wire [7:0] _GEN_3940 = opcode_1 == 4'hf ? _GEN_1890 : _GEN_3426; // @[executor.scala 466:52]
  wire [7:0] _GEN_3941 = opcode_1 == 4'hf ? _GEN_1891 : _GEN_3427; // @[executor.scala 466:52]
  wire [7:0] _GEN_3942 = opcode_1 == 4'hf ? _GEN_1892 : _GEN_3428; // @[executor.scala 466:52]
  wire [7:0] _GEN_3943 = opcode_1 == 4'hf ? _GEN_1893 : _GEN_3429; // @[executor.scala 466:52]
  wire [7:0] _GEN_3944 = opcode_1 == 4'hf ? _GEN_1894 : _GEN_3430; // @[executor.scala 466:52]
  wire [7:0] _GEN_3945 = opcode_1 == 4'hf ? _GEN_1895 : _GEN_3431; // @[executor.scala 466:52]
  wire [7:0] _GEN_3946 = opcode_1 == 4'hf ? _GEN_1896 : _GEN_3432; // @[executor.scala 466:52]
  wire [7:0] _GEN_3947 = opcode_1 == 4'hf ? _GEN_1897 : _GEN_3433; // @[executor.scala 466:52]
  wire [7:0] _GEN_3948 = opcode_1 == 4'hf ? _GEN_1898 : _GEN_3434; // @[executor.scala 466:52]
  wire [7:0] _GEN_3949 = opcode_1 == 4'hf ? _GEN_1899 : _GEN_3435; // @[executor.scala 466:52]
  wire [7:0] _GEN_3950 = opcode_1 == 4'hf ? _GEN_1900 : _GEN_3436; // @[executor.scala 466:52]
  wire [7:0] _GEN_3951 = opcode_1 == 4'hf ? _GEN_1901 : _GEN_3437; // @[executor.scala 466:52]
  wire [7:0] _GEN_3952 = opcode_1 == 4'hf ? _GEN_1902 : _GEN_3438; // @[executor.scala 466:52]
  wire [7:0] _GEN_3953 = opcode_1 == 4'hf ? _GEN_1903 : _GEN_3439; // @[executor.scala 466:52]
  wire [7:0] _GEN_3954 = opcode_1 == 4'hf ? _GEN_1904 : _GEN_3440; // @[executor.scala 466:52]
  wire [7:0] _GEN_3955 = opcode_1 == 4'hf ? _GEN_1905 : _GEN_3441; // @[executor.scala 466:52]
  wire [7:0] _GEN_3956 = opcode_1 == 4'hf ? _GEN_1906 : _GEN_3442; // @[executor.scala 466:52]
  wire [7:0] _GEN_3957 = opcode_1 == 4'hf ? _GEN_1907 : _GEN_3443; // @[executor.scala 466:52]
  wire [7:0] _GEN_3958 = opcode_1 == 4'hf ? _GEN_1908 : _GEN_3444; // @[executor.scala 466:52]
  wire [7:0] _GEN_3959 = opcode_1 == 4'hf ? _GEN_1909 : _GEN_3445; // @[executor.scala 466:52]
  wire [7:0] _GEN_3960 = opcode_1 == 4'hf ? _GEN_1910 : _GEN_3446; // @[executor.scala 466:52]
  wire [7:0] _GEN_3961 = opcode_1 == 4'hf ? _GEN_1911 : _GEN_3447; // @[executor.scala 466:52]
  wire [7:0] _GEN_3962 = opcode_1 == 4'hf ? _GEN_1912 : _GEN_3448; // @[executor.scala 466:52]
  wire [7:0] _GEN_3963 = opcode_1 == 4'hf ? _GEN_1913 : _GEN_3449; // @[executor.scala 466:52]
  wire [7:0] _GEN_3964 = opcode_1 == 4'hf ? _GEN_1914 : _GEN_3450; // @[executor.scala 466:52]
  wire [7:0] _GEN_3965 = opcode_1 == 4'hf ? _GEN_1915 : _GEN_3451; // @[executor.scala 466:52]
  wire [7:0] _GEN_3966 = opcode_1 == 4'hf ? _GEN_1916 : _GEN_3452; // @[executor.scala 466:52]
  wire [7:0] _GEN_3967 = opcode_1 == 4'hf ? _GEN_1917 : _GEN_3453; // @[executor.scala 466:52]
  wire [7:0] _GEN_3968 = opcode_1 == 4'hf ? _GEN_1918 : _GEN_3454; // @[executor.scala 466:52]
  wire [7:0] _GEN_3969 = opcode_1 == 4'hf ? _GEN_1919 : _GEN_3455; // @[executor.scala 466:52]
  wire [7:0] _GEN_3970 = opcode_1 == 4'hf ? _GEN_1920 : _GEN_3456; // @[executor.scala 466:52]
  wire [7:0] _GEN_3971 = opcode_1 == 4'hf ? _GEN_1921 : _GEN_3457; // @[executor.scala 466:52]
  wire [7:0] _GEN_3972 = opcode_1 == 4'hf ? _GEN_1922 : _GEN_3458; // @[executor.scala 466:52]
  wire [7:0] _GEN_3973 = opcode_1 == 4'hf ? _GEN_1923 : _GEN_3459; // @[executor.scala 466:52]
  wire [7:0] _GEN_3974 = opcode_1 == 4'hf ? _GEN_1924 : _GEN_3460; // @[executor.scala 466:52]
  wire [7:0] _GEN_3975 = opcode_1 == 4'hf ? _GEN_1925 : _GEN_3461; // @[executor.scala 466:52]
  wire [7:0] _GEN_3976 = opcode_1 == 4'hf ? _GEN_1926 : _GEN_3462; // @[executor.scala 466:52]
  wire [7:0] _GEN_3977 = opcode_1 == 4'hf ? _GEN_1927 : _GEN_3463; // @[executor.scala 466:52]
  wire [7:0] _GEN_3978 = opcode_1 == 4'hf ? _GEN_1928 : _GEN_3464; // @[executor.scala 466:52]
  wire [7:0] _GEN_3979 = opcode_1 == 4'hf ? _GEN_1929 : _GEN_3465; // @[executor.scala 466:52]
  wire [7:0] _GEN_3980 = opcode_1 == 4'hf ? _GEN_1930 : _GEN_3466; // @[executor.scala 466:52]
  wire [7:0] _GEN_3981 = opcode_1 == 4'hf ? _GEN_1931 : _GEN_3467; // @[executor.scala 466:52]
  wire [7:0] _GEN_3982 = opcode_1 == 4'hf ? _GEN_1932 : _GEN_3468; // @[executor.scala 466:52]
  wire [7:0] _GEN_3983 = opcode_1 == 4'hf ? _GEN_1933 : _GEN_3469; // @[executor.scala 466:52]
  wire [7:0] _GEN_3984 = opcode_1 == 4'hf ? _GEN_1934 : _GEN_3470; // @[executor.scala 466:52]
  wire [7:0] _GEN_3985 = opcode_1 == 4'hf ? _GEN_1935 : _GEN_3471; // @[executor.scala 466:52]
  wire [7:0] _GEN_3986 = opcode_1 == 4'hf ? _GEN_1936 : _GEN_3472; // @[executor.scala 466:52]
  wire [7:0] _GEN_3987 = opcode_1 == 4'hf ? _GEN_1937 : _GEN_3473; // @[executor.scala 466:52]
  wire [7:0] _GEN_3988 = opcode_1 == 4'hf ? _GEN_1938 : _GEN_3474; // @[executor.scala 466:52]
  wire [7:0] _GEN_3989 = opcode_1 == 4'hf ? _GEN_1939 : _GEN_3475; // @[executor.scala 466:52]
  wire [7:0] _GEN_3990 = opcode_1 == 4'hf ? _GEN_1940 : _GEN_3476; // @[executor.scala 466:52]
  wire [7:0] _GEN_3991 = opcode_1 == 4'hf ? _GEN_1941 : _GEN_3477; // @[executor.scala 466:52]
  wire [7:0] _GEN_3992 = opcode_1 == 4'hf ? _GEN_1942 : _GEN_3478; // @[executor.scala 466:52]
  wire [7:0] _GEN_3993 = opcode_1 == 4'hf ? _GEN_1943 : _GEN_3479; // @[executor.scala 466:52]
  wire [7:0] _GEN_3994 = opcode_1 == 4'hf ? _GEN_1944 : _GEN_3480; // @[executor.scala 466:52]
  wire [7:0] _GEN_3995 = opcode_1 == 4'hf ? _GEN_1945 : _GEN_3481; // @[executor.scala 466:52]
  wire [7:0] _GEN_3996 = opcode_1 == 4'hf ? _GEN_1946 : _GEN_3482; // @[executor.scala 466:52]
  wire [7:0] _GEN_3997 = opcode_1 == 4'hf ? _GEN_1947 : _GEN_3483; // @[executor.scala 466:52]
  wire [7:0] _GEN_3998 = opcode_1 == 4'hf ? _GEN_1948 : _GEN_3484; // @[executor.scala 466:52]
  wire [7:0] _GEN_3999 = opcode_1 == 4'hf ? _GEN_1949 : _GEN_3485; // @[executor.scala 466:52]
  wire [7:0] _GEN_4000 = opcode_1 == 4'hf ? _GEN_1950 : _GEN_3486; // @[executor.scala 466:52]
  wire [7:0] _GEN_4001 = opcode_1 == 4'hf ? _GEN_1951 : _GEN_3487; // @[executor.scala 466:52]
  wire [7:0] _GEN_4002 = opcode_1 == 4'hf ? _GEN_1952 : _GEN_3488; // @[executor.scala 466:52]
  wire [7:0] _GEN_4003 = opcode_1 == 4'hf ? _GEN_1953 : _GEN_3489; // @[executor.scala 466:52]
  wire [7:0] _GEN_4004 = opcode_1 == 4'hf ? _GEN_1954 : _GEN_3490; // @[executor.scala 466:52]
  wire [7:0] _GEN_4005 = opcode_1 == 4'hf ? _GEN_1955 : _GEN_3491; // @[executor.scala 466:52]
  wire [7:0] _GEN_4006 = opcode_1 == 4'hf ? _GEN_1956 : _GEN_3492; // @[executor.scala 466:52]
  wire [7:0] _GEN_4007 = opcode_1 == 4'hf ? _GEN_1957 : _GEN_3493; // @[executor.scala 466:52]
  wire [7:0] _GEN_4008 = opcode_1 == 4'hf ? _GEN_1958 : _GEN_3494; // @[executor.scala 466:52]
  wire [7:0] _GEN_4009 = opcode_1 == 4'hf ? _GEN_1959 : _GEN_3495; // @[executor.scala 466:52]
  wire [7:0] _GEN_4010 = opcode_1 == 4'hf ? _GEN_1960 : _GEN_3496; // @[executor.scala 466:52]
  wire [7:0] _GEN_4011 = opcode_1 == 4'hf ? _GEN_1961 : _GEN_3497; // @[executor.scala 466:52]
  wire [7:0] _GEN_4012 = opcode_1 == 4'hf ? _GEN_1962 : _GEN_3498; // @[executor.scala 466:52]
  wire [7:0] _GEN_4013 = opcode_1 == 4'hf ? _GEN_1963 : _GEN_3499; // @[executor.scala 466:52]
  wire [7:0] _GEN_4014 = opcode_1 == 4'hf ? _GEN_1964 : _GEN_3500; // @[executor.scala 466:52]
  wire [7:0] _GEN_4015 = opcode_1 == 4'hf ? _GEN_1965 : _GEN_3501; // @[executor.scala 466:52]
  wire [7:0] _GEN_4016 = opcode_1 == 4'hf ? _GEN_1966 : _GEN_3502; // @[executor.scala 466:52]
  wire [7:0] _GEN_4017 = opcode_1 == 4'hf ? _GEN_1967 : _GEN_3503; // @[executor.scala 466:52]
  wire [7:0] _GEN_4018 = opcode_1 == 4'hf ? _GEN_1968 : _GEN_3504; // @[executor.scala 466:52]
  wire [7:0] _GEN_4019 = opcode_1 == 4'hf ? _GEN_1969 : _GEN_3505; // @[executor.scala 466:52]
  wire [7:0] _GEN_4020 = opcode_1 == 4'hf ? _GEN_1970 : _GEN_3506; // @[executor.scala 466:52]
  wire [7:0] _GEN_4021 = opcode_1 == 4'hf ? _GEN_1971 : _GEN_3507; // @[executor.scala 466:52]
  wire [7:0] _GEN_4022 = opcode_1 == 4'hf ? _GEN_1972 : _GEN_3508; // @[executor.scala 466:52]
  wire [7:0] _GEN_4023 = opcode_1 == 4'hf ? _GEN_1973 : _GEN_3509; // @[executor.scala 466:52]
  wire [7:0] _GEN_4024 = opcode_1 == 4'hf ? _GEN_1974 : _GEN_3510; // @[executor.scala 466:52]
  wire [7:0] _GEN_4025 = opcode_1 == 4'hf ? _GEN_1975 : _GEN_3511; // @[executor.scala 466:52]
  wire [7:0] _GEN_4026 = opcode_1 == 4'hf ? _GEN_1976 : _GEN_3512; // @[executor.scala 466:52]
  wire [7:0] _GEN_4027 = opcode_1 == 4'hf ? _GEN_1977 : _GEN_3513; // @[executor.scala 466:52]
  wire [7:0] _GEN_4028 = opcode_1 == 4'hf ? _GEN_1978 : _GEN_3514; // @[executor.scala 466:52]
  wire [7:0] _GEN_4029 = opcode_1 == 4'hf ? _GEN_1979 : _GEN_3515; // @[executor.scala 466:52]
  wire [7:0] _GEN_4030 = opcode_1 == 4'hf ? _GEN_1980 : _GEN_3516; // @[executor.scala 466:52]
  wire [7:0] _GEN_4031 = opcode_1 == 4'hf ? _GEN_1981 : _GEN_3517; // @[executor.scala 466:52]
  wire [7:0] _GEN_4032 = opcode_1 == 4'hf ? _GEN_1982 : _GEN_3518; // @[executor.scala 466:52]
  wire [7:0] _GEN_4033 = opcode_1 == 4'hf ? _GEN_1983 : _GEN_3519; // @[executor.scala 466:52]
  wire [7:0] _GEN_4034 = opcode_1 == 4'hf ? _GEN_1984 : _GEN_3520; // @[executor.scala 466:52]
  wire [7:0] _GEN_4035 = opcode_1 == 4'hf ? _GEN_1985 : _GEN_3521; // @[executor.scala 466:52]
  wire [7:0] _GEN_4036 = opcode_1 == 4'hf ? _GEN_1986 : _GEN_3522; // @[executor.scala 466:52]
  wire [7:0] _GEN_4037 = opcode_1 == 4'hf ? _GEN_1987 : _GEN_3523; // @[executor.scala 466:52]
  wire [7:0] _GEN_4038 = opcode_1 == 4'hf ? _GEN_1988 : _GEN_3524; // @[executor.scala 466:52]
  wire [7:0] _GEN_4039 = opcode_1 == 4'hf ? _GEN_1989 : _GEN_3525; // @[executor.scala 466:52]
  wire [7:0] _GEN_4040 = opcode_1 == 4'hf ? _GEN_1990 : _GEN_3526; // @[executor.scala 466:52]
  wire [7:0] _GEN_4041 = opcode_1 == 4'hf ? _GEN_1991 : _GEN_3527; // @[executor.scala 466:52]
  wire [7:0] _GEN_4042 = opcode_1 == 4'hf ? _GEN_1992 : _GEN_3528; // @[executor.scala 466:52]
  wire [7:0] _GEN_4043 = opcode_1 == 4'hf ? _GEN_1993 : _GEN_3529; // @[executor.scala 466:52]
  wire [7:0] _GEN_4044 = opcode_1 == 4'hf ? _GEN_1994 : _GEN_3530; // @[executor.scala 466:52]
  wire [7:0] _GEN_4045 = opcode_1 == 4'hf ? _GEN_1995 : _GEN_3531; // @[executor.scala 466:52]
  wire [7:0] _GEN_4046 = opcode_1 == 4'hf ? _GEN_1996 : _GEN_3532; // @[executor.scala 466:52]
  wire [7:0] _GEN_4047 = opcode_1 == 4'hf ? _GEN_1997 : _GEN_3533; // @[executor.scala 466:52]
  wire [7:0] _GEN_4048 = opcode_1 == 4'hf ? _GEN_1998 : _GEN_3534; // @[executor.scala 466:52]
  wire [7:0] _GEN_4049 = opcode_1 == 4'hf ? _GEN_1999 : _GEN_3535; // @[executor.scala 466:52]
  wire [7:0] _GEN_4050 = opcode_1 == 4'hf ? _GEN_2000 : _GEN_3536; // @[executor.scala 466:52]
  wire [7:0] _GEN_4051 = opcode_1 == 4'hf ? _GEN_2001 : _GEN_3537; // @[executor.scala 466:52]
  wire [7:0] _GEN_4052 = opcode_1 == 4'hf ? _GEN_2002 : _GEN_3538; // @[executor.scala 466:52]
  wire [7:0] _GEN_4053 = opcode_1 == 4'hf ? _GEN_2003 : _GEN_3539; // @[executor.scala 466:52]
  wire [7:0] _GEN_4054 = opcode_1 == 4'hf ? _GEN_2004 : _GEN_3540; // @[executor.scala 466:52]
  wire [7:0] _GEN_4055 = opcode_1 == 4'hf ? _GEN_2005 : _GEN_3541; // @[executor.scala 466:52]
  wire [7:0] _GEN_4056 = opcode_1 == 4'hf ? _GEN_2006 : _GEN_3542; // @[executor.scala 466:52]
  wire [7:0] _GEN_4057 = opcode_1 == 4'hf ? _GEN_2007 : _GEN_3543; // @[executor.scala 466:52]
  wire [7:0] _GEN_4058 = opcode_1 == 4'hf ? _GEN_2008 : _GEN_3544; // @[executor.scala 466:52]
  wire [7:0] _GEN_4059 = opcode_1 == 4'hf ? _GEN_2009 : _GEN_3545; // @[executor.scala 466:52]
  wire [7:0] _GEN_4060 = opcode_1 == 4'hf ? _GEN_2010 : _GEN_3546; // @[executor.scala 466:52]
  wire [7:0] _GEN_4061 = opcode_1 == 4'hf ? _GEN_2011 : _GEN_3547; // @[executor.scala 466:52]
  wire [7:0] _GEN_4062 = opcode_1 == 4'hf ? _GEN_2012 : _GEN_3548; // @[executor.scala 466:52]
  wire [7:0] _GEN_4063 = opcode_1 == 4'hf ? _GEN_2013 : _GEN_3549; // @[executor.scala 466:52]
  wire [7:0] _GEN_4064 = opcode_1 == 4'hf ? _GEN_2014 : _GEN_3550; // @[executor.scala 466:52]
  wire [7:0] _GEN_4065 = opcode_1 == 4'hf ? _GEN_2015 : _GEN_3551; // @[executor.scala 466:52]
  wire [7:0] _GEN_4066 = opcode_1 == 4'hf ? _GEN_2016 : _GEN_3552; // @[executor.scala 466:52]
  wire [7:0] _GEN_4067 = opcode_1 == 4'hf ? _GEN_2017 : _GEN_3553; // @[executor.scala 466:52]
  wire [7:0] _GEN_4068 = opcode_1 == 4'hf ? _GEN_2018 : _GEN_3554; // @[executor.scala 466:52]
  wire [7:0] _GEN_4069 = opcode_1 == 4'hf ? _GEN_2019 : _GEN_3555; // @[executor.scala 466:52]
  wire [7:0] _GEN_4070 = opcode_1 == 4'hf ? _GEN_2020 : _GEN_3556; // @[executor.scala 466:52]
  wire [7:0] _GEN_4071 = opcode_1 == 4'hf ? _GEN_2021 : _GEN_3557; // @[executor.scala 466:52]
  wire [7:0] _GEN_4072 = opcode_1 == 4'hf ? _GEN_2022 : _GEN_3558; // @[executor.scala 466:52]
  wire [7:0] _GEN_4073 = opcode_1 == 4'hf ? _GEN_2023 : _GEN_3559; // @[executor.scala 466:52]
  wire [7:0] _GEN_4074 = opcode_1 == 4'hf ? _GEN_2024 : _GEN_3560; // @[executor.scala 466:52]
  wire [7:0] _GEN_4075 = opcode_1 == 4'hf ? _GEN_2025 : _GEN_3561; // @[executor.scala 466:52]
  wire [7:0] _GEN_4076 = opcode_1 == 4'hf ? _GEN_2026 : _GEN_3562; // @[executor.scala 466:52]
  wire [7:0] _GEN_4077 = opcode_1 == 4'hf ? _GEN_2027 : _GEN_3563; // @[executor.scala 466:52]
  wire [7:0] _GEN_4078 = opcode_1 == 4'hf ? _GEN_2028 : _GEN_3564; // @[executor.scala 466:52]
  wire [7:0] _GEN_4079 = opcode_1 == 4'hf ? _GEN_2029 : _GEN_3565; // @[executor.scala 466:52]
  wire [7:0] _GEN_4080 = opcode_1 == 4'hf ? _GEN_2030 : _GEN_3566; // @[executor.scala 466:52]
  wire [7:0] _GEN_4081 = opcode_1 == 4'hf ? _GEN_2031 : _GEN_3567; // @[executor.scala 466:52]
  wire [7:0] _GEN_4082 = opcode_1 == 4'hf ? _GEN_2032 : _GEN_3568; // @[executor.scala 466:52]
  wire [7:0] _GEN_4083 = opcode_1 == 4'hf ? _GEN_2033 : _GEN_3569; // @[executor.scala 466:52]
  wire [7:0] _GEN_4084 = opcode_1 == 4'hf ? _GEN_2034 : _GEN_3570; // @[executor.scala 466:52]
  wire [7:0] _GEN_4085 = opcode_1 == 4'hf ? _GEN_2035 : _GEN_3571; // @[executor.scala 466:52]
  wire [7:0] _GEN_4086 = opcode_1 == 4'hf ? _GEN_2036 : _GEN_3572; // @[executor.scala 466:52]
  wire [7:0] _GEN_4087 = opcode_1 == 4'hf ? _GEN_2037 : _GEN_3573; // @[executor.scala 466:52]
  wire [7:0] _GEN_4088 = opcode_1 == 4'hf ? _GEN_2038 : _GEN_3574; // @[executor.scala 466:52]
  wire [7:0] _GEN_4089 = opcode_1 == 4'hf ? _GEN_2039 : _GEN_3575; // @[executor.scala 466:52]
  wire [7:0] _GEN_4090 = opcode_1 == 4'hf ? _GEN_2040 : _GEN_3576; // @[executor.scala 466:52]
  wire [7:0] _GEN_4091 = opcode_1 == 4'hf ? _GEN_2041 : _GEN_3577; // @[executor.scala 466:52]
  wire [7:0] _GEN_4092 = opcode_1 == 4'hf ? _GEN_2042 : _GEN_3578; // @[executor.scala 466:52]
  wire [7:0] _GEN_4093 = opcode_1 == 4'hf ? _GEN_2043 : _GEN_3579; // @[executor.scala 466:52]
  wire [7:0] _GEN_4094 = opcode_1 == 4'hf ? _GEN_2044 : _GEN_3580; // @[executor.scala 466:52]
  wire [7:0] _GEN_4095 = opcode_1 == 4'hf ? _GEN_2045 : _GEN_3581; // @[executor.scala 466:52]
  wire [7:0] _GEN_4096 = opcode_1 == 4'hf ? _GEN_2046 : _GEN_3582; // @[executor.scala 466:52]
  wire [7:0] _GEN_4097 = opcode_1 == 4'hf ? _GEN_2047 : _GEN_3583; // @[executor.scala 466:52]
  wire [7:0] _GEN_4098 = opcode_1 == 4'hf ? _GEN_2048 : _GEN_3584; // @[executor.scala 466:52]
  wire [7:0] _GEN_4099 = opcode_1 == 4'hf ? _GEN_2049 : _GEN_3585; // @[executor.scala 466:52]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_2 = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_8970 = {{2'd0}, dst_offset_2}; // @[executor.scala 473:49]
  wire [7:0] byte_1024 = field_2[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4100 = mask_2[0] ? byte_1024 : _GEN_3588; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1025 = field_2[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4101 = mask_2[1] ? byte_1025 : _GEN_3589; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1026 = field_2[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4102 = mask_2[2] ? byte_1026 : _GEN_3590; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1027 = field_2[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_4103 = mask_2[3] ? byte_1027 : _GEN_3591; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4104 = _GEN_8970 == 8'h0 ? _GEN_4100 : _GEN_3588; // @[executor.scala 473:84]
  wire [7:0] _GEN_4105 = _GEN_8970 == 8'h0 ? _GEN_4101 : _GEN_3589; // @[executor.scala 473:84]
  wire [7:0] _GEN_4106 = _GEN_8970 == 8'h0 ? _GEN_4102 : _GEN_3590; // @[executor.scala 473:84]
  wire [7:0] _GEN_4107 = _GEN_8970 == 8'h0 ? _GEN_4103 : _GEN_3591; // @[executor.scala 473:84]
  wire [7:0] _GEN_4108 = mask_2[0] ? byte_1024 : _GEN_3592; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4109 = mask_2[1] ? byte_1025 : _GEN_3593; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4110 = mask_2[2] ? byte_1026 : _GEN_3594; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4111 = mask_2[3] ? byte_1027 : _GEN_3595; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4112 = _GEN_8970 == 8'h1 ? _GEN_4108 : _GEN_3592; // @[executor.scala 473:84]
  wire [7:0] _GEN_4113 = _GEN_8970 == 8'h1 ? _GEN_4109 : _GEN_3593; // @[executor.scala 473:84]
  wire [7:0] _GEN_4114 = _GEN_8970 == 8'h1 ? _GEN_4110 : _GEN_3594; // @[executor.scala 473:84]
  wire [7:0] _GEN_4115 = _GEN_8970 == 8'h1 ? _GEN_4111 : _GEN_3595; // @[executor.scala 473:84]
  wire [7:0] _GEN_4116 = mask_2[0] ? byte_1024 : _GEN_3596; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4117 = mask_2[1] ? byte_1025 : _GEN_3597; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4118 = mask_2[2] ? byte_1026 : _GEN_3598; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4119 = mask_2[3] ? byte_1027 : _GEN_3599; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4120 = _GEN_8970 == 8'h2 ? _GEN_4116 : _GEN_3596; // @[executor.scala 473:84]
  wire [7:0] _GEN_4121 = _GEN_8970 == 8'h2 ? _GEN_4117 : _GEN_3597; // @[executor.scala 473:84]
  wire [7:0] _GEN_4122 = _GEN_8970 == 8'h2 ? _GEN_4118 : _GEN_3598; // @[executor.scala 473:84]
  wire [7:0] _GEN_4123 = _GEN_8970 == 8'h2 ? _GEN_4119 : _GEN_3599; // @[executor.scala 473:84]
  wire [7:0] _GEN_4124 = mask_2[0] ? byte_1024 : _GEN_3600; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4125 = mask_2[1] ? byte_1025 : _GEN_3601; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4126 = mask_2[2] ? byte_1026 : _GEN_3602; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4127 = mask_2[3] ? byte_1027 : _GEN_3603; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4128 = _GEN_8970 == 8'h3 ? _GEN_4124 : _GEN_3600; // @[executor.scala 473:84]
  wire [7:0] _GEN_4129 = _GEN_8970 == 8'h3 ? _GEN_4125 : _GEN_3601; // @[executor.scala 473:84]
  wire [7:0] _GEN_4130 = _GEN_8970 == 8'h3 ? _GEN_4126 : _GEN_3602; // @[executor.scala 473:84]
  wire [7:0] _GEN_4131 = _GEN_8970 == 8'h3 ? _GEN_4127 : _GEN_3603; // @[executor.scala 473:84]
  wire [7:0] _GEN_4132 = mask_2[0] ? byte_1024 : _GEN_3604; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4133 = mask_2[1] ? byte_1025 : _GEN_3605; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4134 = mask_2[2] ? byte_1026 : _GEN_3606; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4135 = mask_2[3] ? byte_1027 : _GEN_3607; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4136 = _GEN_8970 == 8'h4 ? _GEN_4132 : _GEN_3604; // @[executor.scala 473:84]
  wire [7:0] _GEN_4137 = _GEN_8970 == 8'h4 ? _GEN_4133 : _GEN_3605; // @[executor.scala 473:84]
  wire [7:0] _GEN_4138 = _GEN_8970 == 8'h4 ? _GEN_4134 : _GEN_3606; // @[executor.scala 473:84]
  wire [7:0] _GEN_4139 = _GEN_8970 == 8'h4 ? _GEN_4135 : _GEN_3607; // @[executor.scala 473:84]
  wire [7:0] _GEN_4140 = mask_2[0] ? byte_1024 : _GEN_3608; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4141 = mask_2[1] ? byte_1025 : _GEN_3609; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4142 = mask_2[2] ? byte_1026 : _GEN_3610; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4143 = mask_2[3] ? byte_1027 : _GEN_3611; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4144 = _GEN_8970 == 8'h5 ? _GEN_4140 : _GEN_3608; // @[executor.scala 473:84]
  wire [7:0] _GEN_4145 = _GEN_8970 == 8'h5 ? _GEN_4141 : _GEN_3609; // @[executor.scala 473:84]
  wire [7:0] _GEN_4146 = _GEN_8970 == 8'h5 ? _GEN_4142 : _GEN_3610; // @[executor.scala 473:84]
  wire [7:0] _GEN_4147 = _GEN_8970 == 8'h5 ? _GEN_4143 : _GEN_3611; // @[executor.scala 473:84]
  wire [7:0] _GEN_4148 = mask_2[0] ? byte_1024 : _GEN_3612; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4149 = mask_2[1] ? byte_1025 : _GEN_3613; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4150 = mask_2[2] ? byte_1026 : _GEN_3614; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4151 = mask_2[3] ? byte_1027 : _GEN_3615; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4152 = _GEN_8970 == 8'h6 ? _GEN_4148 : _GEN_3612; // @[executor.scala 473:84]
  wire [7:0] _GEN_4153 = _GEN_8970 == 8'h6 ? _GEN_4149 : _GEN_3613; // @[executor.scala 473:84]
  wire [7:0] _GEN_4154 = _GEN_8970 == 8'h6 ? _GEN_4150 : _GEN_3614; // @[executor.scala 473:84]
  wire [7:0] _GEN_4155 = _GEN_8970 == 8'h6 ? _GEN_4151 : _GEN_3615; // @[executor.scala 473:84]
  wire [7:0] _GEN_4156 = mask_2[0] ? byte_1024 : _GEN_3616; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4157 = mask_2[1] ? byte_1025 : _GEN_3617; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4158 = mask_2[2] ? byte_1026 : _GEN_3618; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4159 = mask_2[3] ? byte_1027 : _GEN_3619; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4160 = _GEN_8970 == 8'h7 ? _GEN_4156 : _GEN_3616; // @[executor.scala 473:84]
  wire [7:0] _GEN_4161 = _GEN_8970 == 8'h7 ? _GEN_4157 : _GEN_3617; // @[executor.scala 473:84]
  wire [7:0] _GEN_4162 = _GEN_8970 == 8'h7 ? _GEN_4158 : _GEN_3618; // @[executor.scala 473:84]
  wire [7:0] _GEN_4163 = _GEN_8970 == 8'h7 ? _GEN_4159 : _GEN_3619; // @[executor.scala 473:84]
  wire [7:0] _GEN_4164 = mask_2[0] ? byte_1024 : _GEN_3620; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4165 = mask_2[1] ? byte_1025 : _GEN_3621; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4166 = mask_2[2] ? byte_1026 : _GEN_3622; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4167 = mask_2[3] ? byte_1027 : _GEN_3623; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4168 = _GEN_8970 == 8'h8 ? _GEN_4164 : _GEN_3620; // @[executor.scala 473:84]
  wire [7:0] _GEN_4169 = _GEN_8970 == 8'h8 ? _GEN_4165 : _GEN_3621; // @[executor.scala 473:84]
  wire [7:0] _GEN_4170 = _GEN_8970 == 8'h8 ? _GEN_4166 : _GEN_3622; // @[executor.scala 473:84]
  wire [7:0] _GEN_4171 = _GEN_8970 == 8'h8 ? _GEN_4167 : _GEN_3623; // @[executor.scala 473:84]
  wire [7:0] _GEN_4172 = mask_2[0] ? byte_1024 : _GEN_3624; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4173 = mask_2[1] ? byte_1025 : _GEN_3625; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4174 = mask_2[2] ? byte_1026 : _GEN_3626; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4175 = mask_2[3] ? byte_1027 : _GEN_3627; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4176 = _GEN_8970 == 8'h9 ? _GEN_4172 : _GEN_3624; // @[executor.scala 473:84]
  wire [7:0] _GEN_4177 = _GEN_8970 == 8'h9 ? _GEN_4173 : _GEN_3625; // @[executor.scala 473:84]
  wire [7:0] _GEN_4178 = _GEN_8970 == 8'h9 ? _GEN_4174 : _GEN_3626; // @[executor.scala 473:84]
  wire [7:0] _GEN_4179 = _GEN_8970 == 8'h9 ? _GEN_4175 : _GEN_3627; // @[executor.scala 473:84]
  wire [7:0] _GEN_4180 = mask_2[0] ? byte_1024 : _GEN_3628; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4181 = mask_2[1] ? byte_1025 : _GEN_3629; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4182 = mask_2[2] ? byte_1026 : _GEN_3630; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4183 = mask_2[3] ? byte_1027 : _GEN_3631; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4184 = _GEN_8970 == 8'ha ? _GEN_4180 : _GEN_3628; // @[executor.scala 473:84]
  wire [7:0] _GEN_4185 = _GEN_8970 == 8'ha ? _GEN_4181 : _GEN_3629; // @[executor.scala 473:84]
  wire [7:0] _GEN_4186 = _GEN_8970 == 8'ha ? _GEN_4182 : _GEN_3630; // @[executor.scala 473:84]
  wire [7:0] _GEN_4187 = _GEN_8970 == 8'ha ? _GEN_4183 : _GEN_3631; // @[executor.scala 473:84]
  wire [7:0] _GEN_4188 = mask_2[0] ? byte_1024 : _GEN_3632; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4189 = mask_2[1] ? byte_1025 : _GEN_3633; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4190 = mask_2[2] ? byte_1026 : _GEN_3634; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4191 = mask_2[3] ? byte_1027 : _GEN_3635; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4192 = _GEN_8970 == 8'hb ? _GEN_4188 : _GEN_3632; // @[executor.scala 473:84]
  wire [7:0] _GEN_4193 = _GEN_8970 == 8'hb ? _GEN_4189 : _GEN_3633; // @[executor.scala 473:84]
  wire [7:0] _GEN_4194 = _GEN_8970 == 8'hb ? _GEN_4190 : _GEN_3634; // @[executor.scala 473:84]
  wire [7:0] _GEN_4195 = _GEN_8970 == 8'hb ? _GEN_4191 : _GEN_3635; // @[executor.scala 473:84]
  wire [7:0] _GEN_4196 = mask_2[0] ? byte_1024 : _GEN_3636; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4197 = mask_2[1] ? byte_1025 : _GEN_3637; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4198 = mask_2[2] ? byte_1026 : _GEN_3638; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4199 = mask_2[3] ? byte_1027 : _GEN_3639; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4200 = _GEN_8970 == 8'hc ? _GEN_4196 : _GEN_3636; // @[executor.scala 473:84]
  wire [7:0] _GEN_4201 = _GEN_8970 == 8'hc ? _GEN_4197 : _GEN_3637; // @[executor.scala 473:84]
  wire [7:0] _GEN_4202 = _GEN_8970 == 8'hc ? _GEN_4198 : _GEN_3638; // @[executor.scala 473:84]
  wire [7:0] _GEN_4203 = _GEN_8970 == 8'hc ? _GEN_4199 : _GEN_3639; // @[executor.scala 473:84]
  wire [7:0] _GEN_4204 = mask_2[0] ? byte_1024 : _GEN_3640; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4205 = mask_2[1] ? byte_1025 : _GEN_3641; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4206 = mask_2[2] ? byte_1026 : _GEN_3642; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4207 = mask_2[3] ? byte_1027 : _GEN_3643; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4208 = _GEN_8970 == 8'hd ? _GEN_4204 : _GEN_3640; // @[executor.scala 473:84]
  wire [7:0] _GEN_4209 = _GEN_8970 == 8'hd ? _GEN_4205 : _GEN_3641; // @[executor.scala 473:84]
  wire [7:0] _GEN_4210 = _GEN_8970 == 8'hd ? _GEN_4206 : _GEN_3642; // @[executor.scala 473:84]
  wire [7:0] _GEN_4211 = _GEN_8970 == 8'hd ? _GEN_4207 : _GEN_3643; // @[executor.scala 473:84]
  wire [7:0] _GEN_4212 = mask_2[0] ? byte_1024 : _GEN_3644; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4213 = mask_2[1] ? byte_1025 : _GEN_3645; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4214 = mask_2[2] ? byte_1026 : _GEN_3646; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4215 = mask_2[3] ? byte_1027 : _GEN_3647; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4216 = _GEN_8970 == 8'he ? _GEN_4212 : _GEN_3644; // @[executor.scala 473:84]
  wire [7:0] _GEN_4217 = _GEN_8970 == 8'he ? _GEN_4213 : _GEN_3645; // @[executor.scala 473:84]
  wire [7:0] _GEN_4218 = _GEN_8970 == 8'he ? _GEN_4214 : _GEN_3646; // @[executor.scala 473:84]
  wire [7:0] _GEN_4219 = _GEN_8970 == 8'he ? _GEN_4215 : _GEN_3647; // @[executor.scala 473:84]
  wire [7:0] _GEN_4220 = mask_2[0] ? byte_1024 : _GEN_3648; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4221 = mask_2[1] ? byte_1025 : _GEN_3649; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4222 = mask_2[2] ? byte_1026 : _GEN_3650; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4223 = mask_2[3] ? byte_1027 : _GEN_3651; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4224 = _GEN_8970 == 8'hf ? _GEN_4220 : _GEN_3648; // @[executor.scala 473:84]
  wire [7:0] _GEN_4225 = _GEN_8970 == 8'hf ? _GEN_4221 : _GEN_3649; // @[executor.scala 473:84]
  wire [7:0] _GEN_4226 = _GEN_8970 == 8'hf ? _GEN_4222 : _GEN_3650; // @[executor.scala 473:84]
  wire [7:0] _GEN_4227 = _GEN_8970 == 8'hf ? _GEN_4223 : _GEN_3651; // @[executor.scala 473:84]
  wire [7:0] _GEN_4228 = mask_2[0] ? byte_1024 : _GEN_3652; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4229 = mask_2[1] ? byte_1025 : _GEN_3653; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4230 = mask_2[2] ? byte_1026 : _GEN_3654; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4231 = mask_2[3] ? byte_1027 : _GEN_3655; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4232 = _GEN_8970 == 8'h10 ? _GEN_4228 : _GEN_3652; // @[executor.scala 473:84]
  wire [7:0] _GEN_4233 = _GEN_8970 == 8'h10 ? _GEN_4229 : _GEN_3653; // @[executor.scala 473:84]
  wire [7:0] _GEN_4234 = _GEN_8970 == 8'h10 ? _GEN_4230 : _GEN_3654; // @[executor.scala 473:84]
  wire [7:0] _GEN_4235 = _GEN_8970 == 8'h10 ? _GEN_4231 : _GEN_3655; // @[executor.scala 473:84]
  wire [7:0] _GEN_4236 = mask_2[0] ? byte_1024 : _GEN_3656; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4237 = mask_2[1] ? byte_1025 : _GEN_3657; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4238 = mask_2[2] ? byte_1026 : _GEN_3658; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4239 = mask_2[3] ? byte_1027 : _GEN_3659; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4240 = _GEN_8970 == 8'h11 ? _GEN_4236 : _GEN_3656; // @[executor.scala 473:84]
  wire [7:0] _GEN_4241 = _GEN_8970 == 8'h11 ? _GEN_4237 : _GEN_3657; // @[executor.scala 473:84]
  wire [7:0] _GEN_4242 = _GEN_8970 == 8'h11 ? _GEN_4238 : _GEN_3658; // @[executor.scala 473:84]
  wire [7:0] _GEN_4243 = _GEN_8970 == 8'h11 ? _GEN_4239 : _GEN_3659; // @[executor.scala 473:84]
  wire [7:0] _GEN_4244 = mask_2[0] ? byte_1024 : _GEN_3660; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4245 = mask_2[1] ? byte_1025 : _GEN_3661; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4246 = mask_2[2] ? byte_1026 : _GEN_3662; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4247 = mask_2[3] ? byte_1027 : _GEN_3663; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4248 = _GEN_8970 == 8'h12 ? _GEN_4244 : _GEN_3660; // @[executor.scala 473:84]
  wire [7:0] _GEN_4249 = _GEN_8970 == 8'h12 ? _GEN_4245 : _GEN_3661; // @[executor.scala 473:84]
  wire [7:0] _GEN_4250 = _GEN_8970 == 8'h12 ? _GEN_4246 : _GEN_3662; // @[executor.scala 473:84]
  wire [7:0] _GEN_4251 = _GEN_8970 == 8'h12 ? _GEN_4247 : _GEN_3663; // @[executor.scala 473:84]
  wire [7:0] _GEN_4252 = mask_2[0] ? byte_1024 : _GEN_3664; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4253 = mask_2[1] ? byte_1025 : _GEN_3665; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4254 = mask_2[2] ? byte_1026 : _GEN_3666; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4255 = mask_2[3] ? byte_1027 : _GEN_3667; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4256 = _GEN_8970 == 8'h13 ? _GEN_4252 : _GEN_3664; // @[executor.scala 473:84]
  wire [7:0] _GEN_4257 = _GEN_8970 == 8'h13 ? _GEN_4253 : _GEN_3665; // @[executor.scala 473:84]
  wire [7:0] _GEN_4258 = _GEN_8970 == 8'h13 ? _GEN_4254 : _GEN_3666; // @[executor.scala 473:84]
  wire [7:0] _GEN_4259 = _GEN_8970 == 8'h13 ? _GEN_4255 : _GEN_3667; // @[executor.scala 473:84]
  wire [7:0] _GEN_4260 = mask_2[0] ? byte_1024 : _GEN_3668; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4261 = mask_2[1] ? byte_1025 : _GEN_3669; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4262 = mask_2[2] ? byte_1026 : _GEN_3670; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4263 = mask_2[3] ? byte_1027 : _GEN_3671; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4264 = _GEN_8970 == 8'h14 ? _GEN_4260 : _GEN_3668; // @[executor.scala 473:84]
  wire [7:0] _GEN_4265 = _GEN_8970 == 8'h14 ? _GEN_4261 : _GEN_3669; // @[executor.scala 473:84]
  wire [7:0] _GEN_4266 = _GEN_8970 == 8'h14 ? _GEN_4262 : _GEN_3670; // @[executor.scala 473:84]
  wire [7:0] _GEN_4267 = _GEN_8970 == 8'h14 ? _GEN_4263 : _GEN_3671; // @[executor.scala 473:84]
  wire [7:0] _GEN_4268 = mask_2[0] ? byte_1024 : _GEN_3672; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4269 = mask_2[1] ? byte_1025 : _GEN_3673; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4270 = mask_2[2] ? byte_1026 : _GEN_3674; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4271 = mask_2[3] ? byte_1027 : _GEN_3675; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4272 = _GEN_8970 == 8'h15 ? _GEN_4268 : _GEN_3672; // @[executor.scala 473:84]
  wire [7:0] _GEN_4273 = _GEN_8970 == 8'h15 ? _GEN_4269 : _GEN_3673; // @[executor.scala 473:84]
  wire [7:0] _GEN_4274 = _GEN_8970 == 8'h15 ? _GEN_4270 : _GEN_3674; // @[executor.scala 473:84]
  wire [7:0] _GEN_4275 = _GEN_8970 == 8'h15 ? _GEN_4271 : _GEN_3675; // @[executor.scala 473:84]
  wire [7:0] _GEN_4276 = mask_2[0] ? byte_1024 : _GEN_3676; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4277 = mask_2[1] ? byte_1025 : _GEN_3677; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4278 = mask_2[2] ? byte_1026 : _GEN_3678; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4279 = mask_2[3] ? byte_1027 : _GEN_3679; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4280 = _GEN_8970 == 8'h16 ? _GEN_4276 : _GEN_3676; // @[executor.scala 473:84]
  wire [7:0] _GEN_4281 = _GEN_8970 == 8'h16 ? _GEN_4277 : _GEN_3677; // @[executor.scala 473:84]
  wire [7:0] _GEN_4282 = _GEN_8970 == 8'h16 ? _GEN_4278 : _GEN_3678; // @[executor.scala 473:84]
  wire [7:0] _GEN_4283 = _GEN_8970 == 8'h16 ? _GEN_4279 : _GEN_3679; // @[executor.scala 473:84]
  wire [7:0] _GEN_4284 = mask_2[0] ? byte_1024 : _GEN_3680; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4285 = mask_2[1] ? byte_1025 : _GEN_3681; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4286 = mask_2[2] ? byte_1026 : _GEN_3682; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4287 = mask_2[3] ? byte_1027 : _GEN_3683; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4288 = _GEN_8970 == 8'h17 ? _GEN_4284 : _GEN_3680; // @[executor.scala 473:84]
  wire [7:0] _GEN_4289 = _GEN_8970 == 8'h17 ? _GEN_4285 : _GEN_3681; // @[executor.scala 473:84]
  wire [7:0] _GEN_4290 = _GEN_8970 == 8'h17 ? _GEN_4286 : _GEN_3682; // @[executor.scala 473:84]
  wire [7:0] _GEN_4291 = _GEN_8970 == 8'h17 ? _GEN_4287 : _GEN_3683; // @[executor.scala 473:84]
  wire [7:0] _GEN_4292 = mask_2[0] ? byte_1024 : _GEN_3684; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4293 = mask_2[1] ? byte_1025 : _GEN_3685; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4294 = mask_2[2] ? byte_1026 : _GEN_3686; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4295 = mask_2[3] ? byte_1027 : _GEN_3687; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4296 = _GEN_8970 == 8'h18 ? _GEN_4292 : _GEN_3684; // @[executor.scala 473:84]
  wire [7:0] _GEN_4297 = _GEN_8970 == 8'h18 ? _GEN_4293 : _GEN_3685; // @[executor.scala 473:84]
  wire [7:0] _GEN_4298 = _GEN_8970 == 8'h18 ? _GEN_4294 : _GEN_3686; // @[executor.scala 473:84]
  wire [7:0] _GEN_4299 = _GEN_8970 == 8'h18 ? _GEN_4295 : _GEN_3687; // @[executor.scala 473:84]
  wire [7:0] _GEN_4300 = mask_2[0] ? byte_1024 : _GEN_3688; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4301 = mask_2[1] ? byte_1025 : _GEN_3689; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4302 = mask_2[2] ? byte_1026 : _GEN_3690; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4303 = mask_2[3] ? byte_1027 : _GEN_3691; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4304 = _GEN_8970 == 8'h19 ? _GEN_4300 : _GEN_3688; // @[executor.scala 473:84]
  wire [7:0] _GEN_4305 = _GEN_8970 == 8'h19 ? _GEN_4301 : _GEN_3689; // @[executor.scala 473:84]
  wire [7:0] _GEN_4306 = _GEN_8970 == 8'h19 ? _GEN_4302 : _GEN_3690; // @[executor.scala 473:84]
  wire [7:0] _GEN_4307 = _GEN_8970 == 8'h19 ? _GEN_4303 : _GEN_3691; // @[executor.scala 473:84]
  wire [7:0] _GEN_4308 = mask_2[0] ? byte_1024 : _GEN_3692; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4309 = mask_2[1] ? byte_1025 : _GEN_3693; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4310 = mask_2[2] ? byte_1026 : _GEN_3694; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4311 = mask_2[3] ? byte_1027 : _GEN_3695; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4312 = _GEN_8970 == 8'h1a ? _GEN_4308 : _GEN_3692; // @[executor.scala 473:84]
  wire [7:0] _GEN_4313 = _GEN_8970 == 8'h1a ? _GEN_4309 : _GEN_3693; // @[executor.scala 473:84]
  wire [7:0] _GEN_4314 = _GEN_8970 == 8'h1a ? _GEN_4310 : _GEN_3694; // @[executor.scala 473:84]
  wire [7:0] _GEN_4315 = _GEN_8970 == 8'h1a ? _GEN_4311 : _GEN_3695; // @[executor.scala 473:84]
  wire [7:0] _GEN_4316 = mask_2[0] ? byte_1024 : _GEN_3696; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4317 = mask_2[1] ? byte_1025 : _GEN_3697; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4318 = mask_2[2] ? byte_1026 : _GEN_3698; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4319 = mask_2[3] ? byte_1027 : _GEN_3699; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4320 = _GEN_8970 == 8'h1b ? _GEN_4316 : _GEN_3696; // @[executor.scala 473:84]
  wire [7:0] _GEN_4321 = _GEN_8970 == 8'h1b ? _GEN_4317 : _GEN_3697; // @[executor.scala 473:84]
  wire [7:0] _GEN_4322 = _GEN_8970 == 8'h1b ? _GEN_4318 : _GEN_3698; // @[executor.scala 473:84]
  wire [7:0] _GEN_4323 = _GEN_8970 == 8'h1b ? _GEN_4319 : _GEN_3699; // @[executor.scala 473:84]
  wire [7:0] _GEN_4324 = mask_2[0] ? byte_1024 : _GEN_3700; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4325 = mask_2[1] ? byte_1025 : _GEN_3701; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4326 = mask_2[2] ? byte_1026 : _GEN_3702; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4327 = mask_2[3] ? byte_1027 : _GEN_3703; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4328 = _GEN_8970 == 8'h1c ? _GEN_4324 : _GEN_3700; // @[executor.scala 473:84]
  wire [7:0] _GEN_4329 = _GEN_8970 == 8'h1c ? _GEN_4325 : _GEN_3701; // @[executor.scala 473:84]
  wire [7:0] _GEN_4330 = _GEN_8970 == 8'h1c ? _GEN_4326 : _GEN_3702; // @[executor.scala 473:84]
  wire [7:0] _GEN_4331 = _GEN_8970 == 8'h1c ? _GEN_4327 : _GEN_3703; // @[executor.scala 473:84]
  wire [7:0] _GEN_4332 = mask_2[0] ? byte_1024 : _GEN_3704; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4333 = mask_2[1] ? byte_1025 : _GEN_3705; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4334 = mask_2[2] ? byte_1026 : _GEN_3706; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4335 = mask_2[3] ? byte_1027 : _GEN_3707; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4336 = _GEN_8970 == 8'h1d ? _GEN_4332 : _GEN_3704; // @[executor.scala 473:84]
  wire [7:0] _GEN_4337 = _GEN_8970 == 8'h1d ? _GEN_4333 : _GEN_3705; // @[executor.scala 473:84]
  wire [7:0] _GEN_4338 = _GEN_8970 == 8'h1d ? _GEN_4334 : _GEN_3706; // @[executor.scala 473:84]
  wire [7:0] _GEN_4339 = _GEN_8970 == 8'h1d ? _GEN_4335 : _GEN_3707; // @[executor.scala 473:84]
  wire [7:0] _GEN_4340 = mask_2[0] ? byte_1024 : _GEN_3708; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4341 = mask_2[1] ? byte_1025 : _GEN_3709; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4342 = mask_2[2] ? byte_1026 : _GEN_3710; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4343 = mask_2[3] ? byte_1027 : _GEN_3711; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4344 = _GEN_8970 == 8'h1e ? _GEN_4340 : _GEN_3708; // @[executor.scala 473:84]
  wire [7:0] _GEN_4345 = _GEN_8970 == 8'h1e ? _GEN_4341 : _GEN_3709; // @[executor.scala 473:84]
  wire [7:0] _GEN_4346 = _GEN_8970 == 8'h1e ? _GEN_4342 : _GEN_3710; // @[executor.scala 473:84]
  wire [7:0] _GEN_4347 = _GEN_8970 == 8'h1e ? _GEN_4343 : _GEN_3711; // @[executor.scala 473:84]
  wire [7:0] _GEN_4348 = mask_2[0] ? byte_1024 : _GEN_3712; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4349 = mask_2[1] ? byte_1025 : _GEN_3713; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4350 = mask_2[2] ? byte_1026 : _GEN_3714; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4351 = mask_2[3] ? byte_1027 : _GEN_3715; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4352 = _GEN_8970 == 8'h1f ? _GEN_4348 : _GEN_3712; // @[executor.scala 473:84]
  wire [7:0] _GEN_4353 = _GEN_8970 == 8'h1f ? _GEN_4349 : _GEN_3713; // @[executor.scala 473:84]
  wire [7:0] _GEN_4354 = _GEN_8970 == 8'h1f ? _GEN_4350 : _GEN_3714; // @[executor.scala 473:84]
  wire [7:0] _GEN_4355 = _GEN_8970 == 8'h1f ? _GEN_4351 : _GEN_3715; // @[executor.scala 473:84]
  wire [7:0] _GEN_4356 = mask_2[0] ? byte_1024 : _GEN_3716; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4357 = mask_2[1] ? byte_1025 : _GEN_3717; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4358 = mask_2[2] ? byte_1026 : _GEN_3718; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4359 = mask_2[3] ? byte_1027 : _GEN_3719; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4360 = _GEN_8970 == 8'h20 ? _GEN_4356 : _GEN_3716; // @[executor.scala 473:84]
  wire [7:0] _GEN_4361 = _GEN_8970 == 8'h20 ? _GEN_4357 : _GEN_3717; // @[executor.scala 473:84]
  wire [7:0] _GEN_4362 = _GEN_8970 == 8'h20 ? _GEN_4358 : _GEN_3718; // @[executor.scala 473:84]
  wire [7:0] _GEN_4363 = _GEN_8970 == 8'h20 ? _GEN_4359 : _GEN_3719; // @[executor.scala 473:84]
  wire [7:0] _GEN_4364 = mask_2[0] ? byte_1024 : _GEN_3720; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4365 = mask_2[1] ? byte_1025 : _GEN_3721; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4366 = mask_2[2] ? byte_1026 : _GEN_3722; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4367 = mask_2[3] ? byte_1027 : _GEN_3723; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4368 = _GEN_8970 == 8'h21 ? _GEN_4364 : _GEN_3720; // @[executor.scala 473:84]
  wire [7:0] _GEN_4369 = _GEN_8970 == 8'h21 ? _GEN_4365 : _GEN_3721; // @[executor.scala 473:84]
  wire [7:0] _GEN_4370 = _GEN_8970 == 8'h21 ? _GEN_4366 : _GEN_3722; // @[executor.scala 473:84]
  wire [7:0] _GEN_4371 = _GEN_8970 == 8'h21 ? _GEN_4367 : _GEN_3723; // @[executor.scala 473:84]
  wire [7:0] _GEN_4372 = mask_2[0] ? byte_1024 : _GEN_3724; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4373 = mask_2[1] ? byte_1025 : _GEN_3725; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4374 = mask_2[2] ? byte_1026 : _GEN_3726; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4375 = mask_2[3] ? byte_1027 : _GEN_3727; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4376 = _GEN_8970 == 8'h22 ? _GEN_4372 : _GEN_3724; // @[executor.scala 473:84]
  wire [7:0] _GEN_4377 = _GEN_8970 == 8'h22 ? _GEN_4373 : _GEN_3725; // @[executor.scala 473:84]
  wire [7:0] _GEN_4378 = _GEN_8970 == 8'h22 ? _GEN_4374 : _GEN_3726; // @[executor.scala 473:84]
  wire [7:0] _GEN_4379 = _GEN_8970 == 8'h22 ? _GEN_4375 : _GEN_3727; // @[executor.scala 473:84]
  wire [7:0] _GEN_4380 = mask_2[0] ? byte_1024 : _GEN_3728; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4381 = mask_2[1] ? byte_1025 : _GEN_3729; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4382 = mask_2[2] ? byte_1026 : _GEN_3730; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4383 = mask_2[3] ? byte_1027 : _GEN_3731; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4384 = _GEN_8970 == 8'h23 ? _GEN_4380 : _GEN_3728; // @[executor.scala 473:84]
  wire [7:0] _GEN_4385 = _GEN_8970 == 8'h23 ? _GEN_4381 : _GEN_3729; // @[executor.scala 473:84]
  wire [7:0] _GEN_4386 = _GEN_8970 == 8'h23 ? _GEN_4382 : _GEN_3730; // @[executor.scala 473:84]
  wire [7:0] _GEN_4387 = _GEN_8970 == 8'h23 ? _GEN_4383 : _GEN_3731; // @[executor.scala 473:84]
  wire [7:0] _GEN_4388 = mask_2[0] ? byte_1024 : _GEN_3732; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4389 = mask_2[1] ? byte_1025 : _GEN_3733; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4390 = mask_2[2] ? byte_1026 : _GEN_3734; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4391 = mask_2[3] ? byte_1027 : _GEN_3735; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4392 = _GEN_8970 == 8'h24 ? _GEN_4388 : _GEN_3732; // @[executor.scala 473:84]
  wire [7:0] _GEN_4393 = _GEN_8970 == 8'h24 ? _GEN_4389 : _GEN_3733; // @[executor.scala 473:84]
  wire [7:0] _GEN_4394 = _GEN_8970 == 8'h24 ? _GEN_4390 : _GEN_3734; // @[executor.scala 473:84]
  wire [7:0] _GEN_4395 = _GEN_8970 == 8'h24 ? _GEN_4391 : _GEN_3735; // @[executor.scala 473:84]
  wire [7:0] _GEN_4396 = mask_2[0] ? byte_1024 : _GEN_3736; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4397 = mask_2[1] ? byte_1025 : _GEN_3737; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4398 = mask_2[2] ? byte_1026 : _GEN_3738; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4399 = mask_2[3] ? byte_1027 : _GEN_3739; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4400 = _GEN_8970 == 8'h25 ? _GEN_4396 : _GEN_3736; // @[executor.scala 473:84]
  wire [7:0] _GEN_4401 = _GEN_8970 == 8'h25 ? _GEN_4397 : _GEN_3737; // @[executor.scala 473:84]
  wire [7:0] _GEN_4402 = _GEN_8970 == 8'h25 ? _GEN_4398 : _GEN_3738; // @[executor.scala 473:84]
  wire [7:0] _GEN_4403 = _GEN_8970 == 8'h25 ? _GEN_4399 : _GEN_3739; // @[executor.scala 473:84]
  wire [7:0] _GEN_4404 = mask_2[0] ? byte_1024 : _GEN_3740; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4405 = mask_2[1] ? byte_1025 : _GEN_3741; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4406 = mask_2[2] ? byte_1026 : _GEN_3742; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4407 = mask_2[3] ? byte_1027 : _GEN_3743; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4408 = _GEN_8970 == 8'h26 ? _GEN_4404 : _GEN_3740; // @[executor.scala 473:84]
  wire [7:0] _GEN_4409 = _GEN_8970 == 8'h26 ? _GEN_4405 : _GEN_3741; // @[executor.scala 473:84]
  wire [7:0] _GEN_4410 = _GEN_8970 == 8'h26 ? _GEN_4406 : _GEN_3742; // @[executor.scala 473:84]
  wire [7:0] _GEN_4411 = _GEN_8970 == 8'h26 ? _GEN_4407 : _GEN_3743; // @[executor.scala 473:84]
  wire [7:0] _GEN_4412 = mask_2[0] ? byte_1024 : _GEN_3744; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4413 = mask_2[1] ? byte_1025 : _GEN_3745; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4414 = mask_2[2] ? byte_1026 : _GEN_3746; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4415 = mask_2[3] ? byte_1027 : _GEN_3747; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4416 = _GEN_8970 == 8'h27 ? _GEN_4412 : _GEN_3744; // @[executor.scala 473:84]
  wire [7:0] _GEN_4417 = _GEN_8970 == 8'h27 ? _GEN_4413 : _GEN_3745; // @[executor.scala 473:84]
  wire [7:0] _GEN_4418 = _GEN_8970 == 8'h27 ? _GEN_4414 : _GEN_3746; // @[executor.scala 473:84]
  wire [7:0] _GEN_4419 = _GEN_8970 == 8'h27 ? _GEN_4415 : _GEN_3747; // @[executor.scala 473:84]
  wire [7:0] _GEN_4420 = mask_2[0] ? byte_1024 : _GEN_3748; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4421 = mask_2[1] ? byte_1025 : _GEN_3749; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4422 = mask_2[2] ? byte_1026 : _GEN_3750; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4423 = mask_2[3] ? byte_1027 : _GEN_3751; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4424 = _GEN_8970 == 8'h28 ? _GEN_4420 : _GEN_3748; // @[executor.scala 473:84]
  wire [7:0] _GEN_4425 = _GEN_8970 == 8'h28 ? _GEN_4421 : _GEN_3749; // @[executor.scala 473:84]
  wire [7:0] _GEN_4426 = _GEN_8970 == 8'h28 ? _GEN_4422 : _GEN_3750; // @[executor.scala 473:84]
  wire [7:0] _GEN_4427 = _GEN_8970 == 8'h28 ? _GEN_4423 : _GEN_3751; // @[executor.scala 473:84]
  wire [7:0] _GEN_4428 = mask_2[0] ? byte_1024 : _GEN_3752; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4429 = mask_2[1] ? byte_1025 : _GEN_3753; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4430 = mask_2[2] ? byte_1026 : _GEN_3754; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4431 = mask_2[3] ? byte_1027 : _GEN_3755; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4432 = _GEN_8970 == 8'h29 ? _GEN_4428 : _GEN_3752; // @[executor.scala 473:84]
  wire [7:0] _GEN_4433 = _GEN_8970 == 8'h29 ? _GEN_4429 : _GEN_3753; // @[executor.scala 473:84]
  wire [7:0] _GEN_4434 = _GEN_8970 == 8'h29 ? _GEN_4430 : _GEN_3754; // @[executor.scala 473:84]
  wire [7:0] _GEN_4435 = _GEN_8970 == 8'h29 ? _GEN_4431 : _GEN_3755; // @[executor.scala 473:84]
  wire [7:0] _GEN_4436 = mask_2[0] ? byte_1024 : _GEN_3756; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4437 = mask_2[1] ? byte_1025 : _GEN_3757; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4438 = mask_2[2] ? byte_1026 : _GEN_3758; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4439 = mask_2[3] ? byte_1027 : _GEN_3759; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4440 = _GEN_8970 == 8'h2a ? _GEN_4436 : _GEN_3756; // @[executor.scala 473:84]
  wire [7:0] _GEN_4441 = _GEN_8970 == 8'h2a ? _GEN_4437 : _GEN_3757; // @[executor.scala 473:84]
  wire [7:0] _GEN_4442 = _GEN_8970 == 8'h2a ? _GEN_4438 : _GEN_3758; // @[executor.scala 473:84]
  wire [7:0] _GEN_4443 = _GEN_8970 == 8'h2a ? _GEN_4439 : _GEN_3759; // @[executor.scala 473:84]
  wire [7:0] _GEN_4444 = mask_2[0] ? byte_1024 : _GEN_3760; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4445 = mask_2[1] ? byte_1025 : _GEN_3761; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4446 = mask_2[2] ? byte_1026 : _GEN_3762; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4447 = mask_2[3] ? byte_1027 : _GEN_3763; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4448 = _GEN_8970 == 8'h2b ? _GEN_4444 : _GEN_3760; // @[executor.scala 473:84]
  wire [7:0] _GEN_4449 = _GEN_8970 == 8'h2b ? _GEN_4445 : _GEN_3761; // @[executor.scala 473:84]
  wire [7:0] _GEN_4450 = _GEN_8970 == 8'h2b ? _GEN_4446 : _GEN_3762; // @[executor.scala 473:84]
  wire [7:0] _GEN_4451 = _GEN_8970 == 8'h2b ? _GEN_4447 : _GEN_3763; // @[executor.scala 473:84]
  wire [7:0] _GEN_4452 = mask_2[0] ? byte_1024 : _GEN_3764; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4453 = mask_2[1] ? byte_1025 : _GEN_3765; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4454 = mask_2[2] ? byte_1026 : _GEN_3766; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4455 = mask_2[3] ? byte_1027 : _GEN_3767; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4456 = _GEN_8970 == 8'h2c ? _GEN_4452 : _GEN_3764; // @[executor.scala 473:84]
  wire [7:0] _GEN_4457 = _GEN_8970 == 8'h2c ? _GEN_4453 : _GEN_3765; // @[executor.scala 473:84]
  wire [7:0] _GEN_4458 = _GEN_8970 == 8'h2c ? _GEN_4454 : _GEN_3766; // @[executor.scala 473:84]
  wire [7:0] _GEN_4459 = _GEN_8970 == 8'h2c ? _GEN_4455 : _GEN_3767; // @[executor.scala 473:84]
  wire [7:0] _GEN_4460 = mask_2[0] ? byte_1024 : _GEN_3768; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4461 = mask_2[1] ? byte_1025 : _GEN_3769; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4462 = mask_2[2] ? byte_1026 : _GEN_3770; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4463 = mask_2[3] ? byte_1027 : _GEN_3771; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4464 = _GEN_8970 == 8'h2d ? _GEN_4460 : _GEN_3768; // @[executor.scala 473:84]
  wire [7:0] _GEN_4465 = _GEN_8970 == 8'h2d ? _GEN_4461 : _GEN_3769; // @[executor.scala 473:84]
  wire [7:0] _GEN_4466 = _GEN_8970 == 8'h2d ? _GEN_4462 : _GEN_3770; // @[executor.scala 473:84]
  wire [7:0] _GEN_4467 = _GEN_8970 == 8'h2d ? _GEN_4463 : _GEN_3771; // @[executor.scala 473:84]
  wire [7:0] _GEN_4468 = mask_2[0] ? byte_1024 : _GEN_3772; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4469 = mask_2[1] ? byte_1025 : _GEN_3773; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4470 = mask_2[2] ? byte_1026 : _GEN_3774; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4471 = mask_2[3] ? byte_1027 : _GEN_3775; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4472 = _GEN_8970 == 8'h2e ? _GEN_4468 : _GEN_3772; // @[executor.scala 473:84]
  wire [7:0] _GEN_4473 = _GEN_8970 == 8'h2e ? _GEN_4469 : _GEN_3773; // @[executor.scala 473:84]
  wire [7:0] _GEN_4474 = _GEN_8970 == 8'h2e ? _GEN_4470 : _GEN_3774; // @[executor.scala 473:84]
  wire [7:0] _GEN_4475 = _GEN_8970 == 8'h2e ? _GEN_4471 : _GEN_3775; // @[executor.scala 473:84]
  wire [7:0] _GEN_4476 = mask_2[0] ? byte_1024 : _GEN_3776; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4477 = mask_2[1] ? byte_1025 : _GEN_3777; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4478 = mask_2[2] ? byte_1026 : _GEN_3778; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4479 = mask_2[3] ? byte_1027 : _GEN_3779; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4480 = _GEN_8970 == 8'h2f ? _GEN_4476 : _GEN_3776; // @[executor.scala 473:84]
  wire [7:0] _GEN_4481 = _GEN_8970 == 8'h2f ? _GEN_4477 : _GEN_3777; // @[executor.scala 473:84]
  wire [7:0] _GEN_4482 = _GEN_8970 == 8'h2f ? _GEN_4478 : _GEN_3778; // @[executor.scala 473:84]
  wire [7:0] _GEN_4483 = _GEN_8970 == 8'h2f ? _GEN_4479 : _GEN_3779; // @[executor.scala 473:84]
  wire [7:0] _GEN_4484 = mask_2[0] ? byte_1024 : _GEN_3780; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4485 = mask_2[1] ? byte_1025 : _GEN_3781; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4486 = mask_2[2] ? byte_1026 : _GEN_3782; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4487 = mask_2[3] ? byte_1027 : _GEN_3783; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4488 = _GEN_8970 == 8'h30 ? _GEN_4484 : _GEN_3780; // @[executor.scala 473:84]
  wire [7:0] _GEN_4489 = _GEN_8970 == 8'h30 ? _GEN_4485 : _GEN_3781; // @[executor.scala 473:84]
  wire [7:0] _GEN_4490 = _GEN_8970 == 8'h30 ? _GEN_4486 : _GEN_3782; // @[executor.scala 473:84]
  wire [7:0] _GEN_4491 = _GEN_8970 == 8'h30 ? _GEN_4487 : _GEN_3783; // @[executor.scala 473:84]
  wire [7:0] _GEN_4492 = mask_2[0] ? byte_1024 : _GEN_3784; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4493 = mask_2[1] ? byte_1025 : _GEN_3785; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4494 = mask_2[2] ? byte_1026 : _GEN_3786; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4495 = mask_2[3] ? byte_1027 : _GEN_3787; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4496 = _GEN_8970 == 8'h31 ? _GEN_4492 : _GEN_3784; // @[executor.scala 473:84]
  wire [7:0] _GEN_4497 = _GEN_8970 == 8'h31 ? _GEN_4493 : _GEN_3785; // @[executor.scala 473:84]
  wire [7:0] _GEN_4498 = _GEN_8970 == 8'h31 ? _GEN_4494 : _GEN_3786; // @[executor.scala 473:84]
  wire [7:0] _GEN_4499 = _GEN_8970 == 8'h31 ? _GEN_4495 : _GEN_3787; // @[executor.scala 473:84]
  wire [7:0] _GEN_4500 = mask_2[0] ? byte_1024 : _GEN_3788; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4501 = mask_2[1] ? byte_1025 : _GEN_3789; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4502 = mask_2[2] ? byte_1026 : _GEN_3790; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4503 = mask_2[3] ? byte_1027 : _GEN_3791; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4504 = _GEN_8970 == 8'h32 ? _GEN_4500 : _GEN_3788; // @[executor.scala 473:84]
  wire [7:0] _GEN_4505 = _GEN_8970 == 8'h32 ? _GEN_4501 : _GEN_3789; // @[executor.scala 473:84]
  wire [7:0] _GEN_4506 = _GEN_8970 == 8'h32 ? _GEN_4502 : _GEN_3790; // @[executor.scala 473:84]
  wire [7:0] _GEN_4507 = _GEN_8970 == 8'h32 ? _GEN_4503 : _GEN_3791; // @[executor.scala 473:84]
  wire [7:0] _GEN_4508 = mask_2[0] ? byte_1024 : _GEN_3792; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4509 = mask_2[1] ? byte_1025 : _GEN_3793; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4510 = mask_2[2] ? byte_1026 : _GEN_3794; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4511 = mask_2[3] ? byte_1027 : _GEN_3795; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4512 = _GEN_8970 == 8'h33 ? _GEN_4508 : _GEN_3792; // @[executor.scala 473:84]
  wire [7:0] _GEN_4513 = _GEN_8970 == 8'h33 ? _GEN_4509 : _GEN_3793; // @[executor.scala 473:84]
  wire [7:0] _GEN_4514 = _GEN_8970 == 8'h33 ? _GEN_4510 : _GEN_3794; // @[executor.scala 473:84]
  wire [7:0] _GEN_4515 = _GEN_8970 == 8'h33 ? _GEN_4511 : _GEN_3795; // @[executor.scala 473:84]
  wire [7:0] _GEN_4516 = mask_2[0] ? byte_1024 : _GEN_3796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4517 = mask_2[1] ? byte_1025 : _GEN_3797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4518 = mask_2[2] ? byte_1026 : _GEN_3798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4519 = mask_2[3] ? byte_1027 : _GEN_3799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4520 = _GEN_8970 == 8'h34 ? _GEN_4516 : _GEN_3796; // @[executor.scala 473:84]
  wire [7:0] _GEN_4521 = _GEN_8970 == 8'h34 ? _GEN_4517 : _GEN_3797; // @[executor.scala 473:84]
  wire [7:0] _GEN_4522 = _GEN_8970 == 8'h34 ? _GEN_4518 : _GEN_3798; // @[executor.scala 473:84]
  wire [7:0] _GEN_4523 = _GEN_8970 == 8'h34 ? _GEN_4519 : _GEN_3799; // @[executor.scala 473:84]
  wire [7:0] _GEN_4524 = mask_2[0] ? byte_1024 : _GEN_3800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4525 = mask_2[1] ? byte_1025 : _GEN_3801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4526 = mask_2[2] ? byte_1026 : _GEN_3802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4527 = mask_2[3] ? byte_1027 : _GEN_3803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4528 = _GEN_8970 == 8'h35 ? _GEN_4524 : _GEN_3800; // @[executor.scala 473:84]
  wire [7:0] _GEN_4529 = _GEN_8970 == 8'h35 ? _GEN_4525 : _GEN_3801; // @[executor.scala 473:84]
  wire [7:0] _GEN_4530 = _GEN_8970 == 8'h35 ? _GEN_4526 : _GEN_3802; // @[executor.scala 473:84]
  wire [7:0] _GEN_4531 = _GEN_8970 == 8'h35 ? _GEN_4527 : _GEN_3803; // @[executor.scala 473:84]
  wire [7:0] _GEN_4532 = mask_2[0] ? byte_1024 : _GEN_3804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4533 = mask_2[1] ? byte_1025 : _GEN_3805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4534 = mask_2[2] ? byte_1026 : _GEN_3806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4535 = mask_2[3] ? byte_1027 : _GEN_3807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4536 = _GEN_8970 == 8'h36 ? _GEN_4532 : _GEN_3804; // @[executor.scala 473:84]
  wire [7:0] _GEN_4537 = _GEN_8970 == 8'h36 ? _GEN_4533 : _GEN_3805; // @[executor.scala 473:84]
  wire [7:0] _GEN_4538 = _GEN_8970 == 8'h36 ? _GEN_4534 : _GEN_3806; // @[executor.scala 473:84]
  wire [7:0] _GEN_4539 = _GEN_8970 == 8'h36 ? _GEN_4535 : _GEN_3807; // @[executor.scala 473:84]
  wire [7:0] _GEN_4540 = mask_2[0] ? byte_1024 : _GEN_3808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4541 = mask_2[1] ? byte_1025 : _GEN_3809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4542 = mask_2[2] ? byte_1026 : _GEN_3810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4543 = mask_2[3] ? byte_1027 : _GEN_3811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4544 = _GEN_8970 == 8'h37 ? _GEN_4540 : _GEN_3808; // @[executor.scala 473:84]
  wire [7:0] _GEN_4545 = _GEN_8970 == 8'h37 ? _GEN_4541 : _GEN_3809; // @[executor.scala 473:84]
  wire [7:0] _GEN_4546 = _GEN_8970 == 8'h37 ? _GEN_4542 : _GEN_3810; // @[executor.scala 473:84]
  wire [7:0] _GEN_4547 = _GEN_8970 == 8'h37 ? _GEN_4543 : _GEN_3811; // @[executor.scala 473:84]
  wire [7:0] _GEN_4548 = mask_2[0] ? byte_1024 : _GEN_3812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4549 = mask_2[1] ? byte_1025 : _GEN_3813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4550 = mask_2[2] ? byte_1026 : _GEN_3814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4551 = mask_2[3] ? byte_1027 : _GEN_3815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4552 = _GEN_8970 == 8'h38 ? _GEN_4548 : _GEN_3812; // @[executor.scala 473:84]
  wire [7:0] _GEN_4553 = _GEN_8970 == 8'h38 ? _GEN_4549 : _GEN_3813; // @[executor.scala 473:84]
  wire [7:0] _GEN_4554 = _GEN_8970 == 8'h38 ? _GEN_4550 : _GEN_3814; // @[executor.scala 473:84]
  wire [7:0] _GEN_4555 = _GEN_8970 == 8'h38 ? _GEN_4551 : _GEN_3815; // @[executor.scala 473:84]
  wire [7:0] _GEN_4556 = mask_2[0] ? byte_1024 : _GEN_3816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4557 = mask_2[1] ? byte_1025 : _GEN_3817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4558 = mask_2[2] ? byte_1026 : _GEN_3818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4559 = mask_2[3] ? byte_1027 : _GEN_3819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4560 = _GEN_8970 == 8'h39 ? _GEN_4556 : _GEN_3816; // @[executor.scala 473:84]
  wire [7:0] _GEN_4561 = _GEN_8970 == 8'h39 ? _GEN_4557 : _GEN_3817; // @[executor.scala 473:84]
  wire [7:0] _GEN_4562 = _GEN_8970 == 8'h39 ? _GEN_4558 : _GEN_3818; // @[executor.scala 473:84]
  wire [7:0] _GEN_4563 = _GEN_8970 == 8'h39 ? _GEN_4559 : _GEN_3819; // @[executor.scala 473:84]
  wire [7:0] _GEN_4564 = mask_2[0] ? byte_1024 : _GEN_3820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4565 = mask_2[1] ? byte_1025 : _GEN_3821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4566 = mask_2[2] ? byte_1026 : _GEN_3822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4567 = mask_2[3] ? byte_1027 : _GEN_3823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4568 = _GEN_8970 == 8'h3a ? _GEN_4564 : _GEN_3820; // @[executor.scala 473:84]
  wire [7:0] _GEN_4569 = _GEN_8970 == 8'h3a ? _GEN_4565 : _GEN_3821; // @[executor.scala 473:84]
  wire [7:0] _GEN_4570 = _GEN_8970 == 8'h3a ? _GEN_4566 : _GEN_3822; // @[executor.scala 473:84]
  wire [7:0] _GEN_4571 = _GEN_8970 == 8'h3a ? _GEN_4567 : _GEN_3823; // @[executor.scala 473:84]
  wire [7:0] _GEN_4572 = mask_2[0] ? byte_1024 : _GEN_3824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4573 = mask_2[1] ? byte_1025 : _GEN_3825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4574 = mask_2[2] ? byte_1026 : _GEN_3826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4575 = mask_2[3] ? byte_1027 : _GEN_3827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4576 = _GEN_8970 == 8'h3b ? _GEN_4572 : _GEN_3824; // @[executor.scala 473:84]
  wire [7:0] _GEN_4577 = _GEN_8970 == 8'h3b ? _GEN_4573 : _GEN_3825; // @[executor.scala 473:84]
  wire [7:0] _GEN_4578 = _GEN_8970 == 8'h3b ? _GEN_4574 : _GEN_3826; // @[executor.scala 473:84]
  wire [7:0] _GEN_4579 = _GEN_8970 == 8'h3b ? _GEN_4575 : _GEN_3827; // @[executor.scala 473:84]
  wire [7:0] _GEN_4580 = mask_2[0] ? byte_1024 : _GEN_3828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4581 = mask_2[1] ? byte_1025 : _GEN_3829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4582 = mask_2[2] ? byte_1026 : _GEN_3830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4583 = mask_2[3] ? byte_1027 : _GEN_3831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4584 = _GEN_8970 == 8'h3c ? _GEN_4580 : _GEN_3828; // @[executor.scala 473:84]
  wire [7:0] _GEN_4585 = _GEN_8970 == 8'h3c ? _GEN_4581 : _GEN_3829; // @[executor.scala 473:84]
  wire [7:0] _GEN_4586 = _GEN_8970 == 8'h3c ? _GEN_4582 : _GEN_3830; // @[executor.scala 473:84]
  wire [7:0] _GEN_4587 = _GEN_8970 == 8'h3c ? _GEN_4583 : _GEN_3831; // @[executor.scala 473:84]
  wire [7:0] _GEN_4588 = mask_2[0] ? byte_1024 : _GEN_3832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4589 = mask_2[1] ? byte_1025 : _GEN_3833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4590 = mask_2[2] ? byte_1026 : _GEN_3834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4591 = mask_2[3] ? byte_1027 : _GEN_3835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4592 = _GEN_8970 == 8'h3d ? _GEN_4588 : _GEN_3832; // @[executor.scala 473:84]
  wire [7:0] _GEN_4593 = _GEN_8970 == 8'h3d ? _GEN_4589 : _GEN_3833; // @[executor.scala 473:84]
  wire [7:0] _GEN_4594 = _GEN_8970 == 8'h3d ? _GEN_4590 : _GEN_3834; // @[executor.scala 473:84]
  wire [7:0] _GEN_4595 = _GEN_8970 == 8'h3d ? _GEN_4591 : _GEN_3835; // @[executor.scala 473:84]
  wire [7:0] _GEN_4596 = mask_2[0] ? byte_1024 : _GEN_3836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4597 = mask_2[1] ? byte_1025 : _GEN_3837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4598 = mask_2[2] ? byte_1026 : _GEN_3838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4599 = mask_2[3] ? byte_1027 : _GEN_3839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4600 = _GEN_8970 == 8'h3e ? _GEN_4596 : _GEN_3836; // @[executor.scala 473:84]
  wire [7:0] _GEN_4601 = _GEN_8970 == 8'h3e ? _GEN_4597 : _GEN_3837; // @[executor.scala 473:84]
  wire [7:0] _GEN_4602 = _GEN_8970 == 8'h3e ? _GEN_4598 : _GEN_3838; // @[executor.scala 473:84]
  wire [7:0] _GEN_4603 = _GEN_8970 == 8'h3e ? _GEN_4599 : _GEN_3839; // @[executor.scala 473:84]
  wire [7:0] _GEN_4604 = mask_2[0] ? byte_1024 : _GEN_3840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4605 = mask_2[1] ? byte_1025 : _GEN_3841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4606 = mask_2[2] ? byte_1026 : _GEN_3842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4607 = mask_2[3] ? byte_1027 : _GEN_3843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4608 = _GEN_8970 == 8'h3f ? _GEN_4604 : _GEN_3840; // @[executor.scala 473:84]
  wire [7:0] _GEN_4609 = _GEN_8970 == 8'h3f ? _GEN_4605 : _GEN_3841; // @[executor.scala 473:84]
  wire [7:0] _GEN_4610 = _GEN_8970 == 8'h3f ? _GEN_4606 : _GEN_3842; // @[executor.scala 473:84]
  wire [7:0] _GEN_4611 = _GEN_8970 == 8'h3f ? _GEN_4607 : _GEN_3843; // @[executor.scala 473:84]
  wire [7:0] _GEN_4612 = mask_2[0] ? byte_1024 : _GEN_3844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4613 = mask_2[1] ? byte_1025 : _GEN_3845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4614 = mask_2[2] ? byte_1026 : _GEN_3846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4615 = mask_2[3] ? byte_1027 : _GEN_3847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4616 = _GEN_8970 == 8'h40 ? _GEN_4612 : _GEN_3844; // @[executor.scala 473:84]
  wire [7:0] _GEN_4617 = _GEN_8970 == 8'h40 ? _GEN_4613 : _GEN_3845; // @[executor.scala 473:84]
  wire [7:0] _GEN_4618 = _GEN_8970 == 8'h40 ? _GEN_4614 : _GEN_3846; // @[executor.scala 473:84]
  wire [7:0] _GEN_4619 = _GEN_8970 == 8'h40 ? _GEN_4615 : _GEN_3847; // @[executor.scala 473:84]
  wire [7:0] _GEN_4620 = mask_2[0] ? byte_1024 : _GEN_3848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4621 = mask_2[1] ? byte_1025 : _GEN_3849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4622 = mask_2[2] ? byte_1026 : _GEN_3850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4623 = mask_2[3] ? byte_1027 : _GEN_3851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4624 = _GEN_8970 == 8'h41 ? _GEN_4620 : _GEN_3848; // @[executor.scala 473:84]
  wire [7:0] _GEN_4625 = _GEN_8970 == 8'h41 ? _GEN_4621 : _GEN_3849; // @[executor.scala 473:84]
  wire [7:0] _GEN_4626 = _GEN_8970 == 8'h41 ? _GEN_4622 : _GEN_3850; // @[executor.scala 473:84]
  wire [7:0] _GEN_4627 = _GEN_8970 == 8'h41 ? _GEN_4623 : _GEN_3851; // @[executor.scala 473:84]
  wire [7:0] _GEN_4628 = mask_2[0] ? byte_1024 : _GEN_3852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4629 = mask_2[1] ? byte_1025 : _GEN_3853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4630 = mask_2[2] ? byte_1026 : _GEN_3854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4631 = mask_2[3] ? byte_1027 : _GEN_3855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4632 = _GEN_8970 == 8'h42 ? _GEN_4628 : _GEN_3852; // @[executor.scala 473:84]
  wire [7:0] _GEN_4633 = _GEN_8970 == 8'h42 ? _GEN_4629 : _GEN_3853; // @[executor.scala 473:84]
  wire [7:0] _GEN_4634 = _GEN_8970 == 8'h42 ? _GEN_4630 : _GEN_3854; // @[executor.scala 473:84]
  wire [7:0] _GEN_4635 = _GEN_8970 == 8'h42 ? _GEN_4631 : _GEN_3855; // @[executor.scala 473:84]
  wire [7:0] _GEN_4636 = mask_2[0] ? byte_1024 : _GEN_3856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4637 = mask_2[1] ? byte_1025 : _GEN_3857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4638 = mask_2[2] ? byte_1026 : _GEN_3858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4639 = mask_2[3] ? byte_1027 : _GEN_3859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4640 = _GEN_8970 == 8'h43 ? _GEN_4636 : _GEN_3856; // @[executor.scala 473:84]
  wire [7:0] _GEN_4641 = _GEN_8970 == 8'h43 ? _GEN_4637 : _GEN_3857; // @[executor.scala 473:84]
  wire [7:0] _GEN_4642 = _GEN_8970 == 8'h43 ? _GEN_4638 : _GEN_3858; // @[executor.scala 473:84]
  wire [7:0] _GEN_4643 = _GEN_8970 == 8'h43 ? _GEN_4639 : _GEN_3859; // @[executor.scala 473:84]
  wire [7:0] _GEN_4644 = mask_2[0] ? byte_1024 : _GEN_3860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4645 = mask_2[1] ? byte_1025 : _GEN_3861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4646 = mask_2[2] ? byte_1026 : _GEN_3862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4647 = mask_2[3] ? byte_1027 : _GEN_3863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4648 = _GEN_8970 == 8'h44 ? _GEN_4644 : _GEN_3860; // @[executor.scala 473:84]
  wire [7:0] _GEN_4649 = _GEN_8970 == 8'h44 ? _GEN_4645 : _GEN_3861; // @[executor.scala 473:84]
  wire [7:0] _GEN_4650 = _GEN_8970 == 8'h44 ? _GEN_4646 : _GEN_3862; // @[executor.scala 473:84]
  wire [7:0] _GEN_4651 = _GEN_8970 == 8'h44 ? _GEN_4647 : _GEN_3863; // @[executor.scala 473:84]
  wire [7:0] _GEN_4652 = mask_2[0] ? byte_1024 : _GEN_3864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4653 = mask_2[1] ? byte_1025 : _GEN_3865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4654 = mask_2[2] ? byte_1026 : _GEN_3866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4655 = mask_2[3] ? byte_1027 : _GEN_3867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4656 = _GEN_8970 == 8'h45 ? _GEN_4652 : _GEN_3864; // @[executor.scala 473:84]
  wire [7:0] _GEN_4657 = _GEN_8970 == 8'h45 ? _GEN_4653 : _GEN_3865; // @[executor.scala 473:84]
  wire [7:0] _GEN_4658 = _GEN_8970 == 8'h45 ? _GEN_4654 : _GEN_3866; // @[executor.scala 473:84]
  wire [7:0] _GEN_4659 = _GEN_8970 == 8'h45 ? _GEN_4655 : _GEN_3867; // @[executor.scala 473:84]
  wire [7:0] _GEN_4660 = mask_2[0] ? byte_1024 : _GEN_3868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4661 = mask_2[1] ? byte_1025 : _GEN_3869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4662 = mask_2[2] ? byte_1026 : _GEN_3870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4663 = mask_2[3] ? byte_1027 : _GEN_3871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4664 = _GEN_8970 == 8'h46 ? _GEN_4660 : _GEN_3868; // @[executor.scala 473:84]
  wire [7:0] _GEN_4665 = _GEN_8970 == 8'h46 ? _GEN_4661 : _GEN_3869; // @[executor.scala 473:84]
  wire [7:0] _GEN_4666 = _GEN_8970 == 8'h46 ? _GEN_4662 : _GEN_3870; // @[executor.scala 473:84]
  wire [7:0] _GEN_4667 = _GEN_8970 == 8'h46 ? _GEN_4663 : _GEN_3871; // @[executor.scala 473:84]
  wire [7:0] _GEN_4668 = mask_2[0] ? byte_1024 : _GEN_3872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4669 = mask_2[1] ? byte_1025 : _GEN_3873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4670 = mask_2[2] ? byte_1026 : _GEN_3874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4671 = mask_2[3] ? byte_1027 : _GEN_3875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4672 = _GEN_8970 == 8'h47 ? _GEN_4668 : _GEN_3872; // @[executor.scala 473:84]
  wire [7:0] _GEN_4673 = _GEN_8970 == 8'h47 ? _GEN_4669 : _GEN_3873; // @[executor.scala 473:84]
  wire [7:0] _GEN_4674 = _GEN_8970 == 8'h47 ? _GEN_4670 : _GEN_3874; // @[executor.scala 473:84]
  wire [7:0] _GEN_4675 = _GEN_8970 == 8'h47 ? _GEN_4671 : _GEN_3875; // @[executor.scala 473:84]
  wire [7:0] _GEN_4676 = mask_2[0] ? byte_1024 : _GEN_3876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4677 = mask_2[1] ? byte_1025 : _GEN_3877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4678 = mask_2[2] ? byte_1026 : _GEN_3878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4679 = mask_2[3] ? byte_1027 : _GEN_3879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4680 = _GEN_8970 == 8'h48 ? _GEN_4676 : _GEN_3876; // @[executor.scala 473:84]
  wire [7:0] _GEN_4681 = _GEN_8970 == 8'h48 ? _GEN_4677 : _GEN_3877; // @[executor.scala 473:84]
  wire [7:0] _GEN_4682 = _GEN_8970 == 8'h48 ? _GEN_4678 : _GEN_3878; // @[executor.scala 473:84]
  wire [7:0] _GEN_4683 = _GEN_8970 == 8'h48 ? _GEN_4679 : _GEN_3879; // @[executor.scala 473:84]
  wire [7:0] _GEN_4684 = mask_2[0] ? byte_1024 : _GEN_3880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4685 = mask_2[1] ? byte_1025 : _GEN_3881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4686 = mask_2[2] ? byte_1026 : _GEN_3882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4687 = mask_2[3] ? byte_1027 : _GEN_3883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4688 = _GEN_8970 == 8'h49 ? _GEN_4684 : _GEN_3880; // @[executor.scala 473:84]
  wire [7:0] _GEN_4689 = _GEN_8970 == 8'h49 ? _GEN_4685 : _GEN_3881; // @[executor.scala 473:84]
  wire [7:0] _GEN_4690 = _GEN_8970 == 8'h49 ? _GEN_4686 : _GEN_3882; // @[executor.scala 473:84]
  wire [7:0] _GEN_4691 = _GEN_8970 == 8'h49 ? _GEN_4687 : _GEN_3883; // @[executor.scala 473:84]
  wire [7:0] _GEN_4692 = mask_2[0] ? byte_1024 : _GEN_3884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4693 = mask_2[1] ? byte_1025 : _GEN_3885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4694 = mask_2[2] ? byte_1026 : _GEN_3886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4695 = mask_2[3] ? byte_1027 : _GEN_3887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4696 = _GEN_8970 == 8'h4a ? _GEN_4692 : _GEN_3884; // @[executor.scala 473:84]
  wire [7:0] _GEN_4697 = _GEN_8970 == 8'h4a ? _GEN_4693 : _GEN_3885; // @[executor.scala 473:84]
  wire [7:0] _GEN_4698 = _GEN_8970 == 8'h4a ? _GEN_4694 : _GEN_3886; // @[executor.scala 473:84]
  wire [7:0] _GEN_4699 = _GEN_8970 == 8'h4a ? _GEN_4695 : _GEN_3887; // @[executor.scala 473:84]
  wire [7:0] _GEN_4700 = mask_2[0] ? byte_1024 : _GEN_3888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4701 = mask_2[1] ? byte_1025 : _GEN_3889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4702 = mask_2[2] ? byte_1026 : _GEN_3890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4703 = mask_2[3] ? byte_1027 : _GEN_3891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4704 = _GEN_8970 == 8'h4b ? _GEN_4700 : _GEN_3888; // @[executor.scala 473:84]
  wire [7:0] _GEN_4705 = _GEN_8970 == 8'h4b ? _GEN_4701 : _GEN_3889; // @[executor.scala 473:84]
  wire [7:0] _GEN_4706 = _GEN_8970 == 8'h4b ? _GEN_4702 : _GEN_3890; // @[executor.scala 473:84]
  wire [7:0] _GEN_4707 = _GEN_8970 == 8'h4b ? _GEN_4703 : _GEN_3891; // @[executor.scala 473:84]
  wire [7:0] _GEN_4708 = mask_2[0] ? byte_1024 : _GEN_3892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4709 = mask_2[1] ? byte_1025 : _GEN_3893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4710 = mask_2[2] ? byte_1026 : _GEN_3894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4711 = mask_2[3] ? byte_1027 : _GEN_3895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4712 = _GEN_8970 == 8'h4c ? _GEN_4708 : _GEN_3892; // @[executor.scala 473:84]
  wire [7:0] _GEN_4713 = _GEN_8970 == 8'h4c ? _GEN_4709 : _GEN_3893; // @[executor.scala 473:84]
  wire [7:0] _GEN_4714 = _GEN_8970 == 8'h4c ? _GEN_4710 : _GEN_3894; // @[executor.scala 473:84]
  wire [7:0] _GEN_4715 = _GEN_8970 == 8'h4c ? _GEN_4711 : _GEN_3895; // @[executor.scala 473:84]
  wire [7:0] _GEN_4716 = mask_2[0] ? byte_1024 : _GEN_3896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4717 = mask_2[1] ? byte_1025 : _GEN_3897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4718 = mask_2[2] ? byte_1026 : _GEN_3898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4719 = mask_2[3] ? byte_1027 : _GEN_3899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4720 = _GEN_8970 == 8'h4d ? _GEN_4716 : _GEN_3896; // @[executor.scala 473:84]
  wire [7:0] _GEN_4721 = _GEN_8970 == 8'h4d ? _GEN_4717 : _GEN_3897; // @[executor.scala 473:84]
  wire [7:0] _GEN_4722 = _GEN_8970 == 8'h4d ? _GEN_4718 : _GEN_3898; // @[executor.scala 473:84]
  wire [7:0] _GEN_4723 = _GEN_8970 == 8'h4d ? _GEN_4719 : _GEN_3899; // @[executor.scala 473:84]
  wire [7:0] _GEN_4724 = mask_2[0] ? byte_1024 : _GEN_3900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4725 = mask_2[1] ? byte_1025 : _GEN_3901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4726 = mask_2[2] ? byte_1026 : _GEN_3902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4727 = mask_2[3] ? byte_1027 : _GEN_3903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4728 = _GEN_8970 == 8'h4e ? _GEN_4724 : _GEN_3900; // @[executor.scala 473:84]
  wire [7:0] _GEN_4729 = _GEN_8970 == 8'h4e ? _GEN_4725 : _GEN_3901; // @[executor.scala 473:84]
  wire [7:0] _GEN_4730 = _GEN_8970 == 8'h4e ? _GEN_4726 : _GEN_3902; // @[executor.scala 473:84]
  wire [7:0] _GEN_4731 = _GEN_8970 == 8'h4e ? _GEN_4727 : _GEN_3903; // @[executor.scala 473:84]
  wire [7:0] _GEN_4732 = mask_2[0] ? byte_1024 : _GEN_3904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4733 = mask_2[1] ? byte_1025 : _GEN_3905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4734 = mask_2[2] ? byte_1026 : _GEN_3906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4735 = mask_2[3] ? byte_1027 : _GEN_3907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4736 = _GEN_8970 == 8'h4f ? _GEN_4732 : _GEN_3904; // @[executor.scala 473:84]
  wire [7:0] _GEN_4737 = _GEN_8970 == 8'h4f ? _GEN_4733 : _GEN_3905; // @[executor.scala 473:84]
  wire [7:0] _GEN_4738 = _GEN_8970 == 8'h4f ? _GEN_4734 : _GEN_3906; // @[executor.scala 473:84]
  wire [7:0] _GEN_4739 = _GEN_8970 == 8'h4f ? _GEN_4735 : _GEN_3907; // @[executor.scala 473:84]
  wire [7:0] _GEN_4740 = mask_2[0] ? byte_1024 : _GEN_3908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4741 = mask_2[1] ? byte_1025 : _GEN_3909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4742 = mask_2[2] ? byte_1026 : _GEN_3910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4743 = mask_2[3] ? byte_1027 : _GEN_3911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4744 = _GEN_8970 == 8'h50 ? _GEN_4740 : _GEN_3908; // @[executor.scala 473:84]
  wire [7:0] _GEN_4745 = _GEN_8970 == 8'h50 ? _GEN_4741 : _GEN_3909; // @[executor.scala 473:84]
  wire [7:0] _GEN_4746 = _GEN_8970 == 8'h50 ? _GEN_4742 : _GEN_3910; // @[executor.scala 473:84]
  wire [7:0] _GEN_4747 = _GEN_8970 == 8'h50 ? _GEN_4743 : _GEN_3911; // @[executor.scala 473:84]
  wire [7:0] _GEN_4748 = mask_2[0] ? byte_1024 : _GEN_3912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4749 = mask_2[1] ? byte_1025 : _GEN_3913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4750 = mask_2[2] ? byte_1026 : _GEN_3914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4751 = mask_2[3] ? byte_1027 : _GEN_3915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4752 = _GEN_8970 == 8'h51 ? _GEN_4748 : _GEN_3912; // @[executor.scala 473:84]
  wire [7:0] _GEN_4753 = _GEN_8970 == 8'h51 ? _GEN_4749 : _GEN_3913; // @[executor.scala 473:84]
  wire [7:0] _GEN_4754 = _GEN_8970 == 8'h51 ? _GEN_4750 : _GEN_3914; // @[executor.scala 473:84]
  wire [7:0] _GEN_4755 = _GEN_8970 == 8'h51 ? _GEN_4751 : _GEN_3915; // @[executor.scala 473:84]
  wire [7:0] _GEN_4756 = mask_2[0] ? byte_1024 : _GEN_3916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4757 = mask_2[1] ? byte_1025 : _GEN_3917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4758 = mask_2[2] ? byte_1026 : _GEN_3918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4759 = mask_2[3] ? byte_1027 : _GEN_3919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4760 = _GEN_8970 == 8'h52 ? _GEN_4756 : _GEN_3916; // @[executor.scala 473:84]
  wire [7:0] _GEN_4761 = _GEN_8970 == 8'h52 ? _GEN_4757 : _GEN_3917; // @[executor.scala 473:84]
  wire [7:0] _GEN_4762 = _GEN_8970 == 8'h52 ? _GEN_4758 : _GEN_3918; // @[executor.scala 473:84]
  wire [7:0] _GEN_4763 = _GEN_8970 == 8'h52 ? _GEN_4759 : _GEN_3919; // @[executor.scala 473:84]
  wire [7:0] _GEN_4764 = mask_2[0] ? byte_1024 : _GEN_3920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4765 = mask_2[1] ? byte_1025 : _GEN_3921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4766 = mask_2[2] ? byte_1026 : _GEN_3922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4767 = mask_2[3] ? byte_1027 : _GEN_3923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4768 = _GEN_8970 == 8'h53 ? _GEN_4764 : _GEN_3920; // @[executor.scala 473:84]
  wire [7:0] _GEN_4769 = _GEN_8970 == 8'h53 ? _GEN_4765 : _GEN_3921; // @[executor.scala 473:84]
  wire [7:0] _GEN_4770 = _GEN_8970 == 8'h53 ? _GEN_4766 : _GEN_3922; // @[executor.scala 473:84]
  wire [7:0] _GEN_4771 = _GEN_8970 == 8'h53 ? _GEN_4767 : _GEN_3923; // @[executor.scala 473:84]
  wire [7:0] _GEN_4772 = mask_2[0] ? byte_1024 : _GEN_3924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4773 = mask_2[1] ? byte_1025 : _GEN_3925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4774 = mask_2[2] ? byte_1026 : _GEN_3926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4775 = mask_2[3] ? byte_1027 : _GEN_3927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4776 = _GEN_8970 == 8'h54 ? _GEN_4772 : _GEN_3924; // @[executor.scala 473:84]
  wire [7:0] _GEN_4777 = _GEN_8970 == 8'h54 ? _GEN_4773 : _GEN_3925; // @[executor.scala 473:84]
  wire [7:0] _GEN_4778 = _GEN_8970 == 8'h54 ? _GEN_4774 : _GEN_3926; // @[executor.scala 473:84]
  wire [7:0] _GEN_4779 = _GEN_8970 == 8'h54 ? _GEN_4775 : _GEN_3927; // @[executor.scala 473:84]
  wire [7:0] _GEN_4780 = mask_2[0] ? byte_1024 : _GEN_3928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4781 = mask_2[1] ? byte_1025 : _GEN_3929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4782 = mask_2[2] ? byte_1026 : _GEN_3930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4783 = mask_2[3] ? byte_1027 : _GEN_3931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4784 = _GEN_8970 == 8'h55 ? _GEN_4780 : _GEN_3928; // @[executor.scala 473:84]
  wire [7:0] _GEN_4785 = _GEN_8970 == 8'h55 ? _GEN_4781 : _GEN_3929; // @[executor.scala 473:84]
  wire [7:0] _GEN_4786 = _GEN_8970 == 8'h55 ? _GEN_4782 : _GEN_3930; // @[executor.scala 473:84]
  wire [7:0] _GEN_4787 = _GEN_8970 == 8'h55 ? _GEN_4783 : _GEN_3931; // @[executor.scala 473:84]
  wire [7:0] _GEN_4788 = mask_2[0] ? byte_1024 : _GEN_3932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4789 = mask_2[1] ? byte_1025 : _GEN_3933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4790 = mask_2[2] ? byte_1026 : _GEN_3934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4791 = mask_2[3] ? byte_1027 : _GEN_3935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4792 = _GEN_8970 == 8'h56 ? _GEN_4788 : _GEN_3932; // @[executor.scala 473:84]
  wire [7:0] _GEN_4793 = _GEN_8970 == 8'h56 ? _GEN_4789 : _GEN_3933; // @[executor.scala 473:84]
  wire [7:0] _GEN_4794 = _GEN_8970 == 8'h56 ? _GEN_4790 : _GEN_3934; // @[executor.scala 473:84]
  wire [7:0] _GEN_4795 = _GEN_8970 == 8'h56 ? _GEN_4791 : _GEN_3935; // @[executor.scala 473:84]
  wire [7:0] _GEN_4796 = mask_2[0] ? byte_1024 : _GEN_3936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4797 = mask_2[1] ? byte_1025 : _GEN_3937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4798 = mask_2[2] ? byte_1026 : _GEN_3938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4799 = mask_2[3] ? byte_1027 : _GEN_3939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4800 = _GEN_8970 == 8'h57 ? _GEN_4796 : _GEN_3936; // @[executor.scala 473:84]
  wire [7:0] _GEN_4801 = _GEN_8970 == 8'h57 ? _GEN_4797 : _GEN_3937; // @[executor.scala 473:84]
  wire [7:0] _GEN_4802 = _GEN_8970 == 8'h57 ? _GEN_4798 : _GEN_3938; // @[executor.scala 473:84]
  wire [7:0] _GEN_4803 = _GEN_8970 == 8'h57 ? _GEN_4799 : _GEN_3939; // @[executor.scala 473:84]
  wire [7:0] _GEN_4804 = mask_2[0] ? byte_1024 : _GEN_3940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4805 = mask_2[1] ? byte_1025 : _GEN_3941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4806 = mask_2[2] ? byte_1026 : _GEN_3942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4807 = mask_2[3] ? byte_1027 : _GEN_3943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4808 = _GEN_8970 == 8'h58 ? _GEN_4804 : _GEN_3940; // @[executor.scala 473:84]
  wire [7:0] _GEN_4809 = _GEN_8970 == 8'h58 ? _GEN_4805 : _GEN_3941; // @[executor.scala 473:84]
  wire [7:0] _GEN_4810 = _GEN_8970 == 8'h58 ? _GEN_4806 : _GEN_3942; // @[executor.scala 473:84]
  wire [7:0] _GEN_4811 = _GEN_8970 == 8'h58 ? _GEN_4807 : _GEN_3943; // @[executor.scala 473:84]
  wire [7:0] _GEN_4812 = mask_2[0] ? byte_1024 : _GEN_3944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4813 = mask_2[1] ? byte_1025 : _GEN_3945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4814 = mask_2[2] ? byte_1026 : _GEN_3946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4815 = mask_2[3] ? byte_1027 : _GEN_3947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4816 = _GEN_8970 == 8'h59 ? _GEN_4812 : _GEN_3944; // @[executor.scala 473:84]
  wire [7:0] _GEN_4817 = _GEN_8970 == 8'h59 ? _GEN_4813 : _GEN_3945; // @[executor.scala 473:84]
  wire [7:0] _GEN_4818 = _GEN_8970 == 8'h59 ? _GEN_4814 : _GEN_3946; // @[executor.scala 473:84]
  wire [7:0] _GEN_4819 = _GEN_8970 == 8'h59 ? _GEN_4815 : _GEN_3947; // @[executor.scala 473:84]
  wire [7:0] _GEN_4820 = mask_2[0] ? byte_1024 : _GEN_3948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4821 = mask_2[1] ? byte_1025 : _GEN_3949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4822 = mask_2[2] ? byte_1026 : _GEN_3950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4823 = mask_2[3] ? byte_1027 : _GEN_3951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4824 = _GEN_8970 == 8'h5a ? _GEN_4820 : _GEN_3948; // @[executor.scala 473:84]
  wire [7:0] _GEN_4825 = _GEN_8970 == 8'h5a ? _GEN_4821 : _GEN_3949; // @[executor.scala 473:84]
  wire [7:0] _GEN_4826 = _GEN_8970 == 8'h5a ? _GEN_4822 : _GEN_3950; // @[executor.scala 473:84]
  wire [7:0] _GEN_4827 = _GEN_8970 == 8'h5a ? _GEN_4823 : _GEN_3951; // @[executor.scala 473:84]
  wire [7:0] _GEN_4828 = mask_2[0] ? byte_1024 : _GEN_3952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4829 = mask_2[1] ? byte_1025 : _GEN_3953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4830 = mask_2[2] ? byte_1026 : _GEN_3954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4831 = mask_2[3] ? byte_1027 : _GEN_3955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4832 = _GEN_8970 == 8'h5b ? _GEN_4828 : _GEN_3952; // @[executor.scala 473:84]
  wire [7:0] _GEN_4833 = _GEN_8970 == 8'h5b ? _GEN_4829 : _GEN_3953; // @[executor.scala 473:84]
  wire [7:0] _GEN_4834 = _GEN_8970 == 8'h5b ? _GEN_4830 : _GEN_3954; // @[executor.scala 473:84]
  wire [7:0] _GEN_4835 = _GEN_8970 == 8'h5b ? _GEN_4831 : _GEN_3955; // @[executor.scala 473:84]
  wire [7:0] _GEN_4836 = mask_2[0] ? byte_1024 : _GEN_3956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4837 = mask_2[1] ? byte_1025 : _GEN_3957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4838 = mask_2[2] ? byte_1026 : _GEN_3958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4839 = mask_2[3] ? byte_1027 : _GEN_3959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4840 = _GEN_8970 == 8'h5c ? _GEN_4836 : _GEN_3956; // @[executor.scala 473:84]
  wire [7:0] _GEN_4841 = _GEN_8970 == 8'h5c ? _GEN_4837 : _GEN_3957; // @[executor.scala 473:84]
  wire [7:0] _GEN_4842 = _GEN_8970 == 8'h5c ? _GEN_4838 : _GEN_3958; // @[executor.scala 473:84]
  wire [7:0] _GEN_4843 = _GEN_8970 == 8'h5c ? _GEN_4839 : _GEN_3959; // @[executor.scala 473:84]
  wire [7:0] _GEN_4844 = mask_2[0] ? byte_1024 : _GEN_3960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4845 = mask_2[1] ? byte_1025 : _GEN_3961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4846 = mask_2[2] ? byte_1026 : _GEN_3962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4847 = mask_2[3] ? byte_1027 : _GEN_3963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4848 = _GEN_8970 == 8'h5d ? _GEN_4844 : _GEN_3960; // @[executor.scala 473:84]
  wire [7:0] _GEN_4849 = _GEN_8970 == 8'h5d ? _GEN_4845 : _GEN_3961; // @[executor.scala 473:84]
  wire [7:0] _GEN_4850 = _GEN_8970 == 8'h5d ? _GEN_4846 : _GEN_3962; // @[executor.scala 473:84]
  wire [7:0] _GEN_4851 = _GEN_8970 == 8'h5d ? _GEN_4847 : _GEN_3963; // @[executor.scala 473:84]
  wire [7:0] _GEN_4852 = mask_2[0] ? byte_1024 : _GEN_3964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4853 = mask_2[1] ? byte_1025 : _GEN_3965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4854 = mask_2[2] ? byte_1026 : _GEN_3966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4855 = mask_2[3] ? byte_1027 : _GEN_3967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4856 = _GEN_8970 == 8'h5e ? _GEN_4852 : _GEN_3964; // @[executor.scala 473:84]
  wire [7:0] _GEN_4857 = _GEN_8970 == 8'h5e ? _GEN_4853 : _GEN_3965; // @[executor.scala 473:84]
  wire [7:0] _GEN_4858 = _GEN_8970 == 8'h5e ? _GEN_4854 : _GEN_3966; // @[executor.scala 473:84]
  wire [7:0] _GEN_4859 = _GEN_8970 == 8'h5e ? _GEN_4855 : _GEN_3967; // @[executor.scala 473:84]
  wire [7:0] _GEN_4860 = mask_2[0] ? byte_1024 : _GEN_3968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4861 = mask_2[1] ? byte_1025 : _GEN_3969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4862 = mask_2[2] ? byte_1026 : _GEN_3970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4863 = mask_2[3] ? byte_1027 : _GEN_3971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4864 = _GEN_8970 == 8'h5f ? _GEN_4860 : _GEN_3968; // @[executor.scala 473:84]
  wire [7:0] _GEN_4865 = _GEN_8970 == 8'h5f ? _GEN_4861 : _GEN_3969; // @[executor.scala 473:84]
  wire [7:0] _GEN_4866 = _GEN_8970 == 8'h5f ? _GEN_4862 : _GEN_3970; // @[executor.scala 473:84]
  wire [7:0] _GEN_4867 = _GEN_8970 == 8'h5f ? _GEN_4863 : _GEN_3971; // @[executor.scala 473:84]
  wire [7:0] _GEN_4868 = mask_2[0] ? byte_1024 : _GEN_3972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4869 = mask_2[1] ? byte_1025 : _GEN_3973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4870 = mask_2[2] ? byte_1026 : _GEN_3974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4871 = mask_2[3] ? byte_1027 : _GEN_3975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4872 = _GEN_8970 == 8'h60 ? _GEN_4868 : _GEN_3972; // @[executor.scala 473:84]
  wire [7:0] _GEN_4873 = _GEN_8970 == 8'h60 ? _GEN_4869 : _GEN_3973; // @[executor.scala 473:84]
  wire [7:0] _GEN_4874 = _GEN_8970 == 8'h60 ? _GEN_4870 : _GEN_3974; // @[executor.scala 473:84]
  wire [7:0] _GEN_4875 = _GEN_8970 == 8'h60 ? _GEN_4871 : _GEN_3975; // @[executor.scala 473:84]
  wire [7:0] _GEN_4876 = mask_2[0] ? byte_1024 : _GEN_3976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4877 = mask_2[1] ? byte_1025 : _GEN_3977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4878 = mask_2[2] ? byte_1026 : _GEN_3978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4879 = mask_2[3] ? byte_1027 : _GEN_3979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4880 = _GEN_8970 == 8'h61 ? _GEN_4876 : _GEN_3976; // @[executor.scala 473:84]
  wire [7:0] _GEN_4881 = _GEN_8970 == 8'h61 ? _GEN_4877 : _GEN_3977; // @[executor.scala 473:84]
  wire [7:0] _GEN_4882 = _GEN_8970 == 8'h61 ? _GEN_4878 : _GEN_3978; // @[executor.scala 473:84]
  wire [7:0] _GEN_4883 = _GEN_8970 == 8'h61 ? _GEN_4879 : _GEN_3979; // @[executor.scala 473:84]
  wire [7:0] _GEN_4884 = mask_2[0] ? byte_1024 : _GEN_3980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4885 = mask_2[1] ? byte_1025 : _GEN_3981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4886 = mask_2[2] ? byte_1026 : _GEN_3982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4887 = mask_2[3] ? byte_1027 : _GEN_3983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4888 = _GEN_8970 == 8'h62 ? _GEN_4884 : _GEN_3980; // @[executor.scala 473:84]
  wire [7:0] _GEN_4889 = _GEN_8970 == 8'h62 ? _GEN_4885 : _GEN_3981; // @[executor.scala 473:84]
  wire [7:0] _GEN_4890 = _GEN_8970 == 8'h62 ? _GEN_4886 : _GEN_3982; // @[executor.scala 473:84]
  wire [7:0] _GEN_4891 = _GEN_8970 == 8'h62 ? _GEN_4887 : _GEN_3983; // @[executor.scala 473:84]
  wire [7:0] _GEN_4892 = mask_2[0] ? byte_1024 : _GEN_3984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4893 = mask_2[1] ? byte_1025 : _GEN_3985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4894 = mask_2[2] ? byte_1026 : _GEN_3986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4895 = mask_2[3] ? byte_1027 : _GEN_3987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4896 = _GEN_8970 == 8'h63 ? _GEN_4892 : _GEN_3984; // @[executor.scala 473:84]
  wire [7:0] _GEN_4897 = _GEN_8970 == 8'h63 ? _GEN_4893 : _GEN_3985; // @[executor.scala 473:84]
  wire [7:0] _GEN_4898 = _GEN_8970 == 8'h63 ? _GEN_4894 : _GEN_3986; // @[executor.scala 473:84]
  wire [7:0] _GEN_4899 = _GEN_8970 == 8'h63 ? _GEN_4895 : _GEN_3987; // @[executor.scala 473:84]
  wire [7:0] _GEN_4900 = mask_2[0] ? byte_1024 : _GEN_3988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4901 = mask_2[1] ? byte_1025 : _GEN_3989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4902 = mask_2[2] ? byte_1026 : _GEN_3990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4903 = mask_2[3] ? byte_1027 : _GEN_3991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4904 = _GEN_8970 == 8'h64 ? _GEN_4900 : _GEN_3988; // @[executor.scala 473:84]
  wire [7:0] _GEN_4905 = _GEN_8970 == 8'h64 ? _GEN_4901 : _GEN_3989; // @[executor.scala 473:84]
  wire [7:0] _GEN_4906 = _GEN_8970 == 8'h64 ? _GEN_4902 : _GEN_3990; // @[executor.scala 473:84]
  wire [7:0] _GEN_4907 = _GEN_8970 == 8'h64 ? _GEN_4903 : _GEN_3991; // @[executor.scala 473:84]
  wire [7:0] _GEN_4908 = mask_2[0] ? byte_1024 : _GEN_3992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4909 = mask_2[1] ? byte_1025 : _GEN_3993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4910 = mask_2[2] ? byte_1026 : _GEN_3994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4911 = mask_2[3] ? byte_1027 : _GEN_3995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4912 = _GEN_8970 == 8'h65 ? _GEN_4908 : _GEN_3992; // @[executor.scala 473:84]
  wire [7:0] _GEN_4913 = _GEN_8970 == 8'h65 ? _GEN_4909 : _GEN_3993; // @[executor.scala 473:84]
  wire [7:0] _GEN_4914 = _GEN_8970 == 8'h65 ? _GEN_4910 : _GEN_3994; // @[executor.scala 473:84]
  wire [7:0] _GEN_4915 = _GEN_8970 == 8'h65 ? _GEN_4911 : _GEN_3995; // @[executor.scala 473:84]
  wire [7:0] _GEN_4916 = mask_2[0] ? byte_1024 : _GEN_3996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4917 = mask_2[1] ? byte_1025 : _GEN_3997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4918 = mask_2[2] ? byte_1026 : _GEN_3998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4919 = mask_2[3] ? byte_1027 : _GEN_3999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4920 = _GEN_8970 == 8'h66 ? _GEN_4916 : _GEN_3996; // @[executor.scala 473:84]
  wire [7:0] _GEN_4921 = _GEN_8970 == 8'h66 ? _GEN_4917 : _GEN_3997; // @[executor.scala 473:84]
  wire [7:0] _GEN_4922 = _GEN_8970 == 8'h66 ? _GEN_4918 : _GEN_3998; // @[executor.scala 473:84]
  wire [7:0] _GEN_4923 = _GEN_8970 == 8'h66 ? _GEN_4919 : _GEN_3999; // @[executor.scala 473:84]
  wire [7:0] _GEN_4924 = mask_2[0] ? byte_1024 : _GEN_4000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4925 = mask_2[1] ? byte_1025 : _GEN_4001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4926 = mask_2[2] ? byte_1026 : _GEN_4002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4927 = mask_2[3] ? byte_1027 : _GEN_4003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4928 = _GEN_8970 == 8'h67 ? _GEN_4924 : _GEN_4000; // @[executor.scala 473:84]
  wire [7:0] _GEN_4929 = _GEN_8970 == 8'h67 ? _GEN_4925 : _GEN_4001; // @[executor.scala 473:84]
  wire [7:0] _GEN_4930 = _GEN_8970 == 8'h67 ? _GEN_4926 : _GEN_4002; // @[executor.scala 473:84]
  wire [7:0] _GEN_4931 = _GEN_8970 == 8'h67 ? _GEN_4927 : _GEN_4003; // @[executor.scala 473:84]
  wire [7:0] _GEN_4932 = mask_2[0] ? byte_1024 : _GEN_4004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4933 = mask_2[1] ? byte_1025 : _GEN_4005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4934 = mask_2[2] ? byte_1026 : _GEN_4006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4935 = mask_2[3] ? byte_1027 : _GEN_4007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4936 = _GEN_8970 == 8'h68 ? _GEN_4932 : _GEN_4004; // @[executor.scala 473:84]
  wire [7:0] _GEN_4937 = _GEN_8970 == 8'h68 ? _GEN_4933 : _GEN_4005; // @[executor.scala 473:84]
  wire [7:0] _GEN_4938 = _GEN_8970 == 8'h68 ? _GEN_4934 : _GEN_4006; // @[executor.scala 473:84]
  wire [7:0] _GEN_4939 = _GEN_8970 == 8'h68 ? _GEN_4935 : _GEN_4007; // @[executor.scala 473:84]
  wire [7:0] _GEN_4940 = mask_2[0] ? byte_1024 : _GEN_4008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4941 = mask_2[1] ? byte_1025 : _GEN_4009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4942 = mask_2[2] ? byte_1026 : _GEN_4010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4943 = mask_2[3] ? byte_1027 : _GEN_4011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4944 = _GEN_8970 == 8'h69 ? _GEN_4940 : _GEN_4008; // @[executor.scala 473:84]
  wire [7:0] _GEN_4945 = _GEN_8970 == 8'h69 ? _GEN_4941 : _GEN_4009; // @[executor.scala 473:84]
  wire [7:0] _GEN_4946 = _GEN_8970 == 8'h69 ? _GEN_4942 : _GEN_4010; // @[executor.scala 473:84]
  wire [7:0] _GEN_4947 = _GEN_8970 == 8'h69 ? _GEN_4943 : _GEN_4011; // @[executor.scala 473:84]
  wire [7:0] _GEN_4948 = mask_2[0] ? byte_1024 : _GEN_4012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4949 = mask_2[1] ? byte_1025 : _GEN_4013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4950 = mask_2[2] ? byte_1026 : _GEN_4014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4951 = mask_2[3] ? byte_1027 : _GEN_4015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4952 = _GEN_8970 == 8'h6a ? _GEN_4948 : _GEN_4012; // @[executor.scala 473:84]
  wire [7:0] _GEN_4953 = _GEN_8970 == 8'h6a ? _GEN_4949 : _GEN_4013; // @[executor.scala 473:84]
  wire [7:0] _GEN_4954 = _GEN_8970 == 8'h6a ? _GEN_4950 : _GEN_4014; // @[executor.scala 473:84]
  wire [7:0] _GEN_4955 = _GEN_8970 == 8'h6a ? _GEN_4951 : _GEN_4015; // @[executor.scala 473:84]
  wire [7:0] _GEN_4956 = mask_2[0] ? byte_1024 : _GEN_4016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4957 = mask_2[1] ? byte_1025 : _GEN_4017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4958 = mask_2[2] ? byte_1026 : _GEN_4018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4959 = mask_2[3] ? byte_1027 : _GEN_4019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4960 = _GEN_8970 == 8'h6b ? _GEN_4956 : _GEN_4016; // @[executor.scala 473:84]
  wire [7:0] _GEN_4961 = _GEN_8970 == 8'h6b ? _GEN_4957 : _GEN_4017; // @[executor.scala 473:84]
  wire [7:0] _GEN_4962 = _GEN_8970 == 8'h6b ? _GEN_4958 : _GEN_4018; // @[executor.scala 473:84]
  wire [7:0] _GEN_4963 = _GEN_8970 == 8'h6b ? _GEN_4959 : _GEN_4019; // @[executor.scala 473:84]
  wire [7:0] _GEN_4964 = mask_2[0] ? byte_1024 : _GEN_4020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4965 = mask_2[1] ? byte_1025 : _GEN_4021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4966 = mask_2[2] ? byte_1026 : _GEN_4022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4967 = mask_2[3] ? byte_1027 : _GEN_4023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4968 = _GEN_8970 == 8'h6c ? _GEN_4964 : _GEN_4020; // @[executor.scala 473:84]
  wire [7:0] _GEN_4969 = _GEN_8970 == 8'h6c ? _GEN_4965 : _GEN_4021; // @[executor.scala 473:84]
  wire [7:0] _GEN_4970 = _GEN_8970 == 8'h6c ? _GEN_4966 : _GEN_4022; // @[executor.scala 473:84]
  wire [7:0] _GEN_4971 = _GEN_8970 == 8'h6c ? _GEN_4967 : _GEN_4023; // @[executor.scala 473:84]
  wire [7:0] _GEN_4972 = mask_2[0] ? byte_1024 : _GEN_4024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4973 = mask_2[1] ? byte_1025 : _GEN_4025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4974 = mask_2[2] ? byte_1026 : _GEN_4026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4975 = mask_2[3] ? byte_1027 : _GEN_4027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4976 = _GEN_8970 == 8'h6d ? _GEN_4972 : _GEN_4024; // @[executor.scala 473:84]
  wire [7:0] _GEN_4977 = _GEN_8970 == 8'h6d ? _GEN_4973 : _GEN_4025; // @[executor.scala 473:84]
  wire [7:0] _GEN_4978 = _GEN_8970 == 8'h6d ? _GEN_4974 : _GEN_4026; // @[executor.scala 473:84]
  wire [7:0] _GEN_4979 = _GEN_8970 == 8'h6d ? _GEN_4975 : _GEN_4027; // @[executor.scala 473:84]
  wire [7:0] _GEN_4980 = mask_2[0] ? byte_1024 : _GEN_4028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4981 = mask_2[1] ? byte_1025 : _GEN_4029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4982 = mask_2[2] ? byte_1026 : _GEN_4030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4983 = mask_2[3] ? byte_1027 : _GEN_4031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4984 = _GEN_8970 == 8'h6e ? _GEN_4980 : _GEN_4028; // @[executor.scala 473:84]
  wire [7:0] _GEN_4985 = _GEN_8970 == 8'h6e ? _GEN_4981 : _GEN_4029; // @[executor.scala 473:84]
  wire [7:0] _GEN_4986 = _GEN_8970 == 8'h6e ? _GEN_4982 : _GEN_4030; // @[executor.scala 473:84]
  wire [7:0] _GEN_4987 = _GEN_8970 == 8'h6e ? _GEN_4983 : _GEN_4031; // @[executor.scala 473:84]
  wire [7:0] _GEN_4988 = mask_2[0] ? byte_1024 : _GEN_4032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4989 = mask_2[1] ? byte_1025 : _GEN_4033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4990 = mask_2[2] ? byte_1026 : _GEN_4034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4991 = mask_2[3] ? byte_1027 : _GEN_4035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4992 = _GEN_8970 == 8'h6f ? _GEN_4988 : _GEN_4032; // @[executor.scala 473:84]
  wire [7:0] _GEN_4993 = _GEN_8970 == 8'h6f ? _GEN_4989 : _GEN_4033; // @[executor.scala 473:84]
  wire [7:0] _GEN_4994 = _GEN_8970 == 8'h6f ? _GEN_4990 : _GEN_4034; // @[executor.scala 473:84]
  wire [7:0] _GEN_4995 = _GEN_8970 == 8'h6f ? _GEN_4991 : _GEN_4035; // @[executor.scala 473:84]
  wire [7:0] _GEN_4996 = mask_2[0] ? byte_1024 : _GEN_4036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4997 = mask_2[1] ? byte_1025 : _GEN_4037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4998 = mask_2[2] ? byte_1026 : _GEN_4038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_4999 = mask_2[3] ? byte_1027 : _GEN_4039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5000 = _GEN_8970 == 8'h70 ? _GEN_4996 : _GEN_4036; // @[executor.scala 473:84]
  wire [7:0] _GEN_5001 = _GEN_8970 == 8'h70 ? _GEN_4997 : _GEN_4037; // @[executor.scala 473:84]
  wire [7:0] _GEN_5002 = _GEN_8970 == 8'h70 ? _GEN_4998 : _GEN_4038; // @[executor.scala 473:84]
  wire [7:0] _GEN_5003 = _GEN_8970 == 8'h70 ? _GEN_4999 : _GEN_4039; // @[executor.scala 473:84]
  wire [7:0] _GEN_5004 = mask_2[0] ? byte_1024 : _GEN_4040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5005 = mask_2[1] ? byte_1025 : _GEN_4041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5006 = mask_2[2] ? byte_1026 : _GEN_4042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5007 = mask_2[3] ? byte_1027 : _GEN_4043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5008 = _GEN_8970 == 8'h71 ? _GEN_5004 : _GEN_4040; // @[executor.scala 473:84]
  wire [7:0] _GEN_5009 = _GEN_8970 == 8'h71 ? _GEN_5005 : _GEN_4041; // @[executor.scala 473:84]
  wire [7:0] _GEN_5010 = _GEN_8970 == 8'h71 ? _GEN_5006 : _GEN_4042; // @[executor.scala 473:84]
  wire [7:0] _GEN_5011 = _GEN_8970 == 8'h71 ? _GEN_5007 : _GEN_4043; // @[executor.scala 473:84]
  wire [7:0] _GEN_5012 = mask_2[0] ? byte_1024 : _GEN_4044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5013 = mask_2[1] ? byte_1025 : _GEN_4045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5014 = mask_2[2] ? byte_1026 : _GEN_4046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5015 = mask_2[3] ? byte_1027 : _GEN_4047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5016 = _GEN_8970 == 8'h72 ? _GEN_5012 : _GEN_4044; // @[executor.scala 473:84]
  wire [7:0] _GEN_5017 = _GEN_8970 == 8'h72 ? _GEN_5013 : _GEN_4045; // @[executor.scala 473:84]
  wire [7:0] _GEN_5018 = _GEN_8970 == 8'h72 ? _GEN_5014 : _GEN_4046; // @[executor.scala 473:84]
  wire [7:0] _GEN_5019 = _GEN_8970 == 8'h72 ? _GEN_5015 : _GEN_4047; // @[executor.scala 473:84]
  wire [7:0] _GEN_5020 = mask_2[0] ? byte_1024 : _GEN_4048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5021 = mask_2[1] ? byte_1025 : _GEN_4049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5022 = mask_2[2] ? byte_1026 : _GEN_4050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5023 = mask_2[3] ? byte_1027 : _GEN_4051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5024 = _GEN_8970 == 8'h73 ? _GEN_5020 : _GEN_4048; // @[executor.scala 473:84]
  wire [7:0] _GEN_5025 = _GEN_8970 == 8'h73 ? _GEN_5021 : _GEN_4049; // @[executor.scala 473:84]
  wire [7:0] _GEN_5026 = _GEN_8970 == 8'h73 ? _GEN_5022 : _GEN_4050; // @[executor.scala 473:84]
  wire [7:0] _GEN_5027 = _GEN_8970 == 8'h73 ? _GEN_5023 : _GEN_4051; // @[executor.scala 473:84]
  wire [7:0] _GEN_5028 = mask_2[0] ? byte_1024 : _GEN_4052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5029 = mask_2[1] ? byte_1025 : _GEN_4053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5030 = mask_2[2] ? byte_1026 : _GEN_4054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5031 = mask_2[3] ? byte_1027 : _GEN_4055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5032 = _GEN_8970 == 8'h74 ? _GEN_5028 : _GEN_4052; // @[executor.scala 473:84]
  wire [7:0] _GEN_5033 = _GEN_8970 == 8'h74 ? _GEN_5029 : _GEN_4053; // @[executor.scala 473:84]
  wire [7:0] _GEN_5034 = _GEN_8970 == 8'h74 ? _GEN_5030 : _GEN_4054; // @[executor.scala 473:84]
  wire [7:0] _GEN_5035 = _GEN_8970 == 8'h74 ? _GEN_5031 : _GEN_4055; // @[executor.scala 473:84]
  wire [7:0] _GEN_5036 = mask_2[0] ? byte_1024 : _GEN_4056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5037 = mask_2[1] ? byte_1025 : _GEN_4057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5038 = mask_2[2] ? byte_1026 : _GEN_4058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5039 = mask_2[3] ? byte_1027 : _GEN_4059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5040 = _GEN_8970 == 8'h75 ? _GEN_5036 : _GEN_4056; // @[executor.scala 473:84]
  wire [7:0] _GEN_5041 = _GEN_8970 == 8'h75 ? _GEN_5037 : _GEN_4057; // @[executor.scala 473:84]
  wire [7:0] _GEN_5042 = _GEN_8970 == 8'h75 ? _GEN_5038 : _GEN_4058; // @[executor.scala 473:84]
  wire [7:0] _GEN_5043 = _GEN_8970 == 8'h75 ? _GEN_5039 : _GEN_4059; // @[executor.scala 473:84]
  wire [7:0] _GEN_5044 = mask_2[0] ? byte_1024 : _GEN_4060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5045 = mask_2[1] ? byte_1025 : _GEN_4061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5046 = mask_2[2] ? byte_1026 : _GEN_4062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5047 = mask_2[3] ? byte_1027 : _GEN_4063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5048 = _GEN_8970 == 8'h76 ? _GEN_5044 : _GEN_4060; // @[executor.scala 473:84]
  wire [7:0] _GEN_5049 = _GEN_8970 == 8'h76 ? _GEN_5045 : _GEN_4061; // @[executor.scala 473:84]
  wire [7:0] _GEN_5050 = _GEN_8970 == 8'h76 ? _GEN_5046 : _GEN_4062; // @[executor.scala 473:84]
  wire [7:0] _GEN_5051 = _GEN_8970 == 8'h76 ? _GEN_5047 : _GEN_4063; // @[executor.scala 473:84]
  wire [7:0] _GEN_5052 = mask_2[0] ? byte_1024 : _GEN_4064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5053 = mask_2[1] ? byte_1025 : _GEN_4065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5054 = mask_2[2] ? byte_1026 : _GEN_4066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5055 = mask_2[3] ? byte_1027 : _GEN_4067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5056 = _GEN_8970 == 8'h77 ? _GEN_5052 : _GEN_4064; // @[executor.scala 473:84]
  wire [7:0] _GEN_5057 = _GEN_8970 == 8'h77 ? _GEN_5053 : _GEN_4065; // @[executor.scala 473:84]
  wire [7:0] _GEN_5058 = _GEN_8970 == 8'h77 ? _GEN_5054 : _GEN_4066; // @[executor.scala 473:84]
  wire [7:0] _GEN_5059 = _GEN_8970 == 8'h77 ? _GEN_5055 : _GEN_4067; // @[executor.scala 473:84]
  wire [7:0] _GEN_5060 = mask_2[0] ? byte_1024 : _GEN_4068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5061 = mask_2[1] ? byte_1025 : _GEN_4069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5062 = mask_2[2] ? byte_1026 : _GEN_4070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5063 = mask_2[3] ? byte_1027 : _GEN_4071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5064 = _GEN_8970 == 8'h78 ? _GEN_5060 : _GEN_4068; // @[executor.scala 473:84]
  wire [7:0] _GEN_5065 = _GEN_8970 == 8'h78 ? _GEN_5061 : _GEN_4069; // @[executor.scala 473:84]
  wire [7:0] _GEN_5066 = _GEN_8970 == 8'h78 ? _GEN_5062 : _GEN_4070; // @[executor.scala 473:84]
  wire [7:0] _GEN_5067 = _GEN_8970 == 8'h78 ? _GEN_5063 : _GEN_4071; // @[executor.scala 473:84]
  wire [7:0] _GEN_5068 = mask_2[0] ? byte_1024 : _GEN_4072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5069 = mask_2[1] ? byte_1025 : _GEN_4073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5070 = mask_2[2] ? byte_1026 : _GEN_4074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5071 = mask_2[3] ? byte_1027 : _GEN_4075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5072 = _GEN_8970 == 8'h79 ? _GEN_5068 : _GEN_4072; // @[executor.scala 473:84]
  wire [7:0] _GEN_5073 = _GEN_8970 == 8'h79 ? _GEN_5069 : _GEN_4073; // @[executor.scala 473:84]
  wire [7:0] _GEN_5074 = _GEN_8970 == 8'h79 ? _GEN_5070 : _GEN_4074; // @[executor.scala 473:84]
  wire [7:0] _GEN_5075 = _GEN_8970 == 8'h79 ? _GEN_5071 : _GEN_4075; // @[executor.scala 473:84]
  wire [7:0] _GEN_5076 = mask_2[0] ? byte_1024 : _GEN_4076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5077 = mask_2[1] ? byte_1025 : _GEN_4077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5078 = mask_2[2] ? byte_1026 : _GEN_4078; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5079 = mask_2[3] ? byte_1027 : _GEN_4079; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5080 = _GEN_8970 == 8'h7a ? _GEN_5076 : _GEN_4076; // @[executor.scala 473:84]
  wire [7:0] _GEN_5081 = _GEN_8970 == 8'h7a ? _GEN_5077 : _GEN_4077; // @[executor.scala 473:84]
  wire [7:0] _GEN_5082 = _GEN_8970 == 8'h7a ? _GEN_5078 : _GEN_4078; // @[executor.scala 473:84]
  wire [7:0] _GEN_5083 = _GEN_8970 == 8'h7a ? _GEN_5079 : _GEN_4079; // @[executor.scala 473:84]
  wire [7:0] _GEN_5084 = mask_2[0] ? byte_1024 : _GEN_4080; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5085 = mask_2[1] ? byte_1025 : _GEN_4081; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5086 = mask_2[2] ? byte_1026 : _GEN_4082; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5087 = mask_2[3] ? byte_1027 : _GEN_4083; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5088 = _GEN_8970 == 8'h7b ? _GEN_5084 : _GEN_4080; // @[executor.scala 473:84]
  wire [7:0] _GEN_5089 = _GEN_8970 == 8'h7b ? _GEN_5085 : _GEN_4081; // @[executor.scala 473:84]
  wire [7:0] _GEN_5090 = _GEN_8970 == 8'h7b ? _GEN_5086 : _GEN_4082; // @[executor.scala 473:84]
  wire [7:0] _GEN_5091 = _GEN_8970 == 8'h7b ? _GEN_5087 : _GEN_4083; // @[executor.scala 473:84]
  wire [7:0] _GEN_5092 = mask_2[0] ? byte_1024 : _GEN_4084; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5093 = mask_2[1] ? byte_1025 : _GEN_4085; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5094 = mask_2[2] ? byte_1026 : _GEN_4086; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5095 = mask_2[3] ? byte_1027 : _GEN_4087; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5096 = _GEN_8970 == 8'h7c ? _GEN_5092 : _GEN_4084; // @[executor.scala 473:84]
  wire [7:0] _GEN_5097 = _GEN_8970 == 8'h7c ? _GEN_5093 : _GEN_4085; // @[executor.scala 473:84]
  wire [7:0] _GEN_5098 = _GEN_8970 == 8'h7c ? _GEN_5094 : _GEN_4086; // @[executor.scala 473:84]
  wire [7:0] _GEN_5099 = _GEN_8970 == 8'h7c ? _GEN_5095 : _GEN_4087; // @[executor.scala 473:84]
  wire [7:0] _GEN_5100 = mask_2[0] ? byte_1024 : _GEN_4088; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5101 = mask_2[1] ? byte_1025 : _GEN_4089; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5102 = mask_2[2] ? byte_1026 : _GEN_4090; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5103 = mask_2[3] ? byte_1027 : _GEN_4091; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5104 = _GEN_8970 == 8'h7d ? _GEN_5100 : _GEN_4088; // @[executor.scala 473:84]
  wire [7:0] _GEN_5105 = _GEN_8970 == 8'h7d ? _GEN_5101 : _GEN_4089; // @[executor.scala 473:84]
  wire [7:0] _GEN_5106 = _GEN_8970 == 8'h7d ? _GEN_5102 : _GEN_4090; // @[executor.scala 473:84]
  wire [7:0] _GEN_5107 = _GEN_8970 == 8'h7d ? _GEN_5103 : _GEN_4091; // @[executor.scala 473:84]
  wire [7:0] _GEN_5108 = mask_2[0] ? byte_1024 : _GEN_4092; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5109 = mask_2[1] ? byte_1025 : _GEN_4093; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5110 = mask_2[2] ? byte_1026 : _GEN_4094; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5111 = mask_2[3] ? byte_1027 : _GEN_4095; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5112 = _GEN_8970 == 8'h7e ? _GEN_5108 : _GEN_4092; // @[executor.scala 473:84]
  wire [7:0] _GEN_5113 = _GEN_8970 == 8'h7e ? _GEN_5109 : _GEN_4093; // @[executor.scala 473:84]
  wire [7:0] _GEN_5114 = _GEN_8970 == 8'h7e ? _GEN_5110 : _GEN_4094; // @[executor.scala 473:84]
  wire [7:0] _GEN_5115 = _GEN_8970 == 8'h7e ? _GEN_5111 : _GEN_4095; // @[executor.scala 473:84]
  wire [7:0] _GEN_5116 = mask_2[0] ? byte_1024 : _GEN_4096; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5117 = mask_2[1] ? byte_1025 : _GEN_4097; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5118 = mask_2[2] ? byte_1026 : _GEN_4098; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5119 = mask_2[3] ? byte_1027 : _GEN_4099; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_5120 = _GEN_8970 == 8'h7f ? _GEN_5116 : _GEN_4096; // @[executor.scala 473:84]
  wire [7:0] _GEN_5121 = _GEN_8970 == 8'h7f ? _GEN_5117 : _GEN_4097; // @[executor.scala 473:84]
  wire [7:0] _GEN_5122 = _GEN_8970 == 8'h7f ? _GEN_5118 : _GEN_4098; // @[executor.scala 473:84]
  wire [7:0] _GEN_5123 = _GEN_8970 == 8'h7f ? _GEN_5119 : _GEN_4099; // @[executor.scala 473:84]
  wire [7:0] _GEN_5124 = opcode_2 != 4'h0 ? _GEN_4104 : _GEN_3588; // @[executor.scala 470:55]
  wire [7:0] _GEN_5125 = opcode_2 != 4'h0 ? _GEN_4105 : _GEN_3589; // @[executor.scala 470:55]
  wire [7:0] _GEN_5126 = opcode_2 != 4'h0 ? _GEN_4106 : _GEN_3590; // @[executor.scala 470:55]
  wire [7:0] _GEN_5127 = opcode_2 != 4'h0 ? _GEN_4107 : _GEN_3591; // @[executor.scala 470:55]
  wire [7:0] _GEN_5128 = opcode_2 != 4'h0 ? _GEN_4112 : _GEN_3592; // @[executor.scala 470:55]
  wire [7:0] _GEN_5129 = opcode_2 != 4'h0 ? _GEN_4113 : _GEN_3593; // @[executor.scala 470:55]
  wire [7:0] _GEN_5130 = opcode_2 != 4'h0 ? _GEN_4114 : _GEN_3594; // @[executor.scala 470:55]
  wire [7:0] _GEN_5131 = opcode_2 != 4'h0 ? _GEN_4115 : _GEN_3595; // @[executor.scala 470:55]
  wire [7:0] _GEN_5132 = opcode_2 != 4'h0 ? _GEN_4120 : _GEN_3596; // @[executor.scala 470:55]
  wire [7:0] _GEN_5133 = opcode_2 != 4'h0 ? _GEN_4121 : _GEN_3597; // @[executor.scala 470:55]
  wire [7:0] _GEN_5134 = opcode_2 != 4'h0 ? _GEN_4122 : _GEN_3598; // @[executor.scala 470:55]
  wire [7:0] _GEN_5135 = opcode_2 != 4'h0 ? _GEN_4123 : _GEN_3599; // @[executor.scala 470:55]
  wire [7:0] _GEN_5136 = opcode_2 != 4'h0 ? _GEN_4128 : _GEN_3600; // @[executor.scala 470:55]
  wire [7:0] _GEN_5137 = opcode_2 != 4'h0 ? _GEN_4129 : _GEN_3601; // @[executor.scala 470:55]
  wire [7:0] _GEN_5138 = opcode_2 != 4'h0 ? _GEN_4130 : _GEN_3602; // @[executor.scala 470:55]
  wire [7:0] _GEN_5139 = opcode_2 != 4'h0 ? _GEN_4131 : _GEN_3603; // @[executor.scala 470:55]
  wire [7:0] _GEN_5140 = opcode_2 != 4'h0 ? _GEN_4136 : _GEN_3604; // @[executor.scala 470:55]
  wire [7:0] _GEN_5141 = opcode_2 != 4'h0 ? _GEN_4137 : _GEN_3605; // @[executor.scala 470:55]
  wire [7:0] _GEN_5142 = opcode_2 != 4'h0 ? _GEN_4138 : _GEN_3606; // @[executor.scala 470:55]
  wire [7:0] _GEN_5143 = opcode_2 != 4'h0 ? _GEN_4139 : _GEN_3607; // @[executor.scala 470:55]
  wire [7:0] _GEN_5144 = opcode_2 != 4'h0 ? _GEN_4144 : _GEN_3608; // @[executor.scala 470:55]
  wire [7:0] _GEN_5145 = opcode_2 != 4'h0 ? _GEN_4145 : _GEN_3609; // @[executor.scala 470:55]
  wire [7:0] _GEN_5146 = opcode_2 != 4'h0 ? _GEN_4146 : _GEN_3610; // @[executor.scala 470:55]
  wire [7:0] _GEN_5147 = opcode_2 != 4'h0 ? _GEN_4147 : _GEN_3611; // @[executor.scala 470:55]
  wire [7:0] _GEN_5148 = opcode_2 != 4'h0 ? _GEN_4152 : _GEN_3612; // @[executor.scala 470:55]
  wire [7:0] _GEN_5149 = opcode_2 != 4'h0 ? _GEN_4153 : _GEN_3613; // @[executor.scala 470:55]
  wire [7:0] _GEN_5150 = opcode_2 != 4'h0 ? _GEN_4154 : _GEN_3614; // @[executor.scala 470:55]
  wire [7:0] _GEN_5151 = opcode_2 != 4'h0 ? _GEN_4155 : _GEN_3615; // @[executor.scala 470:55]
  wire [7:0] _GEN_5152 = opcode_2 != 4'h0 ? _GEN_4160 : _GEN_3616; // @[executor.scala 470:55]
  wire [7:0] _GEN_5153 = opcode_2 != 4'h0 ? _GEN_4161 : _GEN_3617; // @[executor.scala 470:55]
  wire [7:0] _GEN_5154 = opcode_2 != 4'h0 ? _GEN_4162 : _GEN_3618; // @[executor.scala 470:55]
  wire [7:0] _GEN_5155 = opcode_2 != 4'h0 ? _GEN_4163 : _GEN_3619; // @[executor.scala 470:55]
  wire [7:0] _GEN_5156 = opcode_2 != 4'h0 ? _GEN_4168 : _GEN_3620; // @[executor.scala 470:55]
  wire [7:0] _GEN_5157 = opcode_2 != 4'h0 ? _GEN_4169 : _GEN_3621; // @[executor.scala 470:55]
  wire [7:0] _GEN_5158 = opcode_2 != 4'h0 ? _GEN_4170 : _GEN_3622; // @[executor.scala 470:55]
  wire [7:0] _GEN_5159 = opcode_2 != 4'h0 ? _GEN_4171 : _GEN_3623; // @[executor.scala 470:55]
  wire [7:0] _GEN_5160 = opcode_2 != 4'h0 ? _GEN_4176 : _GEN_3624; // @[executor.scala 470:55]
  wire [7:0] _GEN_5161 = opcode_2 != 4'h0 ? _GEN_4177 : _GEN_3625; // @[executor.scala 470:55]
  wire [7:0] _GEN_5162 = opcode_2 != 4'h0 ? _GEN_4178 : _GEN_3626; // @[executor.scala 470:55]
  wire [7:0] _GEN_5163 = opcode_2 != 4'h0 ? _GEN_4179 : _GEN_3627; // @[executor.scala 470:55]
  wire [7:0] _GEN_5164 = opcode_2 != 4'h0 ? _GEN_4184 : _GEN_3628; // @[executor.scala 470:55]
  wire [7:0] _GEN_5165 = opcode_2 != 4'h0 ? _GEN_4185 : _GEN_3629; // @[executor.scala 470:55]
  wire [7:0] _GEN_5166 = opcode_2 != 4'h0 ? _GEN_4186 : _GEN_3630; // @[executor.scala 470:55]
  wire [7:0] _GEN_5167 = opcode_2 != 4'h0 ? _GEN_4187 : _GEN_3631; // @[executor.scala 470:55]
  wire [7:0] _GEN_5168 = opcode_2 != 4'h0 ? _GEN_4192 : _GEN_3632; // @[executor.scala 470:55]
  wire [7:0] _GEN_5169 = opcode_2 != 4'h0 ? _GEN_4193 : _GEN_3633; // @[executor.scala 470:55]
  wire [7:0] _GEN_5170 = opcode_2 != 4'h0 ? _GEN_4194 : _GEN_3634; // @[executor.scala 470:55]
  wire [7:0] _GEN_5171 = opcode_2 != 4'h0 ? _GEN_4195 : _GEN_3635; // @[executor.scala 470:55]
  wire [7:0] _GEN_5172 = opcode_2 != 4'h0 ? _GEN_4200 : _GEN_3636; // @[executor.scala 470:55]
  wire [7:0] _GEN_5173 = opcode_2 != 4'h0 ? _GEN_4201 : _GEN_3637; // @[executor.scala 470:55]
  wire [7:0] _GEN_5174 = opcode_2 != 4'h0 ? _GEN_4202 : _GEN_3638; // @[executor.scala 470:55]
  wire [7:0] _GEN_5175 = opcode_2 != 4'h0 ? _GEN_4203 : _GEN_3639; // @[executor.scala 470:55]
  wire [7:0] _GEN_5176 = opcode_2 != 4'h0 ? _GEN_4208 : _GEN_3640; // @[executor.scala 470:55]
  wire [7:0] _GEN_5177 = opcode_2 != 4'h0 ? _GEN_4209 : _GEN_3641; // @[executor.scala 470:55]
  wire [7:0] _GEN_5178 = opcode_2 != 4'h0 ? _GEN_4210 : _GEN_3642; // @[executor.scala 470:55]
  wire [7:0] _GEN_5179 = opcode_2 != 4'h0 ? _GEN_4211 : _GEN_3643; // @[executor.scala 470:55]
  wire [7:0] _GEN_5180 = opcode_2 != 4'h0 ? _GEN_4216 : _GEN_3644; // @[executor.scala 470:55]
  wire [7:0] _GEN_5181 = opcode_2 != 4'h0 ? _GEN_4217 : _GEN_3645; // @[executor.scala 470:55]
  wire [7:0] _GEN_5182 = opcode_2 != 4'h0 ? _GEN_4218 : _GEN_3646; // @[executor.scala 470:55]
  wire [7:0] _GEN_5183 = opcode_2 != 4'h0 ? _GEN_4219 : _GEN_3647; // @[executor.scala 470:55]
  wire [7:0] _GEN_5184 = opcode_2 != 4'h0 ? _GEN_4224 : _GEN_3648; // @[executor.scala 470:55]
  wire [7:0] _GEN_5185 = opcode_2 != 4'h0 ? _GEN_4225 : _GEN_3649; // @[executor.scala 470:55]
  wire [7:0] _GEN_5186 = opcode_2 != 4'h0 ? _GEN_4226 : _GEN_3650; // @[executor.scala 470:55]
  wire [7:0] _GEN_5187 = opcode_2 != 4'h0 ? _GEN_4227 : _GEN_3651; // @[executor.scala 470:55]
  wire [7:0] _GEN_5188 = opcode_2 != 4'h0 ? _GEN_4232 : _GEN_3652; // @[executor.scala 470:55]
  wire [7:0] _GEN_5189 = opcode_2 != 4'h0 ? _GEN_4233 : _GEN_3653; // @[executor.scala 470:55]
  wire [7:0] _GEN_5190 = opcode_2 != 4'h0 ? _GEN_4234 : _GEN_3654; // @[executor.scala 470:55]
  wire [7:0] _GEN_5191 = opcode_2 != 4'h0 ? _GEN_4235 : _GEN_3655; // @[executor.scala 470:55]
  wire [7:0] _GEN_5192 = opcode_2 != 4'h0 ? _GEN_4240 : _GEN_3656; // @[executor.scala 470:55]
  wire [7:0] _GEN_5193 = opcode_2 != 4'h0 ? _GEN_4241 : _GEN_3657; // @[executor.scala 470:55]
  wire [7:0] _GEN_5194 = opcode_2 != 4'h0 ? _GEN_4242 : _GEN_3658; // @[executor.scala 470:55]
  wire [7:0] _GEN_5195 = opcode_2 != 4'h0 ? _GEN_4243 : _GEN_3659; // @[executor.scala 470:55]
  wire [7:0] _GEN_5196 = opcode_2 != 4'h0 ? _GEN_4248 : _GEN_3660; // @[executor.scala 470:55]
  wire [7:0] _GEN_5197 = opcode_2 != 4'h0 ? _GEN_4249 : _GEN_3661; // @[executor.scala 470:55]
  wire [7:0] _GEN_5198 = opcode_2 != 4'h0 ? _GEN_4250 : _GEN_3662; // @[executor.scala 470:55]
  wire [7:0] _GEN_5199 = opcode_2 != 4'h0 ? _GEN_4251 : _GEN_3663; // @[executor.scala 470:55]
  wire [7:0] _GEN_5200 = opcode_2 != 4'h0 ? _GEN_4256 : _GEN_3664; // @[executor.scala 470:55]
  wire [7:0] _GEN_5201 = opcode_2 != 4'h0 ? _GEN_4257 : _GEN_3665; // @[executor.scala 470:55]
  wire [7:0] _GEN_5202 = opcode_2 != 4'h0 ? _GEN_4258 : _GEN_3666; // @[executor.scala 470:55]
  wire [7:0] _GEN_5203 = opcode_2 != 4'h0 ? _GEN_4259 : _GEN_3667; // @[executor.scala 470:55]
  wire [7:0] _GEN_5204 = opcode_2 != 4'h0 ? _GEN_4264 : _GEN_3668; // @[executor.scala 470:55]
  wire [7:0] _GEN_5205 = opcode_2 != 4'h0 ? _GEN_4265 : _GEN_3669; // @[executor.scala 470:55]
  wire [7:0] _GEN_5206 = opcode_2 != 4'h0 ? _GEN_4266 : _GEN_3670; // @[executor.scala 470:55]
  wire [7:0] _GEN_5207 = opcode_2 != 4'h0 ? _GEN_4267 : _GEN_3671; // @[executor.scala 470:55]
  wire [7:0] _GEN_5208 = opcode_2 != 4'h0 ? _GEN_4272 : _GEN_3672; // @[executor.scala 470:55]
  wire [7:0] _GEN_5209 = opcode_2 != 4'h0 ? _GEN_4273 : _GEN_3673; // @[executor.scala 470:55]
  wire [7:0] _GEN_5210 = opcode_2 != 4'h0 ? _GEN_4274 : _GEN_3674; // @[executor.scala 470:55]
  wire [7:0] _GEN_5211 = opcode_2 != 4'h0 ? _GEN_4275 : _GEN_3675; // @[executor.scala 470:55]
  wire [7:0] _GEN_5212 = opcode_2 != 4'h0 ? _GEN_4280 : _GEN_3676; // @[executor.scala 470:55]
  wire [7:0] _GEN_5213 = opcode_2 != 4'h0 ? _GEN_4281 : _GEN_3677; // @[executor.scala 470:55]
  wire [7:0] _GEN_5214 = opcode_2 != 4'h0 ? _GEN_4282 : _GEN_3678; // @[executor.scala 470:55]
  wire [7:0] _GEN_5215 = opcode_2 != 4'h0 ? _GEN_4283 : _GEN_3679; // @[executor.scala 470:55]
  wire [7:0] _GEN_5216 = opcode_2 != 4'h0 ? _GEN_4288 : _GEN_3680; // @[executor.scala 470:55]
  wire [7:0] _GEN_5217 = opcode_2 != 4'h0 ? _GEN_4289 : _GEN_3681; // @[executor.scala 470:55]
  wire [7:0] _GEN_5218 = opcode_2 != 4'h0 ? _GEN_4290 : _GEN_3682; // @[executor.scala 470:55]
  wire [7:0] _GEN_5219 = opcode_2 != 4'h0 ? _GEN_4291 : _GEN_3683; // @[executor.scala 470:55]
  wire [7:0] _GEN_5220 = opcode_2 != 4'h0 ? _GEN_4296 : _GEN_3684; // @[executor.scala 470:55]
  wire [7:0] _GEN_5221 = opcode_2 != 4'h0 ? _GEN_4297 : _GEN_3685; // @[executor.scala 470:55]
  wire [7:0] _GEN_5222 = opcode_2 != 4'h0 ? _GEN_4298 : _GEN_3686; // @[executor.scala 470:55]
  wire [7:0] _GEN_5223 = opcode_2 != 4'h0 ? _GEN_4299 : _GEN_3687; // @[executor.scala 470:55]
  wire [7:0] _GEN_5224 = opcode_2 != 4'h0 ? _GEN_4304 : _GEN_3688; // @[executor.scala 470:55]
  wire [7:0] _GEN_5225 = opcode_2 != 4'h0 ? _GEN_4305 : _GEN_3689; // @[executor.scala 470:55]
  wire [7:0] _GEN_5226 = opcode_2 != 4'h0 ? _GEN_4306 : _GEN_3690; // @[executor.scala 470:55]
  wire [7:0] _GEN_5227 = opcode_2 != 4'h0 ? _GEN_4307 : _GEN_3691; // @[executor.scala 470:55]
  wire [7:0] _GEN_5228 = opcode_2 != 4'h0 ? _GEN_4312 : _GEN_3692; // @[executor.scala 470:55]
  wire [7:0] _GEN_5229 = opcode_2 != 4'h0 ? _GEN_4313 : _GEN_3693; // @[executor.scala 470:55]
  wire [7:0] _GEN_5230 = opcode_2 != 4'h0 ? _GEN_4314 : _GEN_3694; // @[executor.scala 470:55]
  wire [7:0] _GEN_5231 = opcode_2 != 4'h0 ? _GEN_4315 : _GEN_3695; // @[executor.scala 470:55]
  wire [7:0] _GEN_5232 = opcode_2 != 4'h0 ? _GEN_4320 : _GEN_3696; // @[executor.scala 470:55]
  wire [7:0] _GEN_5233 = opcode_2 != 4'h0 ? _GEN_4321 : _GEN_3697; // @[executor.scala 470:55]
  wire [7:0] _GEN_5234 = opcode_2 != 4'h0 ? _GEN_4322 : _GEN_3698; // @[executor.scala 470:55]
  wire [7:0] _GEN_5235 = opcode_2 != 4'h0 ? _GEN_4323 : _GEN_3699; // @[executor.scala 470:55]
  wire [7:0] _GEN_5236 = opcode_2 != 4'h0 ? _GEN_4328 : _GEN_3700; // @[executor.scala 470:55]
  wire [7:0] _GEN_5237 = opcode_2 != 4'h0 ? _GEN_4329 : _GEN_3701; // @[executor.scala 470:55]
  wire [7:0] _GEN_5238 = opcode_2 != 4'h0 ? _GEN_4330 : _GEN_3702; // @[executor.scala 470:55]
  wire [7:0] _GEN_5239 = opcode_2 != 4'h0 ? _GEN_4331 : _GEN_3703; // @[executor.scala 470:55]
  wire [7:0] _GEN_5240 = opcode_2 != 4'h0 ? _GEN_4336 : _GEN_3704; // @[executor.scala 470:55]
  wire [7:0] _GEN_5241 = opcode_2 != 4'h0 ? _GEN_4337 : _GEN_3705; // @[executor.scala 470:55]
  wire [7:0] _GEN_5242 = opcode_2 != 4'h0 ? _GEN_4338 : _GEN_3706; // @[executor.scala 470:55]
  wire [7:0] _GEN_5243 = opcode_2 != 4'h0 ? _GEN_4339 : _GEN_3707; // @[executor.scala 470:55]
  wire [7:0] _GEN_5244 = opcode_2 != 4'h0 ? _GEN_4344 : _GEN_3708; // @[executor.scala 470:55]
  wire [7:0] _GEN_5245 = opcode_2 != 4'h0 ? _GEN_4345 : _GEN_3709; // @[executor.scala 470:55]
  wire [7:0] _GEN_5246 = opcode_2 != 4'h0 ? _GEN_4346 : _GEN_3710; // @[executor.scala 470:55]
  wire [7:0] _GEN_5247 = opcode_2 != 4'h0 ? _GEN_4347 : _GEN_3711; // @[executor.scala 470:55]
  wire [7:0] _GEN_5248 = opcode_2 != 4'h0 ? _GEN_4352 : _GEN_3712; // @[executor.scala 470:55]
  wire [7:0] _GEN_5249 = opcode_2 != 4'h0 ? _GEN_4353 : _GEN_3713; // @[executor.scala 470:55]
  wire [7:0] _GEN_5250 = opcode_2 != 4'h0 ? _GEN_4354 : _GEN_3714; // @[executor.scala 470:55]
  wire [7:0] _GEN_5251 = opcode_2 != 4'h0 ? _GEN_4355 : _GEN_3715; // @[executor.scala 470:55]
  wire [7:0] _GEN_5252 = opcode_2 != 4'h0 ? _GEN_4360 : _GEN_3716; // @[executor.scala 470:55]
  wire [7:0] _GEN_5253 = opcode_2 != 4'h0 ? _GEN_4361 : _GEN_3717; // @[executor.scala 470:55]
  wire [7:0] _GEN_5254 = opcode_2 != 4'h0 ? _GEN_4362 : _GEN_3718; // @[executor.scala 470:55]
  wire [7:0] _GEN_5255 = opcode_2 != 4'h0 ? _GEN_4363 : _GEN_3719; // @[executor.scala 470:55]
  wire [7:0] _GEN_5256 = opcode_2 != 4'h0 ? _GEN_4368 : _GEN_3720; // @[executor.scala 470:55]
  wire [7:0] _GEN_5257 = opcode_2 != 4'h0 ? _GEN_4369 : _GEN_3721; // @[executor.scala 470:55]
  wire [7:0] _GEN_5258 = opcode_2 != 4'h0 ? _GEN_4370 : _GEN_3722; // @[executor.scala 470:55]
  wire [7:0] _GEN_5259 = opcode_2 != 4'h0 ? _GEN_4371 : _GEN_3723; // @[executor.scala 470:55]
  wire [7:0] _GEN_5260 = opcode_2 != 4'h0 ? _GEN_4376 : _GEN_3724; // @[executor.scala 470:55]
  wire [7:0] _GEN_5261 = opcode_2 != 4'h0 ? _GEN_4377 : _GEN_3725; // @[executor.scala 470:55]
  wire [7:0] _GEN_5262 = opcode_2 != 4'h0 ? _GEN_4378 : _GEN_3726; // @[executor.scala 470:55]
  wire [7:0] _GEN_5263 = opcode_2 != 4'h0 ? _GEN_4379 : _GEN_3727; // @[executor.scala 470:55]
  wire [7:0] _GEN_5264 = opcode_2 != 4'h0 ? _GEN_4384 : _GEN_3728; // @[executor.scala 470:55]
  wire [7:0] _GEN_5265 = opcode_2 != 4'h0 ? _GEN_4385 : _GEN_3729; // @[executor.scala 470:55]
  wire [7:0] _GEN_5266 = opcode_2 != 4'h0 ? _GEN_4386 : _GEN_3730; // @[executor.scala 470:55]
  wire [7:0] _GEN_5267 = opcode_2 != 4'h0 ? _GEN_4387 : _GEN_3731; // @[executor.scala 470:55]
  wire [7:0] _GEN_5268 = opcode_2 != 4'h0 ? _GEN_4392 : _GEN_3732; // @[executor.scala 470:55]
  wire [7:0] _GEN_5269 = opcode_2 != 4'h0 ? _GEN_4393 : _GEN_3733; // @[executor.scala 470:55]
  wire [7:0] _GEN_5270 = opcode_2 != 4'h0 ? _GEN_4394 : _GEN_3734; // @[executor.scala 470:55]
  wire [7:0] _GEN_5271 = opcode_2 != 4'h0 ? _GEN_4395 : _GEN_3735; // @[executor.scala 470:55]
  wire [7:0] _GEN_5272 = opcode_2 != 4'h0 ? _GEN_4400 : _GEN_3736; // @[executor.scala 470:55]
  wire [7:0] _GEN_5273 = opcode_2 != 4'h0 ? _GEN_4401 : _GEN_3737; // @[executor.scala 470:55]
  wire [7:0] _GEN_5274 = opcode_2 != 4'h0 ? _GEN_4402 : _GEN_3738; // @[executor.scala 470:55]
  wire [7:0] _GEN_5275 = opcode_2 != 4'h0 ? _GEN_4403 : _GEN_3739; // @[executor.scala 470:55]
  wire [7:0] _GEN_5276 = opcode_2 != 4'h0 ? _GEN_4408 : _GEN_3740; // @[executor.scala 470:55]
  wire [7:0] _GEN_5277 = opcode_2 != 4'h0 ? _GEN_4409 : _GEN_3741; // @[executor.scala 470:55]
  wire [7:0] _GEN_5278 = opcode_2 != 4'h0 ? _GEN_4410 : _GEN_3742; // @[executor.scala 470:55]
  wire [7:0] _GEN_5279 = opcode_2 != 4'h0 ? _GEN_4411 : _GEN_3743; // @[executor.scala 470:55]
  wire [7:0] _GEN_5280 = opcode_2 != 4'h0 ? _GEN_4416 : _GEN_3744; // @[executor.scala 470:55]
  wire [7:0] _GEN_5281 = opcode_2 != 4'h0 ? _GEN_4417 : _GEN_3745; // @[executor.scala 470:55]
  wire [7:0] _GEN_5282 = opcode_2 != 4'h0 ? _GEN_4418 : _GEN_3746; // @[executor.scala 470:55]
  wire [7:0] _GEN_5283 = opcode_2 != 4'h0 ? _GEN_4419 : _GEN_3747; // @[executor.scala 470:55]
  wire [7:0] _GEN_5284 = opcode_2 != 4'h0 ? _GEN_4424 : _GEN_3748; // @[executor.scala 470:55]
  wire [7:0] _GEN_5285 = opcode_2 != 4'h0 ? _GEN_4425 : _GEN_3749; // @[executor.scala 470:55]
  wire [7:0] _GEN_5286 = opcode_2 != 4'h0 ? _GEN_4426 : _GEN_3750; // @[executor.scala 470:55]
  wire [7:0] _GEN_5287 = opcode_2 != 4'h0 ? _GEN_4427 : _GEN_3751; // @[executor.scala 470:55]
  wire [7:0] _GEN_5288 = opcode_2 != 4'h0 ? _GEN_4432 : _GEN_3752; // @[executor.scala 470:55]
  wire [7:0] _GEN_5289 = opcode_2 != 4'h0 ? _GEN_4433 : _GEN_3753; // @[executor.scala 470:55]
  wire [7:0] _GEN_5290 = opcode_2 != 4'h0 ? _GEN_4434 : _GEN_3754; // @[executor.scala 470:55]
  wire [7:0] _GEN_5291 = opcode_2 != 4'h0 ? _GEN_4435 : _GEN_3755; // @[executor.scala 470:55]
  wire [7:0] _GEN_5292 = opcode_2 != 4'h0 ? _GEN_4440 : _GEN_3756; // @[executor.scala 470:55]
  wire [7:0] _GEN_5293 = opcode_2 != 4'h0 ? _GEN_4441 : _GEN_3757; // @[executor.scala 470:55]
  wire [7:0] _GEN_5294 = opcode_2 != 4'h0 ? _GEN_4442 : _GEN_3758; // @[executor.scala 470:55]
  wire [7:0] _GEN_5295 = opcode_2 != 4'h0 ? _GEN_4443 : _GEN_3759; // @[executor.scala 470:55]
  wire [7:0] _GEN_5296 = opcode_2 != 4'h0 ? _GEN_4448 : _GEN_3760; // @[executor.scala 470:55]
  wire [7:0] _GEN_5297 = opcode_2 != 4'h0 ? _GEN_4449 : _GEN_3761; // @[executor.scala 470:55]
  wire [7:0] _GEN_5298 = opcode_2 != 4'h0 ? _GEN_4450 : _GEN_3762; // @[executor.scala 470:55]
  wire [7:0] _GEN_5299 = opcode_2 != 4'h0 ? _GEN_4451 : _GEN_3763; // @[executor.scala 470:55]
  wire [7:0] _GEN_5300 = opcode_2 != 4'h0 ? _GEN_4456 : _GEN_3764; // @[executor.scala 470:55]
  wire [7:0] _GEN_5301 = opcode_2 != 4'h0 ? _GEN_4457 : _GEN_3765; // @[executor.scala 470:55]
  wire [7:0] _GEN_5302 = opcode_2 != 4'h0 ? _GEN_4458 : _GEN_3766; // @[executor.scala 470:55]
  wire [7:0] _GEN_5303 = opcode_2 != 4'h0 ? _GEN_4459 : _GEN_3767; // @[executor.scala 470:55]
  wire [7:0] _GEN_5304 = opcode_2 != 4'h0 ? _GEN_4464 : _GEN_3768; // @[executor.scala 470:55]
  wire [7:0] _GEN_5305 = opcode_2 != 4'h0 ? _GEN_4465 : _GEN_3769; // @[executor.scala 470:55]
  wire [7:0] _GEN_5306 = opcode_2 != 4'h0 ? _GEN_4466 : _GEN_3770; // @[executor.scala 470:55]
  wire [7:0] _GEN_5307 = opcode_2 != 4'h0 ? _GEN_4467 : _GEN_3771; // @[executor.scala 470:55]
  wire [7:0] _GEN_5308 = opcode_2 != 4'h0 ? _GEN_4472 : _GEN_3772; // @[executor.scala 470:55]
  wire [7:0] _GEN_5309 = opcode_2 != 4'h0 ? _GEN_4473 : _GEN_3773; // @[executor.scala 470:55]
  wire [7:0] _GEN_5310 = opcode_2 != 4'h0 ? _GEN_4474 : _GEN_3774; // @[executor.scala 470:55]
  wire [7:0] _GEN_5311 = opcode_2 != 4'h0 ? _GEN_4475 : _GEN_3775; // @[executor.scala 470:55]
  wire [7:0] _GEN_5312 = opcode_2 != 4'h0 ? _GEN_4480 : _GEN_3776; // @[executor.scala 470:55]
  wire [7:0] _GEN_5313 = opcode_2 != 4'h0 ? _GEN_4481 : _GEN_3777; // @[executor.scala 470:55]
  wire [7:0] _GEN_5314 = opcode_2 != 4'h0 ? _GEN_4482 : _GEN_3778; // @[executor.scala 470:55]
  wire [7:0] _GEN_5315 = opcode_2 != 4'h0 ? _GEN_4483 : _GEN_3779; // @[executor.scala 470:55]
  wire [7:0] _GEN_5316 = opcode_2 != 4'h0 ? _GEN_4488 : _GEN_3780; // @[executor.scala 470:55]
  wire [7:0] _GEN_5317 = opcode_2 != 4'h0 ? _GEN_4489 : _GEN_3781; // @[executor.scala 470:55]
  wire [7:0] _GEN_5318 = opcode_2 != 4'h0 ? _GEN_4490 : _GEN_3782; // @[executor.scala 470:55]
  wire [7:0] _GEN_5319 = opcode_2 != 4'h0 ? _GEN_4491 : _GEN_3783; // @[executor.scala 470:55]
  wire [7:0] _GEN_5320 = opcode_2 != 4'h0 ? _GEN_4496 : _GEN_3784; // @[executor.scala 470:55]
  wire [7:0] _GEN_5321 = opcode_2 != 4'h0 ? _GEN_4497 : _GEN_3785; // @[executor.scala 470:55]
  wire [7:0] _GEN_5322 = opcode_2 != 4'h0 ? _GEN_4498 : _GEN_3786; // @[executor.scala 470:55]
  wire [7:0] _GEN_5323 = opcode_2 != 4'h0 ? _GEN_4499 : _GEN_3787; // @[executor.scala 470:55]
  wire [7:0] _GEN_5324 = opcode_2 != 4'h0 ? _GEN_4504 : _GEN_3788; // @[executor.scala 470:55]
  wire [7:0] _GEN_5325 = opcode_2 != 4'h0 ? _GEN_4505 : _GEN_3789; // @[executor.scala 470:55]
  wire [7:0] _GEN_5326 = opcode_2 != 4'h0 ? _GEN_4506 : _GEN_3790; // @[executor.scala 470:55]
  wire [7:0] _GEN_5327 = opcode_2 != 4'h0 ? _GEN_4507 : _GEN_3791; // @[executor.scala 470:55]
  wire [7:0] _GEN_5328 = opcode_2 != 4'h0 ? _GEN_4512 : _GEN_3792; // @[executor.scala 470:55]
  wire [7:0] _GEN_5329 = opcode_2 != 4'h0 ? _GEN_4513 : _GEN_3793; // @[executor.scala 470:55]
  wire [7:0] _GEN_5330 = opcode_2 != 4'h0 ? _GEN_4514 : _GEN_3794; // @[executor.scala 470:55]
  wire [7:0] _GEN_5331 = opcode_2 != 4'h0 ? _GEN_4515 : _GEN_3795; // @[executor.scala 470:55]
  wire [7:0] _GEN_5332 = opcode_2 != 4'h0 ? _GEN_4520 : _GEN_3796; // @[executor.scala 470:55]
  wire [7:0] _GEN_5333 = opcode_2 != 4'h0 ? _GEN_4521 : _GEN_3797; // @[executor.scala 470:55]
  wire [7:0] _GEN_5334 = opcode_2 != 4'h0 ? _GEN_4522 : _GEN_3798; // @[executor.scala 470:55]
  wire [7:0] _GEN_5335 = opcode_2 != 4'h0 ? _GEN_4523 : _GEN_3799; // @[executor.scala 470:55]
  wire [7:0] _GEN_5336 = opcode_2 != 4'h0 ? _GEN_4528 : _GEN_3800; // @[executor.scala 470:55]
  wire [7:0] _GEN_5337 = opcode_2 != 4'h0 ? _GEN_4529 : _GEN_3801; // @[executor.scala 470:55]
  wire [7:0] _GEN_5338 = opcode_2 != 4'h0 ? _GEN_4530 : _GEN_3802; // @[executor.scala 470:55]
  wire [7:0] _GEN_5339 = opcode_2 != 4'h0 ? _GEN_4531 : _GEN_3803; // @[executor.scala 470:55]
  wire [7:0] _GEN_5340 = opcode_2 != 4'h0 ? _GEN_4536 : _GEN_3804; // @[executor.scala 470:55]
  wire [7:0] _GEN_5341 = opcode_2 != 4'h0 ? _GEN_4537 : _GEN_3805; // @[executor.scala 470:55]
  wire [7:0] _GEN_5342 = opcode_2 != 4'h0 ? _GEN_4538 : _GEN_3806; // @[executor.scala 470:55]
  wire [7:0] _GEN_5343 = opcode_2 != 4'h0 ? _GEN_4539 : _GEN_3807; // @[executor.scala 470:55]
  wire [7:0] _GEN_5344 = opcode_2 != 4'h0 ? _GEN_4544 : _GEN_3808; // @[executor.scala 470:55]
  wire [7:0] _GEN_5345 = opcode_2 != 4'h0 ? _GEN_4545 : _GEN_3809; // @[executor.scala 470:55]
  wire [7:0] _GEN_5346 = opcode_2 != 4'h0 ? _GEN_4546 : _GEN_3810; // @[executor.scala 470:55]
  wire [7:0] _GEN_5347 = opcode_2 != 4'h0 ? _GEN_4547 : _GEN_3811; // @[executor.scala 470:55]
  wire [7:0] _GEN_5348 = opcode_2 != 4'h0 ? _GEN_4552 : _GEN_3812; // @[executor.scala 470:55]
  wire [7:0] _GEN_5349 = opcode_2 != 4'h0 ? _GEN_4553 : _GEN_3813; // @[executor.scala 470:55]
  wire [7:0] _GEN_5350 = opcode_2 != 4'h0 ? _GEN_4554 : _GEN_3814; // @[executor.scala 470:55]
  wire [7:0] _GEN_5351 = opcode_2 != 4'h0 ? _GEN_4555 : _GEN_3815; // @[executor.scala 470:55]
  wire [7:0] _GEN_5352 = opcode_2 != 4'h0 ? _GEN_4560 : _GEN_3816; // @[executor.scala 470:55]
  wire [7:0] _GEN_5353 = opcode_2 != 4'h0 ? _GEN_4561 : _GEN_3817; // @[executor.scala 470:55]
  wire [7:0] _GEN_5354 = opcode_2 != 4'h0 ? _GEN_4562 : _GEN_3818; // @[executor.scala 470:55]
  wire [7:0] _GEN_5355 = opcode_2 != 4'h0 ? _GEN_4563 : _GEN_3819; // @[executor.scala 470:55]
  wire [7:0] _GEN_5356 = opcode_2 != 4'h0 ? _GEN_4568 : _GEN_3820; // @[executor.scala 470:55]
  wire [7:0] _GEN_5357 = opcode_2 != 4'h0 ? _GEN_4569 : _GEN_3821; // @[executor.scala 470:55]
  wire [7:0] _GEN_5358 = opcode_2 != 4'h0 ? _GEN_4570 : _GEN_3822; // @[executor.scala 470:55]
  wire [7:0] _GEN_5359 = opcode_2 != 4'h0 ? _GEN_4571 : _GEN_3823; // @[executor.scala 470:55]
  wire [7:0] _GEN_5360 = opcode_2 != 4'h0 ? _GEN_4576 : _GEN_3824; // @[executor.scala 470:55]
  wire [7:0] _GEN_5361 = opcode_2 != 4'h0 ? _GEN_4577 : _GEN_3825; // @[executor.scala 470:55]
  wire [7:0] _GEN_5362 = opcode_2 != 4'h0 ? _GEN_4578 : _GEN_3826; // @[executor.scala 470:55]
  wire [7:0] _GEN_5363 = opcode_2 != 4'h0 ? _GEN_4579 : _GEN_3827; // @[executor.scala 470:55]
  wire [7:0] _GEN_5364 = opcode_2 != 4'h0 ? _GEN_4584 : _GEN_3828; // @[executor.scala 470:55]
  wire [7:0] _GEN_5365 = opcode_2 != 4'h0 ? _GEN_4585 : _GEN_3829; // @[executor.scala 470:55]
  wire [7:0] _GEN_5366 = opcode_2 != 4'h0 ? _GEN_4586 : _GEN_3830; // @[executor.scala 470:55]
  wire [7:0] _GEN_5367 = opcode_2 != 4'h0 ? _GEN_4587 : _GEN_3831; // @[executor.scala 470:55]
  wire [7:0] _GEN_5368 = opcode_2 != 4'h0 ? _GEN_4592 : _GEN_3832; // @[executor.scala 470:55]
  wire [7:0] _GEN_5369 = opcode_2 != 4'h0 ? _GEN_4593 : _GEN_3833; // @[executor.scala 470:55]
  wire [7:0] _GEN_5370 = opcode_2 != 4'h0 ? _GEN_4594 : _GEN_3834; // @[executor.scala 470:55]
  wire [7:0] _GEN_5371 = opcode_2 != 4'h0 ? _GEN_4595 : _GEN_3835; // @[executor.scala 470:55]
  wire [7:0] _GEN_5372 = opcode_2 != 4'h0 ? _GEN_4600 : _GEN_3836; // @[executor.scala 470:55]
  wire [7:0] _GEN_5373 = opcode_2 != 4'h0 ? _GEN_4601 : _GEN_3837; // @[executor.scala 470:55]
  wire [7:0] _GEN_5374 = opcode_2 != 4'h0 ? _GEN_4602 : _GEN_3838; // @[executor.scala 470:55]
  wire [7:0] _GEN_5375 = opcode_2 != 4'h0 ? _GEN_4603 : _GEN_3839; // @[executor.scala 470:55]
  wire [7:0] _GEN_5376 = opcode_2 != 4'h0 ? _GEN_4608 : _GEN_3840; // @[executor.scala 470:55]
  wire [7:0] _GEN_5377 = opcode_2 != 4'h0 ? _GEN_4609 : _GEN_3841; // @[executor.scala 470:55]
  wire [7:0] _GEN_5378 = opcode_2 != 4'h0 ? _GEN_4610 : _GEN_3842; // @[executor.scala 470:55]
  wire [7:0] _GEN_5379 = opcode_2 != 4'h0 ? _GEN_4611 : _GEN_3843; // @[executor.scala 470:55]
  wire [7:0] _GEN_5380 = opcode_2 != 4'h0 ? _GEN_4616 : _GEN_3844; // @[executor.scala 470:55]
  wire [7:0] _GEN_5381 = opcode_2 != 4'h0 ? _GEN_4617 : _GEN_3845; // @[executor.scala 470:55]
  wire [7:0] _GEN_5382 = opcode_2 != 4'h0 ? _GEN_4618 : _GEN_3846; // @[executor.scala 470:55]
  wire [7:0] _GEN_5383 = opcode_2 != 4'h0 ? _GEN_4619 : _GEN_3847; // @[executor.scala 470:55]
  wire [7:0] _GEN_5384 = opcode_2 != 4'h0 ? _GEN_4624 : _GEN_3848; // @[executor.scala 470:55]
  wire [7:0] _GEN_5385 = opcode_2 != 4'h0 ? _GEN_4625 : _GEN_3849; // @[executor.scala 470:55]
  wire [7:0] _GEN_5386 = opcode_2 != 4'h0 ? _GEN_4626 : _GEN_3850; // @[executor.scala 470:55]
  wire [7:0] _GEN_5387 = opcode_2 != 4'h0 ? _GEN_4627 : _GEN_3851; // @[executor.scala 470:55]
  wire [7:0] _GEN_5388 = opcode_2 != 4'h0 ? _GEN_4632 : _GEN_3852; // @[executor.scala 470:55]
  wire [7:0] _GEN_5389 = opcode_2 != 4'h0 ? _GEN_4633 : _GEN_3853; // @[executor.scala 470:55]
  wire [7:0] _GEN_5390 = opcode_2 != 4'h0 ? _GEN_4634 : _GEN_3854; // @[executor.scala 470:55]
  wire [7:0] _GEN_5391 = opcode_2 != 4'h0 ? _GEN_4635 : _GEN_3855; // @[executor.scala 470:55]
  wire [7:0] _GEN_5392 = opcode_2 != 4'h0 ? _GEN_4640 : _GEN_3856; // @[executor.scala 470:55]
  wire [7:0] _GEN_5393 = opcode_2 != 4'h0 ? _GEN_4641 : _GEN_3857; // @[executor.scala 470:55]
  wire [7:0] _GEN_5394 = opcode_2 != 4'h0 ? _GEN_4642 : _GEN_3858; // @[executor.scala 470:55]
  wire [7:0] _GEN_5395 = opcode_2 != 4'h0 ? _GEN_4643 : _GEN_3859; // @[executor.scala 470:55]
  wire [7:0] _GEN_5396 = opcode_2 != 4'h0 ? _GEN_4648 : _GEN_3860; // @[executor.scala 470:55]
  wire [7:0] _GEN_5397 = opcode_2 != 4'h0 ? _GEN_4649 : _GEN_3861; // @[executor.scala 470:55]
  wire [7:0] _GEN_5398 = opcode_2 != 4'h0 ? _GEN_4650 : _GEN_3862; // @[executor.scala 470:55]
  wire [7:0] _GEN_5399 = opcode_2 != 4'h0 ? _GEN_4651 : _GEN_3863; // @[executor.scala 470:55]
  wire [7:0] _GEN_5400 = opcode_2 != 4'h0 ? _GEN_4656 : _GEN_3864; // @[executor.scala 470:55]
  wire [7:0] _GEN_5401 = opcode_2 != 4'h0 ? _GEN_4657 : _GEN_3865; // @[executor.scala 470:55]
  wire [7:0] _GEN_5402 = opcode_2 != 4'h0 ? _GEN_4658 : _GEN_3866; // @[executor.scala 470:55]
  wire [7:0] _GEN_5403 = opcode_2 != 4'h0 ? _GEN_4659 : _GEN_3867; // @[executor.scala 470:55]
  wire [7:0] _GEN_5404 = opcode_2 != 4'h0 ? _GEN_4664 : _GEN_3868; // @[executor.scala 470:55]
  wire [7:0] _GEN_5405 = opcode_2 != 4'h0 ? _GEN_4665 : _GEN_3869; // @[executor.scala 470:55]
  wire [7:0] _GEN_5406 = opcode_2 != 4'h0 ? _GEN_4666 : _GEN_3870; // @[executor.scala 470:55]
  wire [7:0] _GEN_5407 = opcode_2 != 4'h0 ? _GEN_4667 : _GEN_3871; // @[executor.scala 470:55]
  wire [7:0] _GEN_5408 = opcode_2 != 4'h0 ? _GEN_4672 : _GEN_3872; // @[executor.scala 470:55]
  wire [7:0] _GEN_5409 = opcode_2 != 4'h0 ? _GEN_4673 : _GEN_3873; // @[executor.scala 470:55]
  wire [7:0] _GEN_5410 = opcode_2 != 4'h0 ? _GEN_4674 : _GEN_3874; // @[executor.scala 470:55]
  wire [7:0] _GEN_5411 = opcode_2 != 4'h0 ? _GEN_4675 : _GEN_3875; // @[executor.scala 470:55]
  wire [7:0] _GEN_5412 = opcode_2 != 4'h0 ? _GEN_4680 : _GEN_3876; // @[executor.scala 470:55]
  wire [7:0] _GEN_5413 = opcode_2 != 4'h0 ? _GEN_4681 : _GEN_3877; // @[executor.scala 470:55]
  wire [7:0] _GEN_5414 = opcode_2 != 4'h0 ? _GEN_4682 : _GEN_3878; // @[executor.scala 470:55]
  wire [7:0] _GEN_5415 = opcode_2 != 4'h0 ? _GEN_4683 : _GEN_3879; // @[executor.scala 470:55]
  wire [7:0] _GEN_5416 = opcode_2 != 4'h0 ? _GEN_4688 : _GEN_3880; // @[executor.scala 470:55]
  wire [7:0] _GEN_5417 = opcode_2 != 4'h0 ? _GEN_4689 : _GEN_3881; // @[executor.scala 470:55]
  wire [7:0] _GEN_5418 = opcode_2 != 4'h0 ? _GEN_4690 : _GEN_3882; // @[executor.scala 470:55]
  wire [7:0] _GEN_5419 = opcode_2 != 4'h0 ? _GEN_4691 : _GEN_3883; // @[executor.scala 470:55]
  wire [7:0] _GEN_5420 = opcode_2 != 4'h0 ? _GEN_4696 : _GEN_3884; // @[executor.scala 470:55]
  wire [7:0] _GEN_5421 = opcode_2 != 4'h0 ? _GEN_4697 : _GEN_3885; // @[executor.scala 470:55]
  wire [7:0] _GEN_5422 = opcode_2 != 4'h0 ? _GEN_4698 : _GEN_3886; // @[executor.scala 470:55]
  wire [7:0] _GEN_5423 = opcode_2 != 4'h0 ? _GEN_4699 : _GEN_3887; // @[executor.scala 470:55]
  wire [7:0] _GEN_5424 = opcode_2 != 4'h0 ? _GEN_4704 : _GEN_3888; // @[executor.scala 470:55]
  wire [7:0] _GEN_5425 = opcode_2 != 4'h0 ? _GEN_4705 : _GEN_3889; // @[executor.scala 470:55]
  wire [7:0] _GEN_5426 = opcode_2 != 4'h0 ? _GEN_4706 : _GEN_3890; // @[executor.scala 470:55]
  wire [7:0] _GEN_5427 = opcode_2 != 4'h0 ? _GEN_4707 : _GEN_3891; // @[executor.scala 470:55]
  wire [7:0] _GEN_5428 = opcode_2 != 4'h0 ? _GEN_4712 : _GEN_3892; // @[executor.scala 470:55]
  wire [7:0] _GEN_5429 = opcode_2 != 4'h0 ? _GEN_4713 : _GEN_3893; // @[executor.scala 470:55]
  wire [7:0] _GEN_5430 = opcode_2 != 4'h0 ? _GEN_4714 : _GEN_3894; // @[executor.scala 470:55]
  wire [7:0] _GEN_5431 = opcode_2 != 4'h0 ? _GEN_4715 : _GEN_3895; // @[executor.scala 470:55]
  wire [7:0] _GEN_5432 = opcode_2 != 4'h0 ? _GEN_4720 : _GEN_3896; // @[executor.scala 470:55]
  wire [7:0] _GEN_5433 = opcode_2 != 4'h0 ? _GEN_4721 : _GEN_3897; // @[executor.scala 470:55]
  wire [7:0] _GEN_5434 = opcode_2 != 4'h0 ? _GEN_4722 : _GEN_3898; // @[executor.scala 470:55]
  wire [7:0] _GEN_5435 = opcode_2 != 4'h0 ? _GEN_4723 : _GEN_3899; // @[executor.scala 470:55]
  wire [7:0] _GEN_5436 = opcode_2 != 4'h0 ? _GEN_4728 : _GEN_3900; // @[executor.scala 470:55]
  wire [7:0] _GEN_5437 = opcode_2 != 4'h0 ? _GEN_4729 : _GEN_3901; // @[executor.scala 470:55]
  wire [7:0] _GEN_5438 = opcode_2 != 4'h0 ? _GEN_4730 : _GEN_3902; // @[executor.scala 470:55]
  wire [7:0] _GEN_5439 = opcode_2 != 4'h0 ? _GEN_4731 : _GEN_3903; // @[executor.scala 470:55]
  wire [7:0] _GEN_5440 = opcode_2 != 4'h0 ? _GEN_4736 : _GEN_3904; // @[executor.scala 470:55]
  wire [7:0] _GEN_5441 = opcode_2 != 4'h0 ? _GEN_4737 : _GEN_3905; // @[executor.scala 470:55]
  wire [7:0] _GEN_5442 = opcode_2 != 4'h0 ? _GEN_4738 : _GEN_3906; // @[executor.scala 470:55]
  wire [7:0] _GEN_5443 = opcode_2 != 4'h0 ? _GEN_4739 : _GEN_3907; // @[executor.scala 470:55]
  wire [7:0] _GEN_5444 = opcode_2 != 4'h0 ? _GEN_4744 : _GEN_3908; // @[executor.scala 470:55]
  wire [7:0] _GEN_5445 = opcode_2 != 4'h0 ? _GEN_4745 : _GEN_3909; // @[executor.scala 470:55]
  wire [7:0] _GEN_5446 = opcode_2 != 4'h0 ? _GEN_4746 : _GEN_3910; // @[executor.scala 470:55]
  wire [7:0] _GEN_5447 = opcode_2 != 4'h0 ? _GEN_4747 : _GEN_3911; // @[executor.scala 470:55]
  wire [7:0] _GEN_5448 = opcode_2 != 4'h0 ? _GEN_4752 : _GEN_3912; // @[executor.scala 470:55]
  wire [7:0] _GEN_5449 = opcode_2 != 4'h0 ? _GEN_4753 : _GEN_3913; // @[executor.scala 470:55]
  wire [7:0] _GEN_5450 = opcode_2 != 4'h0 ? _GEN_4754 : _GEN_3914; // @[executor.scala 470:55]
  wire [7:0] _GEN_5451 = opcode_2 != 4'h0 ? _GEN_4755 : _GEN_3915; // @[executor.scala 470:55]
  wire [7:0] _GEN_5452 = opcode_2 != 4'h0 ? _GEN_4760 : _GEN_3916; // @[executor.scala 470:55]
  wire [7:0] _GEN_5453 = opcode_2 != 4'h0 ? _GEN_4761 : _GEN_3917; // @[executor.scala 470:55]
  wire [7:0] _GEN_5454 = opcode_2 != 4'h0 ? _GEN_4762 : _GEN_3918; // @[executor.scala 470:55]
  wire [7:0] _GEN_5455 = opcode_2 != 4'h0 ? _GEN_4763 : _GEN_3919; // @[executor.scala 470:55]
  wire [7:0] _GEN_5456 = opcode_2 != 4'h0 ? _GEN_4768 : _GEN_3920; // @[executor.scala 470:55]
  wire [7:0] _GEN_5457 = opcode_2 != 4'h0 ? _GEN_4769 : _GEN_3921; // @[executor.scala 470:55]
  wire [7:0] _GEN_5458 = opcode_2 != 4'h0 ? _GEN_4770 : _GEN_3922; // @[executor.scala 470:55]
  wire [7:0] _GEN_5459 = opcode_2 != 4'h0 ? _GEN_4771 : _GEN_3923; // @[executor.scala 470:55]
  wire [7:0] _GEN_5460 = opcode_2 != 4'h0 ? _GEN_4776 : _GEN_3924; // @[executor.scala 470:55]
  wire [7:0] _GEN_5461 = opcode_2 != 4'h0 ? _GEN_4777 : _GEN_3925; // @[executor.scala 470:55]
  wire [7:0] _GEN_5462 = opcode_2 != 4'h0 ? _GEN_4778 : _GEN_3926; // @[executor.scala 470:55]
  wire [7:0] _GEN_5463 = opcode_2 != 4'h0 ? _GEN_4779 : _GEN_3927; // @[executor.scala 470:55]
  wire [7:0] _GEN_5464 = opcode_2 != 4'h0 ? _GEN_4784 : _GEN_3928; // @[executor.scala 470:55]
  wire [7:0] _GEN_5465 = opcode_2 != 4'h0 ? _GEN_4785 : _GEN_3929; // @[executor.scala 470:55]
  wire [7:0] _GEN_5466 = opcode_2 != 4'h0 ? _GEN_4786 : _GEN_3930; // @[executor.scala 470:55]
  wire [7:0] _GEN_5467 = opcode_2 != 4'h0 ? _GEN_4787 : _GEN_3931; // @[executor.scala 470:55]
  wire [7:0] _GEN_5468 = opcode_2 != 4'h0 ? _GEN_4792 : _GEN_3932; // @[executor.scala 470:55]
  wire [7:0] _GEN_5469 = opcode_2 != 4'h0 ? _GEN_4793 : _GEN_3933; // @[executor.scala 470:55]
  wire [7:0] _GEN_5470 = opcode_2 != 4'h0 ? _GEN_4794 : _GEN_3934; // @[executor.scala 470:55]
  wire [7:0] _GEN_5471 = opcode_2 != 4'h0 ? _GEN_4795 : _GEN_3935; // @[executor.scala 470:55]
  wire [7:0] _GEN_5472 = opcode_2 != 4'h0 ? _GEN_4800 : _GEN_3936; // @[executor.scala 470:55]
  wire [7:0] _GEN_5473 = opcode_2 != 4'h0 ? _GEN_4801 : _GEN_3937; // @[executor.scala 470:55]
  wire [7:0] _GEN_5474 = opcode_2 != 4'h0 ? _GEN_4802 : _GEN_3938; // @[executor.scala 470:55]
  wire [7:0] _GEN_5475 = opcode_2 != 4'h0 ? _GEN_4803 : _GEN_3939; // @[executor.scala 470:55]
  wire [7:0] _GEN_5476 = opcode_2 != 4'h0 ? _GEN_4808 : _GEN_3940; // @[executor.scala 470:55]
  wire [7:0] _GEN_5477 = opcode_2 != 4'h0 ? _GEN_4809 : _GEN_3941; // @[executor.scala 470:55]
  wire [7:0] _GEN_5478 = opcode_2 != 4'h0 ? _GEN_4810 : _GEN_3942; // @[executor.scala 470:55]
  wire [7:0] _GEN_5479 = opcode_2 != 4'h0 ? _GEN_4811 : _GEN_3943; // @[executor.scala 470:55]
  wire [7:0] _GEN_5480 = opcode_2 != 4'h0 ? _GEN_4816 : _GEN_3944; // @[executor.scala 470:55]
  wire [7:0] _GEN_5481 = opcode_2 != 4'h0 ? _GEN_4817 : _GEN_3945; // @[executor.scala 470:55]
  wire [7:0] _GEN_5482 = opcode_2 != 4'h0 ? _GEN_4818 : _GEN_3946; // @[executor.scala 470:55]
  wire [7:0] _GEN_5483 = opcode_2 != 4'h0 ? _GEN_4819 : _GEN_3947; // @[executor.scala 470:55]
  wire [7:0] _GEN_5484 = opcode_2 != 4'h0 ? _GEN_4824 : _GEN_3948; // @[executor.scala 470:55]
  wire [7:0] _GEN_5485 = opcode_2 != 4'h0 ? _GEN_4825 : _GEN_3949; // @[executor.scala 470:55]
  wire [7:0] _GEN_5486 = opcode_2 != 4'h0 ? _GEN_4826 : _GEN_3950; // @[executor.scala 470:55]
  wire [7:0] _GEN_5487 = opcode_2 != 4'h0 ? _GEN_4827 : _GEN_3951; // @[executor.scala 470:55]
  wire [7:0] _GEN_5488 = opcode_2 != 4'h0 ? _GEN_4832 : _GEN_3952; // @[executor.scala 470:55]
  wire [7:0] _GEN_5489 = opcode_2 != 4'h0 ? _GEN_4833 : _GEN_3953; // @[executor.scala 470:55]
  wire [7:0] _GEN_5490 = opcode_2 != 4'h0 ? _GEN_4834 : _GEN_3954; // @[executor.scala 470:55]
  wire [7:0] _GEN_5491 = opcode_2 != 4'h0 ? _GEN_4835 : _GEN_3955; // @[executor.scala 470:55]
  wire [7:0] _GEN_5492 = opcode_2 != 4'h0 ? _GEN_4840 : _GEN_3956; // @[executor.scala 470:55]
  wire [7:0] _GEN_5493 = opcode_2 != 4'h0 ? _GEN_4841 : _GEN_3957; // @[executor.scala 470:55]
  wire [7:0] _GEN_5494 = opcode_2 != 4'h0 ? _GEN_4842 : _GEN_3958; // @[executor.scala 470:55]
  wire [7:0] _GEN_5495 = opcode_2 != 4'h0 ? _GEN_4843 : _GEN_3959; // @[executor.scala 470:55]
  wire [7:0] _GEN_5496 = opcode_2 != 4'h0 ? _GEN_4848 : _GEN_3960; // @[executor.scala 470:55]
  wire [7:0] _GEN_5497 = opcode_2 != 4'h0 ? _GEN_4849 : _GEN_3961; // @[executor.scala 470:55]
  wire [7:0] _GEN_5498 = opcode_2 != 4'h0 ? _GEN_4850 : _GEN_3962; // @[executor.scala 470:55]
  wire [7:0] _GEN_5499 = opcode_2 != 4'h0 ? _GEN_4851 : _GEN_3963; // @[executor.scala 470:55]
  wire [7:0] _GEN_5500 = opcode_2 != 4'h0 ? _GEN_4856 : _GEN_3964; // @[executor.scala 470:55]
  wire [7:0] _GEN_5501 = opcode_2 != 4'h0 ? _GEN_4857 : _GEN_3965; // @[executor.scala 470:55]
  wire [7:0] _GEN_5502 = opcode_2 != 4'h0 ? _GEN_4858 : _GEN_3966; // @[executor.scala 470:55]
  wire [7:0] _GEN_5503 = opcode_2 != 4'h0 ? _GEN_4859 : _GEN_3967; // @[executor.scala 470:55]
  wire [7:0] _GEN_5504 = opcode_2 != 4'h0 ? _GEN_4864 : _GEN_3968; // @[executor.scala 470:55]
  wire [7:0] _GEN_5505 = opcode_2 != 4'h0 ? _GEN_4865 : _GEN_3969; // @[executor.scala 470:55]
  wire [7:0] _GEN_5506 = opcode_2 != 4'h0 ? _GEN_4866 : _GEN_3970; // @[executor.scala 470:55]
  wire [7:0] _GEN_5507 = opcode_2 != 4'h0 ? _GEN_4867 : _GEN_3971; // @[executor.scala 470:55]
  wire [7:0] _GEN_5508 = opcode_2 != 4'h0 ? _GEN_4872 : _GEN_3972; // @[executor.scala 470:55]
  wire [7:0] _GEN_5509 = opcode_2 != 4'h0 ? _GEN_4873 : _GEN_3973; // @[executor.scala 470:55]
  wire [7:0] _GEN_5510 = opcode_2 != 4'h0 ? _GEN_4874 : _GEN_3974; // @[executor.scala 470:55]
  wire [7:0] _GEN_5511 = opcode_2 != 4'h0 ? _GEN_4875 : _GEN_3975; // @[executor.scala 470:55]
  wire [7:0] _GEN_5512 = opcode_2 != 4'h0 ? _GEN_4880 : _GEN_3976; // @[executor.scala 470:55]
  wire [7:0] _GEN_5513 = opcode_2 != 4'h0 ? _GEN_4881 : _GEN_3977; // @[executor.scala 470:55]
  wire [7:0] _GEN_5514 = opcode_2 != 4'h0 ? _GEN_4882 : _GEN_3978; // @[executor.scala 470:55]
  wire [7:0] _GEN_5515 = opcode_2 != 4'h0 ? _GEN_4883 : _GEN_3979; // @[executor.scala 470:55]
  wire [7:0] _GEN_5516 = opcode_2 != 4'h0 ? _GEN_4888 : _GEN_3980; // @[executor.scala 470:55]
  wire [7:0] _GEN_5517 = opcode_2 != 4'h0 ? _GEN_4889 : _GEN_3981; // @[executor.scala 470:55]
  wire [7:0] _GEN_5518 = opcode_2 != 4'h0 ? _GEN_4890 : _GEN_3982; // @[executor.scala 470:55]
  wire [7:0] _GEN_5519 = opcode_2 != 4'h0 ? _GEN_4891 : _GEN_3983; // @[executor.scala 470:55]
  wire [7:0] _GEN_5520 = opcode_2 != 4'h0 ? _GEN_4896 : _GEN_3984; // @[executor.scala 470:55]
  wire [7:0] _GEN_5521 = opcode_2 != 4'h0 ? _GEN_4897 : _GEN_3985; // @[executor.scala 470:55]
  wire [7:0] _GEN_5522 = opcode_2 != 4'h0 ? _GEN_4898 : _GEN_3986; // @[executor.scala 470:55]
  wire [7:0] _GEN_5523 = opcode_2 != 4'h0 ? _GEN_4899 : _GEN_3987; // @[executor.scala 470:55]
  wire [7:0] _GEN_5524 = opcode_2 != 4'h0 ? _GEN_4904 : _GEN_3988; // @[executor.scala 470:55]
  wire [7:0] _GEN_5525 = opcode_2 != 4'h0 ? _GEN_4905 : _GEN_3989; // @[executor.scala 470:55]
  wire [7:0] _GEN_5526 = opcode_2 != 4'h0 ? _GEN_4906 : _GEN_3990; // @[executor.scala 470:55]
  wire [7:0] _GEN_5527 = opcode_2 != 4'h0 ? _GEN_4907 : _GEN_3991; // @[executor.scala 470:55]
  wire [7:0] _GEN_5528 = opcode_2 != 4'h0 ? _GEN_4912 : _GEN_3992; // @[executor.scala 470:55]
  wire [7:0] _GEN_5529 = opcode_2 != 4'h0 ? _GEN_4913 : _GEN_3993; // @[executor.scala 470:55]
  wire [7:0] _GEN_5530 = opcode_2 != 4'h0 ? _GEN_4914 : _GEN_3994; // @[executor.scala 470:55]
  wire [7:0] _GEN_5531 = opcode_2 != 4'h0 ? _GEN_4915 : _GEN_3995; // @[executor.scala 470:55]
  wire [7:0] _GEN_5532 = opcode_2 != 4'h0 ? _GEN_4920 : _GEN_3996; // @[executor.scala 470:55]
  wire [7:0] _GEN_5533 = opcode_2 != 4'h0 ? _GEN_4921 : _GEN_3997; // @[executor.scala 470:55]
  wire [7:0] _GEN_5534 = opcode_2 != 4'h0 ? _GEN_4922 : _GEN_3998; // @[executor.scala 470:55]
  wire [7:0] _GEN_5535 = opcode_2 != 4'h0 ? _GEN_4923 : _GEN_3999; // @[executor.scala 470:55]
  wire [7:0] _GEN_5536 = opcode_2 != 4'h0 ? _GEN_4928 : _GEN_4000; // @[executor.scala 470:55]
  wire [7:0] _GEN_5537 = opcode_2 != 4'h0 ? _GEN_4929 : _GEN_4001; // @[executor.scala 470:55]
  wire [7:0] _GEN_5538 = opcode_2 != 4'h0 ? _GEN_4930 : _GEN_4002; // @[executor.scala 470:55]
  wire [7:0] _GEN_5539 = opcode_2 != 4'h0 ? _GEN_4931 : _GEN_4003; // @[executor.scala 470:55]
  wire [7:0] _GEN_5540 = opcode_2 != 4'h0 ? _GEN_4936 : _GEN_4004; // @[executor.scala 470:55]
  wire [7:0] _GEN_5541 = opcode_2 != 4'h0 ? _GEN_4937 : _GEN_4005; // @[executor.scala 470:55]
  wire [7:0] _GEN_5542 = opcode_2 != 4'h0 ? _GEN_4938 : _GEN_4006; // @[executor.scala 470:55]
  wire [7:0] _GEN_5543 = opcode_2 != 4'h0 ? _GEN_4939 : _GEN_4007; // @[executor.scala 470:55]
  wire [7:0] _GEN_5544 = opcode_2 != 4'h0 ? _GEN_4944 : _GEN_4008; // @[executor.scala 470:55]
  wire [7:0] _GEN_5545 = opcode_2 != 4'h0 ? _GEN_4945 : _GEN_4009; // @[executor.scala 470:55]
  wire [7:0] _GEN_5546 = opcode_2 != 4'h0 ? _GEN_4946 : _GEN_4010; // @[executor.scala 470:55]
  wire [7:0] _GEN_5547 = opcode_2 != 4'h0 ? _GEN_4947 : _GEN_4011; // @[executor.scala 470:55]
  wire [7:0] _GEN_5548 = opcode_2 != 4'h0 ? _GEN_4952 : _GEN_4012; // @[executor.scala 470:55]
  wire [7:0] _GEN_5549 = opcode_2 != 4'h0 ? _GEN_4953 : _GEN_4013; // @[executor.scala 470:55]
  wire [7:0] _GEN_5550 = opcode_2 != 4'h0 ? _GEN_4954 : _GEN_4014; // @[executor.scala 470:55]
  wire [7:0] _GEN_5551 = opcode_2 != 4'h0 ? _GEN_4955 : _GEN_4015; // @[executor.scala 470:55]
  wire [7:0] _GEN_5552 = opcode_2 != 4'h0 ? _GEN_4960 : _GEN_4016; // @[executor.scala 470:55]
  wire [7:0] _GEN_5553 = opcode_2 != 4'h0 ? _GEN_4961 : _GEN_4017; // @[executor.scala 470:55]
  wire [7:0] _GEN_5554 = opcode_2 != 4'h0 ? _GEN_4962 : _GEN_4018; // @[executor.scala 470:55]
  wire [7:0] _GEN_5555 = opcode_2 != 4'h0 ? _GEN_4963 : _GEN_4019; // @[executor.scala 470:55]
  wire [7:0] _GEN_5556 = opcode_2 != 4'h0 ? _GEN_4968 : _GEN_4020; // @[executor.scala 470:55]
  wire [7:0] _GEN_5557 = opcode_2 != 4'h0 ? _GEN_4969 : _GEN_4021; // @[executor.scala 470:55]
  wire [7:0] _GEN_5558 = opcode_2 != 4'h0 ? _GEN_4970 : _GEN_4022; // @[executor.scala 470:55]
  wire [7:0] _GEN_5559 = opcode_2 != 4'h0 ? _GEN_4971 : _GEN_4023; // @[executor.scala 470:55]
  wire [7:0] _GEN_5560 = opcode_2 != 4'h0 ? _GEN_4976 : _GEN_4024; // @[executor.scala 470:55]
  wire [7:0] _GEN_5561 = opcode_2 != 4'h0 ? _GEN_4977 : _GEN_4025; // @[executor.scala 470:55]
  wire [7:0] _GEN_5562 = opcode_2 != 4'h0 ? _GEN_4978 : _GEN_4026; // @[executor.scala 470:55]
  wire [7:0] _GEN_5563 = opcode_2 != 4'h0 ? _GEN_4979 : _GEN_4027; // @[executor.scala 470:55]
  wire [7:0] _GEN_5564 = opcode_2 != 4'h0 ? _GEN_4984 : _GEN_4028; // @[executor.scala 470:55]
  wire [7:0] _GEN_5565 = opcode_2 != 4'h0 ? _GEN_4985 : _GEN_4029; // @[executor.scala 470:55]
  wire [7:0] _GEN_5566 = opcode_2 != 4'h0 ? _GEN_4986 : _GEN_4030; // @[executor.scala 470:55]
  wire [7:0] _GEN_5567 = opcode_2 != 4'h0 ? _GEN_4987 : _GEN_4031; // @[executor.scala 470:55]
  wire [7:0] _GEN_5568 = opcode_2 != 4'h0 ? _GEN_4992 : _GEN_4032; // @[executor.scala 470:55]
  wire [7:0] _GEN_5569 = opcode_2 != 4'h0 ? _GEN_4993 : _GEN_4033; // @[executor.scala 470:55]
  wire [7:0] _GEN_5570 = opcode_2 != 4'h0 ? _GEN_4994 : _GEN_4034; // @[executor.scala 470:55]
  wire [7:0] _GEN_5571 = opcode_2 != 4'h0 ? _GEN_4995 : _GEN_4035; // @[executor.scala 470:55]
  wire [7:0] _GEN_5572 = opcode_2 != 4'h0 ? _GEN_5000 : _GEN_4036; // @[executor.scala 470:55]
  wire [7:0] _GEN_5573 = opcode_2 != 4'h0 ? _GEN_5001 : _GEN_4037; // @[executor.scala 470:55]
  wire [7:0] _GEN_5574 = opcode_2 != 4'h0 ? _GEN_5002 : _GEN_4038; // @[executor.scala 470:55]
  wire [7:0] _GEN_5575 = opcode_2 != 4'h0 ? _GEN_5003 : _GEN_4039; // @[executor.scala 470:55]
  wire [7:0] _GEN_5576 = opcode_2 != 4'h0 ? _GEN_5008 : _GEN_4040; // @[executor.scala 470:55]
  wire [7:0] _GEN_5577 = opcode_2 != 4'h0 ? _GEN_5009 : _GEN_4041; // @[executor.scala 470:55]
  wire [7:0] _GEN_5578 = opcode_2 != 4'h0 ? _GEN_5010 : _GEN_4042; // @[executor.scala 470:55]
  wire [7:0] _GEN_5579 = opcode_2 != 4'h0 ? _GEN_5011 : _GEN_4043; // @[executor.scala 470:55]
  wire [7:0] _GEN_5580 = opcode_2 != 4'h0 ? _GEN_5016 : _GEN_4044; // @[executor.scala 470:55]
  wire [7:0] _GEN_5581 = opcode_2 != 4'h0 ? _GEN_5017 : _GEN_4045; // @[executor.scala 470:55]
  wire [7:0] _GEN_5582 = opcode_2 != 4'h0 ? _GEN_5018 : _GEN_4046; // @[executor.scala 470:55]
  wire [7:0] _GEN_5583 = opcode_2 != 4'h0 ? _GEN_5019 : _GEN_4047; // @[executor.scala 470:55]
  wire [7:0] _GEN_5584 = opcode_2 != 4'h0 ? _GEN_5024 : _GEN_4048; // @[executor.scala 470:55]
  wire [7:0] _GEN_5585 = opcode_2 != 4'h0 ? _GEN_5025 : _GEN_4049; // @[executor.scala 470:55]
  wire [7:0] _GEN_5586 = opcode_2 != 4'h0 ? _GEN_5026 : _GEN_4050; // @[executor.scala 470:55]
  wire [7:0] _GEN_5587 = opcode_2 != 4'h0 ? _GEN_5027 : _GEN_4051; // @[executor.scala 470:55]
  wire [7:0] _GEN_5588 = opcode_2 != 4'h0 ? _GEN_5032 : _GEN_4052; // @[executor.scala 470:55]
  wire [7:0] _GEN_5589 = opcode_2 != 4'h0 ? _GEN_5033 : _GEN_4053; // @[executor.scala 470:55]
  wire [7:0] _GEN_5590 = opcode_2 != 4'h0 ? _GEN_5034 : _GEN_4054; // @[executor.scala 470:55]
  wire [7:0] _GEN_5591 = opcode_2 != 4'h0 ? _GEN_5035 : _GEN_4055; // @[executor.scala 470:55]
  wire [7:0] _GEN_5592 = opcode_2 != 4'h0 ? _GEN_5040 : _GEN_4056; // @[executor.scala 470:55]
  wire [7:0] _GEN_5593 = opcode_2 != 4'h0 ? _GEN_5041 : _GEN_4057; // @[executor.scala 470:55]
  wire [7:0] _GEN_5594 = opcode_2 != 4'h0 ? _GEN_5042 : _GEN_4058; // @[executor.scala 470:55]
  wire [7:0] _GEN_5595 = opcode_2 != 4'h0 ? _GEN_5043 : _GEN_4059; // @[executor.scala 470:55]
  wire [7:0] _GEN_5596 = opcode_2 != 4'h0 ? _GEN_5048 : _GEN_4060; // @[executor.scala 470:55]
  wire [7:0] _GEN_5597 = opcode_2 != 4'h0 ? _GEN_5049 : _GEN_4061; // @[executor.scala 470:55]
  wire [7:0] _GEN_5598 = opcode_2 != 4'h0 ? _GEN_5050 : _GEN_4062; // @[executor.scala 470:55]
  wire [7:0] _GEN_5599 = opcode_2 != 4'h0 ? _GEN_5051 : _GEN_4063; // @[executor.scala 470:55]
  wire [7:0] _GEN_5600 = opcode_2 != 4'h0 ? _GEN_5056 : _GEN_4064; // @[executor.scala 470:55]
  wire [7:0] _GEN_5601 = opcode_2 != 4'h0 ? _GEN_5057 : _GEN_4065; // @[executor.scala 470:55]
  wire [7:0] _GEN_5602 = opcode_2 != 4'h0 ? _GEN_5058 : _GEN_4066; // @[executor.scala 470:55]
  wire [7:0] _GEN_5603 = opcode_2 != 4'h0 ? _GEN_5059 : _GEN_4067; // @[executor.scala 470:55]
  wire [7:0] _GEN_5604 = opcode_2 != 4'h0 ? _GEN_5064 : _GEN_4068; // @[executor.scala 470:55]
  wire [7:0] _GEN_5605 = opcode_2 != 4'h0 ? _GEN_5065 : _GEN_4069; // @[executor.scala 470:55]
  wire [7:0] _GEN_5606 = opcode_2 != 4'h0 ? _GEN_5066 : _GEN_4070; // @[executor.scala 470:55]
  wire [7:0] _GEN_5607 = opcode_2 != 4'h0 ? _GEN_5067 : _GEN_4071; // @[executor.scala 470:55]
  wire [7:0] _GEN_5608 = opcode_2 != 4'h0 ? _GEN_5072 : _GEN_4072; // @[executor.scala 470:55]
  wire [7:0] _GEN_5609 = opcode_2 != 4'h0 ? _GEN_5073 : _GEN_4073; // @[executor.scala 470:55]
  wire [7:0] _GEN_5610 = opcode_2 != 4'h0 ? _GEN_5074 : _GEN_4074; // @[executor.scala 470:55]
  wire [7:0] _GEN_5611 = opcode_2 != 4'h0 ? _GEN_5075 : _GEN_4075; // @[executor.scala 470:55]
  wire [7:0] _GEN_5612 = opcode_2 != 4'h0 ? _GEN_5080 : _GEN_4076; // @[executor.scala 470:55]
  wire [7:0] _GEN_5613 = opcode_2 != 4'h0 ? _GEN_5081 : _GEN_4077; // @[executor.scala 470:55]
  wire [7:0] _GEN_5614 = opcode_2 != 4'h0 ? _GEN_5082 : _GEN_4078; // @[executor.scala 470:55]
  wire [7:0] _GEN_5615 = opcode_2 != 4'h0 ? _GEN_5083 : _GEN_4079; // @[executor.scala 470:55]
  wire [7:0] _GEN_5616 = opcode_2 != 4'h0 ? _GEN_5088 : _GEN_4080; // @[executor.scala 470:55]
  wire [7:0] _GEN_5617 = opcode_2 != 4'h0 ? _GEN_5089 : _GEN_4081; // @[executor.scala 470:55]
  wire [7:0] _GEN_5618 = opcode_2 != 4'h0 ? _GEN_5090 : _GEN_4082; // @[executor.scala 470:55]
  wire [7:0] _GEN_5619 = opcode_2 != 4'h0 ? _GEN_5091 : _GEN_4083; // @[executor.scala 470:55]
  wire [7:0] _GEN_5620 = opcode_2 != 4'h0 ? _GEN_5096 : _GEN_4084; // @[executor.scala 470:55]
  wire [7:0] _GEN_5621 = opcode_2 != 4'h0 ? _GEN_5097 : _GEN_4085; // @[executor.scala 470:55]
  wire [7:0] _GEN_5622 = opcode_2 != 4'h0 ? _GEN_5098 : _GEN_4086; // @[executor.scala 470:55]
  wire [7:0] _GEN_5623 = opcode_2 != 4'h0 ? _GEN_5099 : _GEN_4087; // @[executor.scala 470:55]
  wire [7:0] _GEN_5624 = opcode_2 != 4'h0 ? _GEN_5104 : _GEN_4088; // @[executor.scala 470:55]
  wire [7:0] _GEN_5625 = opcode_2 != 4'h0 ? _GEN_5105 : _GEN_4089; // @[executor.scala 470:55]
  wire [7:0] _GEN_5626 = opcode_2 != 4'h0 ? _GEN_5106 : _GEN_4090; // @[executor.scala 470:55]
  wire [7:0] _GEN_5627 = opcode_2 != 4'h0 ? _GEN_5107 : _GEN_4091; // @[executor.scala 470:55]
  wire [7:0] _GEN_5628 = opcode_2 != 4'h0 ? _GEN_5112 : _GEN_4092; // @[executor.scala 470:55]
  wire [7:0] _GEN_5629 = opcode_2 != 4'h0 ? _GEN_5113 : _GEN_4093; // @[executor.scala 470:55]
  wire [7:0] _GEN_5630 = opcode_2 != 4'h0 ? _GEN_5114 : _GEN_4094; // @[executor.scala 470:55]
  wire [7:0] _GEN_5631 = opcode_2 != 4'h0 ? _GEN_5115 : _GEN_4095; // @[executor.scala 470:55]
  wire [7:0] _GEN_5632 = opcode_2 != 4'h0 ? _GEN_5120 : _GEN_4096; // @[executor.scala 470:55]
  wire [7:0] _GEN_5633 = opcode_2 != 4'h0 ? _GEN_5121 : _GEN_4097; // @[executor.scala 470:55]
  wire [7:0] _GEN_5634 = opcode_2 != 4'h0 ? _GEN_5122 : _GEN_4098; // @[executor.scala 470:55]
  wire [7:0] _GEN_5635 = opcode_2 != 4'h0 ? _GEN_5123 : _GEN_4099; // @[executor.scala 470:55]
  wire [3:0] _GEN_5636 = opcode_2 == 4'hf ? parameter_2_2[13:10] : _GEN_3586; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_5637 = opcode_2 == 4'hf ? parameter_2_2[0] : _GEN_3587; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_5638 = opcode_2 == 4'hf ? _GEN_3588 : _GEN_5124; // @[executor.scala 466:52]
  wire [7:0] _GEN_5639 = opcode_2 == 4'hf ? _GEN_3589 : _GEN_5125; // @[executor.scala 466:52]
  wire [7:0] _GEN_5640 = opcode_2 == 4'hf ? _GEN_3590 : _GEN_5126; // @[executor.scala 466:52]
  wire [7:0] _GEN_5641 = opcode_2 == 4'hf ? _GEN_3591 : _GEN_5127; // @[executor.scala 466:52]
  wire [7:0] _GEN_5642 = opcode_2 == 4'hf ? _GEN_3592 : _GEN_5128; // @[executor.scala 466:52]
  wire [7:0] _GEN_5643 = opcode_2 == 4'hf ? _GEN_3593 : _GEN_5129; // @[executor.scala 466:52]
  wire [7:0] _GEN_5644 = opcode_2 == 4'hf ? _GEN_3594 : _GEN_5130; // @[executor.scala 466:52]
  wire [7:0] _GEN_5645 = opcode_2 == 4'hf ? _GEN_3595 : _GEN_5131; // @[executor.scala 466:52]
  wire [7:0] _GEN_5646 = opcode_2 == 4'hf ? _GEN_3596 : _GEN_5132; // @[executor.scala 466:52]
  wire [7:0] _GEN_5647 = opcode_2 == 4'hf ? _GEN_3597 : _GEN_5133; // @[executor.scala 466:52]
  wire [7:0] _GEN_5648 = opcode_2 == 4'hf ? _GEN_3598 : _GEN_5134; // @[executor.scala 466:52]
  wire [7:0] _GEN_5649 = opcode_2 == 4'hf ? _GEN_3599 : _GEN_5135; // @[executor.scala 466:52]
  wire [7:0] _GEN_5650 = opcode_2 == 4'hf ? _GEN_3600 : _GEN_5136; // @[executor.scala 466:52]
  wire [7:0] _GEN_5651 = opcode_2 == 4'hf ? _GEN_3601 : _GEN_5137; // @[executor.scala 466:52]
  wire [7:0] _GEN_5652 = opcode_2 == 4'hf ? _GEN_3602 : _GEN_5138; // @[executor.scala 466:52]
  wire [7:0] _GEN_5653 = opcode_2 == 4'hf ? _GEN_3603 : _GEN_5139; // @[executor.scala 466:52]
  wire [7:0] _GEN_5654 = opcode_2 == 4'hf ? _GEN_3604 : _GEN_5140; // @[executor.scala 466:52]
  wire [7:0] _GEN_5655 = opcode_2 == 4'hf ? _GEN_3605 : _GEN_5141; // @[executor.scala 466:52]
  wire [7:0] _GEN_5656 = opcode_2 == 4'hf ? _GEN_3606 : _GEN_5142; // @[executor.scala 466:52]
  wire [7:0] _GEN_5657 = opcode_2 == 4'hf ? _GEN_3607 : _GEN_5143; // @[executor.scala 466:52]
  wire [7:0] _GEN_5658 = opcode_2 == 4'hf ? _GEN_3608 : _GEN_5144; // @[executor.scala 466:52]
  wire [7:0] _GEN_5659 = opcode_2 == 4'hf ? _GEN_3609 : _GEN_5145; // @[executor.scala 466:52]
  wire [7:0] _GEN_5660 = opcode_2 == 4'hf ? _GEN_3610 : _GEN_5146; // @[executor.scala 466:52]
  wire [7:0] _GEN_5661 = opcode_2 == 4'hf ? _GEN_3611 : _GEN_5147; // @[executor.scala 466:52]
  wire [7:0] _GEN_5662 = opcode_2 == 4'hf ? _GEN_3612 : _GEN_5148; // @[executor.scala 466:52]
  wire [7:0] _GEN_5663 = opcode_2 == 4'hf ? _GEN_3613 : _GEN_5149; // @[executor.scala 466:52]
  wire [7:0] _GEN_5664 = opcode_2 == 4'hf ? _GEN_3614 : _GEN_5150; // @[executor.scala 466:52]
  wire [7:0] _GEN_5665 = opcode_2 == 4'hf ? _GEN_3615 : _GEN_5151; // @[executor.scala 466:52]
  wire [7:0] _GEN_5666 = opcode_2 == 4'hf ? _GEN_3616 : _GEN_5152; // @[executor.scala 466:52]
  wire [7:0] _GEN_5667 = opcode_2 == 4'hf ? _GEN_3617 : _GEN_5153; // @[executor.scala 466:52]
  wire [7:0] _GEN_5668 = opcode_2 == 4'hf ? _GEN_3618 : _GEN_5154; // @[executor.scala 466:52]
  wire [7:0] _GEN_5669 = opcode_2 == 4'hf ? _GEN_3619 : _GEN_5155; // @[executor.scala 466:52]
  wire [7:0] _GEN_5670 = opcode_2 == 4'hf ? _GEN_3620 : _GEN_5156; // @[executor.scala 466:52]
  wire [7:0] _GEN_5671 = opcode_2 == 4'hf ? _GEN_3621 : _GEN_5157; // @[executor.scala 466:52]
  wire [7:0] _GEN_5672 = opcode_2 == 4'hf ? _GEN_3622 : _GEN_5158; // @[executor.scala 466:52]
  wire [7:0] _GEN_5673 = opcode_2 == 4'hf ? _GEN_3623 : _GEN_5159; // @[executor.scala 466:52]
  wire [7:0] _GEN_5674 = opcode_2 == 4'hf ? _GEN_3624 : _GEN_5160; // @[executor.scala 466:52]
  wire [7:0] _GEN_5675 = opcode_2 == 4'hf ? _GEN_3625 : _GEN_5161; // @[executor.scala 466:52]
  wire [7:0] _GEN_5676 = opcode_2 == 4'hf ? _GEN_3626 : _GEN_5162; // @[executor.scala 466:52]
  wire [7:0] _GEN_5677 = opcode_2 == 4'hf ? _GEN_3627 : _GEN_5163; // @[executor.scala 466:52]
  wire [7:0] _GEN_5678 = opcode_2 == 4'hf ? _GEN_3628 : _GEN_5164; // @[executor.scala 466:52]
  wire [7:0] _GEN_5679 = opcode_2 == 4'hf ? _GEN_3629 : _GEN_5165; // @[executor.scala 466:52]
  wire [7:0] _GEN_5680 = opcode_2 == 4'hf ? _GEN_3630 : _GEN_5166; // @[executor.scala 466:52]
  wire [7:0] _GEN_5681 = opcode_2 == 4'hf ? _GEN_3631 : _GEN_5167; // @[executor.scala 466:52]
  wire [7:0] _GEN_5682 = opcode_2 == 4'hf ? _GEN_3632 : _GEN_5168; // @[executor.scala 466:52]
  wire [7:0] _GEN_5683 = opcode_2 == 4'hf ? _GEN_3633 : _GEN_5169; // @[executor.scala 466:52]
  wire [7:0] _GEN_5684 = opcode_2 == 4'hf ? _GEN_3634 : _GEN_5170; // @[executor.scala 466:52]
  wire [7:0] _GEN_5685 = opcode_2 == 4'hf ? _GEN_3635 : _GEN_5171; // @[executor.scala 466:52]
  wire [7:0] _GEN_5686 = opcode_2 == 4'hf ? _GEN_3636 : _GEN_5172; // @[executor.scala 466:52]
  wire [7:0] _GEN_5687 = opcode_2 == 4'hf ? _GEN_3637 : _GEN_5173; // @[executor.scala 466:52]
  wire [7:0] _GEN_5688 = opcode_2 == 4'hf ? _GEN_3638 : _GEN_5174; // @[executor.scala 466:52]
  wire [7:0] _GEN_5689 = opcode_2 == 4'hf ? _GEN_3639 : _GEN_5175; // @[executor.scala 466:52]
  wire [7:0] _GEN_5690 = opcode_2 == 4'hf ? _GEN_3640 : _GEN_5176; // @[executor.scala 466:52]
  wire [7:0] _GEN_5691 = opcode_2 == 4'hf ? _GEN_3641 : _GEN_5177; // @[executor.scala 466:52]
  wire [7:0] _GEN_5692 = opcode_2 == 4'hf ? _GEN_3642 : _GEN_5178; // @[executor.scala 466:52]
  wire [7:0] _GEN_5693 = opcode_2 == 4'hf ? _GEN_3643 : _GEN_5179; // @[executor.scala 466:52]
  wire [7:0] _GEN_5694 = opcode_2 == 4'hf ? _GEN_3644 : _GEN_5180; // @[executor.scala 466:52]
  wire [7:0] _GEN_5695 = opcode_2 == 4'hf ? _GEN_3645 : _GEN_5181; // @[executor.scala 466:52]
  wire [7:0] _GEN_5696 = opcode_2 == 4'hf ? _GEN_3646 : _GEN_5182; // @[executor.scala 466:52]
  wire [7:0] _GEN_5697 = opcode_2 == 4'hf ? _GEN_3647 : _GEN_5183; // @[executor.scala 466:52]
  wire [7:0] _GEN_5698 = opcode_2 == 4'hf ? _GEN_3648 : _GEN_5184; // @[executor.scala 466:52]
  wire [7:0] _GEN_5699 = opcode_2 == 4'hf ? _GEN_3649 : _GEN_5185; // @[executor.scala 466:52]
  wire [7:0] _GEN_5700 = opcode_2 == 4'hf ? _GEN_3650 : _GEN_5186; // @[executor.scala 466:52]
  wire [7:0] _GEN_5701 = opcode_2 == 4'hf ? _GEN_3651 : _GEN_5187; // @[executor.scala 466:52]
  wire [7:0] _GEN_5702 = opcode_2 == 4'hf ? _GEN_3652 : _GEN_5188; // @[executor.scala 466:52]
  wire [7:0] _GEN_5703 = opcode_2 == 4'hf ? _GEN_3653 : _GEN_5189; // @[executor.scala 466:52]
  wire [7:0] _GEN_5704 = opcode_2 == 4'hf ? _GEN_3654 : _GEN_5190; // @[executor.scala 466:52]
  wire [7:0] _GEN_5705 = opcode_2 == 4'hf ? _GEN_3655 : _GEN_5191; // @[executor.scala 466:52]
  wire [7:0] _GEN_5706 = opcode_2 == 4'hf ? _GEN_3656 : _GEN_5192; // @[executor.scala 466:52]
  wire [7:0] _GEN_5707 = opcode_2 == 4'hf ? _GEN_3657 : _GEN_5193; // @[executor.scala 466:52]
  wire [7:0] _GEN_5708 = opcode_2 == 4'hf ? _GEN_3658 : _GEN_5194; // @[executor.scala 466:52]
  wire [7:0] _GEN_5709 = opcode_2 == 4'hf ? _GEN_3659 : _GEN_5195; // @[executor.scala 466:52]
  wire [7:0] _GEN_5710 = opcode_2 == 4'hf ? _GEN_3660 : _GEN_5196; // @[executor.scala 466:52]
  wire [7:0] _GEN_5711 = opcode_2 == 4'hf ? _GEN_3661 : _GEN_5197; // @[executor.scala 466:52]
  wire [7:0] _GEN_5712 = opcode_2 == 4'hf ? _GEN_3662 : _GEN_5198; // @[executor.scala 466:52]
  wire [7:0] _GEN_5713 = opcode_2 == 4'hf ? _GEN_3663 : _GEN_5199; // @[executor.scala 466:52]
  wire [7:0] _GEN_5714 = opcode_2 == 4'hf ? _GEN_3664 : _GEN_5200; // @[executor.scala 466:52]
  wire [7:0] _GEN_5715 = opcode_2 == 4'hf ? _GEN_3665 : _GEN_5201; // @[executor.scala 466:52]
  wire [7:0] _GEN_5716 = opcode_2 == 4'hf ? _GEN_3666 : _GEN_5202; // @[executor.scala 466:52]
  wire [7:0] _GEN_5717 = opcode_2 == 4'hf ? _GEN_3667 : _GEN_5203; // @[executor.scala 466:52]
  wire [7:0] _GEN_5718 = opcode_2 == 4'hf ? _GEN_3668 : _GEN_5204; // @[executor.scala 466:52]
  wire [7:0] _GEN_5719 = opcode_2 == 4'hf ? _GEN_3669 : _GEN_5205; // @[executor.scala 466:52]
  wire [7:0] _GEN_5720 = opcode_2 == 4'hf ? _GEN_3670 : _GEN_5206; // @[executor.scala 466:52]
  wire [7:0] _GEN_5721 = opcode_2 == 4'hf ? _GEN_3671 : _GEN_5207; // @[executor.scala 466:52]
  wire [7:0] _GEN_5722 = opcode_2 == 4'hf ? _GEN_3672 : _GEN_5208; // @[executor.scala 466:52]
  wire [7:0] _GEN_5723 = opcode_2 == 4'hf ? _GEN_3673 : _GEN_5209; // @[executor.scala 466:52]
  wire [7:0] _GEN_5724 = opcode_2 == 4'hf ? _GEN_3674 : _GEN_5210; // @[executor.scala 466:52]
  wire [7:0] _GEN_5725 = opcode_2 == 4'hf ? _GEN_3675 : _GEN_5211; // @[executor.scala 466:52]
  wire [7:0] _GEN_5726 = opcode_2 == 4'hf ? _GEN_3676 : _GEN_5212; // @[executor.scala 466:52]
  wire [7:0] _GEN_5727 = opcode_2 == 4'hf ? _GEN_3677 : _GEN_5213; // @[executor.scala 466:52]
  wire [7:0] _GEN_5728 = opcode_2 == 4'hf ? _GEN_3678 : _GEN_5214; // @[executor.scala 466:52]
  wire [7:0] _GEN_5729 = opcode_2 == 4'hf ? _GEN_3679 : _GEN_5215; // @[executor.scala 466:52]
  wire [7:0] _GEN_5730 = opcode_2 == 4'hf ? _GEN_3680 : _GEN_5216; // @[executor.scala 466:52]
  wire [7:0] _GEN_5731 = opcode_2 == 4'hf ? _GEN_3681 : _GEN_5217; // @[executor.scala 466:52]
  wire [7:0] _GEN_5732 = opcode_2 == 4'hf ? _GEN_3682 : _GEN_5218; // @[executor.scala 466:52]
  wire [7:0] _GEN_5733 = opcode_2 == 4'hf ? _GEN_3683 : _GEN_5219; // @[executor.scala 466:52]
  wire [7:0] _GEN_5734 = opcode_2 == 4'hf ? _GEN_3684 : _GEN_5220; // @[executor.scala 466:52]
  wire [7:0] _GEN_5735 = opcode_2 == 4'hf ? _GEN_3685 : _GEN_5221; // @[executor.scala 466:52]
  wire [7:0] _GEN_5736 = opcode_2 == 4'hf ? _GEN_3686 : _GEN_5222; // @[executor.scala 466:52]
  wire [7:0] _GEN_5737 = opcode_2 == 4'hf ? _GEN_3687 : _GEN_5223; // @[executor.scala 466:52]
  wire [7:0] _GEN_5738 = opcode_2 == 4'hf ? _GEN_3688 : _GEN_5224; // @[executor.scala 466:52]
  wire [7:0] _GEN_5739 = opcode_2 == 4'hf ? _GEN_3689 : _GEN_5225; // @[executor.scala 466:52]
  wire [7:0] _GEN_5740 = opcode_2 == 4'hf ? _GEN_3690 : _GEN_5226; // @[executor.scala 466:52]
  wire [7:0] _GEN_5741 = opcode_2 == 4'hf ? _GEN_3691 : _GEN_5227; // @[executor.scala 466:52]
  wire [7:0] _GEN_5742 = opcode_2 == 4'hf ? _GEN_3692 : _GEN_5228; // @[executor.scala 466:52]
  wire [7:0] _GEN_5743 = opcode_2 == 4'hf ? _GEN_3693 : _GEN_5229; // @[executor.scala 466:52]
  wire [7:0] _GEN_5744 = opcode_2 == 4'hf ? _GEN_3694 : _GEN_5230; // @[executor.scala 466:52]
  wire [7:0] _GEN_5745 = opcode_2 == 4'hf ? _GEN_3695 : _GEN_5231; // @[executor.scala 466:52]
  wire [7:0] _GEN_5746 = opcode_2 == 4'hf ? _GEN_3696 : _GEN_5232; // @[executor.scala 466:52]
  wire [7:0] _GEN_5747 = opcode_2 == 4'hf ? _GEN_3697 : _GEN_5233; // @[executor.scala 466:52]
  wire [7:0] _GEN_5748 = opcode_2 == 4'hf ? _GEN_3698 : _GEN_5234; // @[executor.scala 466:52]
  wire [7:0] _GEN_5749 = opcode_2 == 4'hf ? _GEN_3699 : _GEN_5235; // @[executor.scala 466:52]
  wire [7:0] _GEN_5750 = opcode_2 == 4'hf ? _GEN_3700 : _GEN_5236; // @[executor.scala 466:52]
  wire [7:0] _GEN_5751 = opcode_2 == 4'hf ? _GEN_3701 : _GEN_5237; // @[executor.scala 466:52]
  wire [7:0] _GEN_5752 = opcode_2 == 4'hf ? _GEN_3702 : _GEN_5238; // @[executor.scala 466:52]
  wire [7:0] _GEN_5753 = opcode_2 == 4'hf ? _GEN_3703 : _GEN_5239; // @[executor.scala 466:52]
  wire [7:0] _GEN_5754 = opcode_2 == 4'hf ? _GEN_3704 : _GEN_5240; // @[executor.scala 466:52]
  wire [7:0] _GEN_5755 = opcode_2 == 4'hf ? _GEN_3705 : _GEN_5241; // @[executor.scala 466:52]
  wire [7:0] _GEN_5756 = opcode_2 == 4'hf ? _GEN_3706 : _GEN_5242; // @[executor.scala 466:52]
  wire [7:0] _GEN_5757 = opcode_2 == 4'hf ? _GEN_3707 : _GEN_5243; // @[executor.scala 466:52]
  wire [7:0] _GEN_5758 = opcode_2 == 4'hf ? _GEN_3708 : _GEN_5244; // @[executor.scala 466:52]
  wire [7:0] _GEN_5759 = opcode_2 == 4'hf ? _GEN_3709 : _GEN_5245; // @[executor.scala 466:52]
  wire [7:0] _GEN_5760 = opcode_2 == 4'hf ? _GEN_3710 : _GEN_5246; // @[executor.scala 466:52]
  wire [7:0] _GEN_5761 = opcode_2 == 4'hf ? _GEN_3711 : _GEN_5247; // @[executor.scala 466:52]
  wire [7:0] _GEN_5762 = opcode_2 == 4'hf ? _GEN_3712 : _GEN_5248; // @[executor.scala 466:52]
  wire [7:0] _GEN_5763 = opcode_2 == 4'hf ? _GEN_3713 : _GEN_5249; // @[executor.scala 466:52]
  wire [7:0] _GEN_5764 = opcode_2 == 4'hf ? _GEN_3714 : _GEN_5250; // @[executor.scala 466:52]
  wire [7:0] _GEN_5765 = opcode_2 == 4'hf ? _GEN_3715 : _GEN_5251; // @[executor.scala 466:52]
  wire [7:0] _GEN_5766 = opcode_2 == 4'hf ? _GEN_3716 : _GEN_5252; // @[executor.scala 466:52]
  wire [7:0] _GEN_5767 = opcode_2 == 4'hf ? _GEN_3717 : _GEN_5253; // @[executor.scala 466:52]
  wire [7:0] _GEN_5768 = opcode_2 == 4'hf ? _GEN_3718 : _GEN_5254; // @[executor.scala 466:52]
  wire [7:0] _GEN_5769 = opcode_2 == 4'hf ? _GEN_3719 : _GEN_5255; // @[executor.scala 466:52]
  wire [7:0] _GEN_5770 = opcode_2 == 4'hf ? _GEN_3720 : _GEN_5256; // @[executor.scala 466:52]
  wire [7:0] _GEN_5771 = opcode_2 == 4'hf ? _GEN_3721 : _GEN_5257; // @[executor.scala 466:52]
  wire [7:0] _GEN_5772 = opcode_2 == 4'hf ? _GEN_3722 : _GEN_5258; // @[executor.scala 466:52]
  wire [7:0] _GEN_5773 = opcode_2 == 4'hf ? _GEN_3723 : _GEN_5259; // @[executor.scala 466:52]
  wire [7:0] _GEN_5774 = opcode_2 == 4'hf ? _GEN_3724 : _GEN_5260; // @[executor.scala 466:52]
  wire [7:0] _GEN_5775 = opcode_2 == 4'hf ? _GEN_3725 : _GEN_5261; // @[executor.scala 466:52]
  wire [7:0] _GEN_5776 = opcode_2 == 4'hf ? _GEN_3726 : _GEN_5262; // @[executor.scala 466:52]
  wire [7:0] _GEN_5777 = opcode_2 == 4'hf ? _GEN_3727 : _GEN_5263; // @[executor.scala 466:52]
  wire [7:0] _GEN_5778 = opcode_2 == 4'hf ? _GEN_3728 : _GEN_5264; // @[executor.scala 466:52]
  wire [7:0] _GEN_5779 = opcode_2 == 4'hf ? _GEN_3729 : _GEN_5265; // @[executor.scala 466:52]
  wire [7:0] _GEN_5780 = opcode_2 == 4'hf ? _GEN_3730 : _GEN_5266; // @[executor.scala 466:52]
  wire [7:0] _GEN_5781 = opcode_2 == 4'hf ? _GEN_3731 : _GEN_5267; // @[executor.scala 466:52]
  wire [7:0] _GEN_5782 = opcode_2 == 4'hf ? _GEN_3732 : _GEN_5268; // @[executor.scala 466:52]
  wire [7:0] _GEN_5783 = opcode_2 == 4'hf ? _GEN_3733 : _GEN_5269; // @[executor.scala 466:52]
  wire [7:0] _GEN_5784 = opcode_2 == 4'hf ? _GEN_3734 : _GEN_5270; // @[executor.scala 466:52]
  wire [7:0] _GEN_5785 = opcode_2 == 4'hf ? _GEN_3735 : _GEN_5271; // @[executor.scala 466:52]
  wire [7:0] _GEN_5786 = opcode_2 == 4'hf ? _GEN_3736 : _GEN_5272; // @[executor.scala 466:52]
  wire [7:0] _GEN_5787 = opcode_2 == 4'hf ? _GEN_3737 : _GEN_5273; // @[executor.scala 466:52]
  wire [7:0] _GEN_5788 = opcode_2 == 4'hf ? _GEN_3738 : _GEN_5274; // @[executor.scala 466:52]
  wire [7:0] _GEN_5789 = opcode_2 == 4'hf ? _GEN_3739 : _GEN_5275; // @[executor.scala 466:52]
  wire [7:0] _GEN_5790 = opcode_2 == 4'hf ? _GEN_3740 : _GEN_5276; // @[executor.scala 466:52]
  wire [7:0] _GEN_5791 = opcode_2 == 4'hf ? _GEN_3741 : _GEN_5277; // @[executor.scala 466:52]
  wire [7:0] _GEN_5792 = opcode_2 == 4'hf ? _GEN_3742 : _GEN_5278; // @[executor.scala 466:52]
  wire [7:0] _GEN_5793 = opcode_2 == 4'hf ? _GEN_3743 : _GEN_5279; // @[executor.scala 466:52]
  wire [7:0] _GEN_5794 = opcode_2 == 4'hf ? _GEN_3744 : _GEN_5280; // @[executor.scala 466:52]
  wire [7:0] _GEN_5795 = opcode_2 == 4'hf ? _GEN_3745 : _GEN_5281; // @[executor.scala 466:52]
  wire [7:0] _GEN_5796 = opcode_2 == 4'hf ? _GEN_3746 : _GEN_5282; // @[executor.scala 466:52]
  wire [7:0] _GEN_5797 = opcode_2 == 4'hf ? _GEN_3747 : _GEN_5283; // @[executor.scala 466:52]
  wire [7:0] _GEN_5798 = opcode_2 == 4'hf ? _GEN_3748 : _GEN_5284; // @[executor.scala 466:52]
  wire [7:0] _GEN_5799 = opcode_2 == 4'hf ? _GEN_3749 : _GEN_5285; // @[executor.scala 466:52]
  wire [7:0] _GEN_5800 = opcode_2 == 4'hf ? _GEN_3750 : _GEN_5286; // @[executor.scala 466:52]
  wire [7:0] _GEN_5801 = opcode_2 == 4'hf ? _GEN_3751 : _GEN_5287; // @[executor.scala 466:52]
  wire [7:0] _GEN_5802 = opcode_2 == 4'hf ? _GEN_3752 : _GEN_5288; // @[executor.scala 466:52]
  wire [7:0] _GEN_5803 = opcode_2 == 4'hf ? _GEN_3753 : _GEN_5289; // @[executor.scala 466:52]
  wire [7:0] _GEN_5804 = opcode_2 == 4'hf ? _GEN_3754 : _GEN_5290; // @[executor.scala 466:52]
  wire [7:0] _GEN_5805 = opcode_2 == 4'hf ? _GEN_3755 : _GEN_5291; // @[executor.scala 466:52]
  wire [7:0] _GEN_5806 = opcode_2 == 4'hf ? _GEN_3756 : _GEN_5292; // @[executor.scala 466:52]
  wire [7:0] _GEN_5807 = opcode_2 == 4'hf ? _GEN_3757 : _GEN_5293; // @[executor.scala 466:52]
  wire [7:0] _GEN_5808 = opcode_2 == 4'hf ? _GEN_3758 : _GEN_5294; // @[executor.scala 466:52]
  wire [7:0] _GEN_5809 = opcode_2 == 4'hf ? _GEN_3759 : _GEN_5295; // @[executor.scala 466:52]
  wire [7:0] _GEN_5810 = opcode_2 == 4'hf ? _GEN_3760 : _GEN_5296; // @[executor.scala 466:52]
  wire [7:0] _GEN_5811 = opcode_2 == 4'hf ? _GEN_3761 : _GEN_5297; // @[executor.scala 466:52]
  wire [7:0] _GEN_5812 = opcode_2 == 4'hf ? _GEN_3762 : _GEN_5298; // @[executor.scala 466:52]
  wire [7:0] _GEN_5813 = opcode_2 == 4'hf ? _GEN_3763 : _GEN_5299; // @[executor.scala 466:52]
  wire [7:0] _GEN_5814 = opcode_2 == 4'hf ? _GEN_3764 : _GEN_5300; // @[executor.scala 466:52]
  wire [7:0] _GEN_5815 = opcode_2 == 4'hf ? _GEN_3765 : _GEN_5301; // @[executor.scala 466:52]
  wire [7:0] _GEN_5816 = opcode_2 == 4'hf ? _GEN_3766 : _GEN_5302; // @[executor.scala 466:52]
  wire [7:0] _GEN_5817 = opcode_2 == 4'hf ? _GEN_3767 : _GEN_5303; // @[executor.scala 466:52]
  wire [7:0] _GEN_5818 = opcode_2 == 4'hf ? _GEN_3768 : _GEN_5304; // @[executor.scala 466:52]
  wire [7:0] _GEN_5819 = opcode_2 == 4'hf ? _GEN_3769 : _GEN_5305; // @[executor.scala 466:52]
  wire [7:0] _GEN_5820 = opcode_2 == 4'hf ? _GEN_3770 : _GEN_5306; // @[executor.scala 466:52]
  wire [7:0] _GEN_5821 = opcode_2 == 4'hf ? _GEN_3771 : _GEN_5307; // @[executor.scala 466:52]
  wire [7:0] _GEN_5822 = opcode_2 == 4'hf ? _GEN_3772 : _GEN_5308; // @[executor.scala 466:52]
  wire [7:0] _GEN_5823 = opcode_2 == 4'hf ? _GEN_3773 : _GEN_5309; // @[executor.scala 466:52]
  wire [7:0] _GEN_5824 = opcode_2 == 4'hf ? _GEN_3774 : _GEN_5310; // @[executor.scala 466:52]
  wire [7:0] _GEN_5825 = opcode_2 == 4'hf ? _GEN_3775 : _GEN_5311; // @[executor.scala 466:52]
  wire [7:0] _GEN_5826 = opcode_2 == 4'hf ? _GEN_3776 : _GEN_5312; // @[executor.scala 466:52]
  wire [7:0] _GEN_5827 = opcode_2 == 4'hf ? _GEN_3777 : _GEN_5313; // @[executor.scala 466:52]
  wire [7:0] _GEN_5828 = opcode_2 == 4'hf ? _GEN_3778 : _GEN_5314; // @[executor.scala 466:52]
  wire [7:0] _GEN_5829 = opcode_2 == 4'hf ? _GEN_3779 : _GEN_5315; // @[executor.scala 466:52]
  wire [7:0] _GEN_5830 = opcode_2 == 4'hf ? _GEN_3780 : _GEN_5316; // @[executor.scala 466:52]
  wire [7:0] _GEN_5831 = opcode_2 == 4'hf ? _GEN_3781 : _GEN_5317; // @[executor.scala 466:52]
  wire [7:0] _GEN_5832 = opcode_2 == 4'hf ? _GEN_3782 : _GEN_5318; // @[executor.scala 466:52]
  wire [7:0] _GEN_5833 = opcode_2 == 4'hf ? _GEN_3783 : _GEN_5319; // @[executor.scala 466:52]
  wire [7:0] _GEN_5834 = opcode_2 == 4'hf ? _GEN_3784 : _GEN_5320; // @[executor.scala 466:52]
  wire [7:0] _GEN_5835 = opcode_2 == 4'hf ? _GEN_3785 : _GEN_5321; // @[executor.scala 466:52]
  wire [7:0] _GEN_5836 = opcode_2 == 4'hf ? _GEN_3786 : _GEN_5322; // @[executor.scala 466:52]
  wire [7:0] _GEN_5837 = opcode_2 == 4'hf ? _GEN_3787 : _GEN_5323; // @[executor.scala 466:52]
  wire [7:0] _GEN_5838 = opcode_2 == 4'hf ? _GEN_3788 : _GEN_5324; // @[executor.scala 466:52]
  wire [7:0] _GEN_5839 = opcode_2 == 4'hf ? _GEN_3789 : _GEN_5325; // @[executor.scala 466:52]
  wire [7:0] _GEN_5840 = opcode_2 == 4'hf ? _GEN_3790 : _GEN_5326; // @[executor.scala 466:52]
  wire [7:0] _GEN_5841 = opcode_2 == 4'hf ? _GEN_3791 : _GEN_5327; // @[executor.scala 466:52]
  wire [7:0] _GEN_5842 = opcode_2 == 4'hf ? _GEN_3792 : _GEN_5328; // @[executor.scala 466:52]
  wire [7:0] _GEN_5843 = opcode_2 == 4'hf ? _GEN_3793 : _GEN_5329; // @[executor.scala 466:52]
  wire [7:0] _GEN_5844 = opcode_2 == 4'hf ? _GEN_3794 : _GEN_5330; // @[executor.scala 466:52]
  wire [7:0] _GEN_5845 = opcode_2 == 4'hf ? _GEN_3795 : _GEN_5331; // @[executor.scala 466:52]
  wire [7:0] _GEN_5846 = opcode_2 == 4'hf ? _GEN_3796 : _GEN_5332; // @[executor.scala 466:52]
  wire [7:0] _GEN_5847 = opcode_2 == 4'hf ? _GEN_3797 : _GEN_5333; // @[executor.scala 466:52]
  wire [7:0] _GEN_5848 = opcode_2 == 4'hf ? _GEN_3798 : _GEN_5334; // @[executor.scala 466:52]
  wire [7:0] _GEN_5849 = opcode_2 == 4'hf ? _GEN_3799 : _GEN_5335; // @[executor.scala 466:52]
  wire [7:0] _GEN_5850 = opcode_2 == 4'hf ? _GEN_3800 : _GEN_5336; // @[executor.scala 466:52]
  wire [7:0] _GEN_5851 = opcode_2 == 4'hf ? _GEN_3801 : _GEN_5337; // @[executor.scala 466:52]
  wire [7:0] _GEN_5852 = opcode_2 == 4'hf ? _GEN_3802 : _GEN_5338; // @[executor.scala 466:52]
  wire [7:0] _GEN_5853 = opcode_2 == 4'hf ? _GEN_3803 : _GEN_5339; // @[executor.scala 466:52]
  wire [7:0] _GEN_5854 = opcode_2 == 4'hf ? _GEN_3804 : _GEN_5340; // @[executor.scala 466:52]
  wire [7:0] _GEN_5855 = opcode_2 == 4'hf ? _GEN_3805 : _GEN_5341; // @[executor.scala 466:52]
  wire [7:0] _GEN_5856 = opcode_2 == 4'hf ? _GEN_3806 : _GEN_5342; // @[executor.scala 466:52]
  wire [7:0] _GEN_5857 = opcode_2 == 4'hf ? _GEN_3807 : _GEN_5343; // @[executor.scala 466:52]
  wire [7:0] _GEN_5858 = opcode_2 == 4'hf ? _GEN_3808 : _GEN_5344; // @[executor.scala 466:52]
  wire [7:0] _GEN_5859 = opcode_2 == 4'hf ? _GEN_3809 : _GEN_5345; // @[executor.scala 466:52]
  wire [7:0] _GEN_5860 = opcode_2 == 4'hf ? _GEN_3810 : _GEN_5346; // @[executor.scala 466:52]
  wire [7:0] _GEN_5861 = opcode_2 == 4'hf ? _GEN_3811 : _GEN_5347; // @[executor.scala 466:52]
  wire [7:0] _GEN_5862 = opcode_2 == 4'hf ? _GEN_3812 : _GEN_5348; // @[executor.scala 466:52]
  wire [7:0] _GEN_5863 = opcode_2 == 4'hf ? _GEN_3813 : _GEN_5349; // @[executor.scala 466:52]
  wire [7:0] _GEN_5864 = opcode_2 == 4'hf ? _GEN_3814 : _GEN_5350; // @[executor.scala 466:52]
  wire [7:0] _GEN_5865 = opcode_2 == 4'hf ? _GEN_3815 : _GEN_5351; // @[executor.scala 466:52]
  wire [7:0] _GEN_5866 = opcode_2 == 4'hf ? _GEN_3816 : _GEN_5352; // @[executor.scala 466:52]
  wire [7:0] _GEN_5867 = opcode_2 == 4'hf ? _GEN_3817 : _GEN_5353; // @[executor.scala 466:52]
  wire [7:0] _GEN_5868 = opcode_2 == 4'hf ? _GEN_3818 : _GEN_5354; // @[executor.scala 466:52]
  wire [7:0] _GEN_5869 = opcode_2 == 4'hf ? _GEN_3819 : _GEN_5355; // @[executor.scala 466:52]
  wire [7:0] _GEN_5870 = opcode_2 == 4'hf ? _GEN_3820 : _GEN_5356; // @[executor.scala 466:52]
  wire [7:0] _GEN_5871 = opcode_2 == 4'hf ? _GEN_3821 : _GEN_5357; // @[executor.scala 466:52]
  wire [7:0] _GEN_5872 = opcode_2 == 4'hf ? _GEN_3822 : _GEN_5358; // @[executor.scala 466:52]
  wire [7:0] _GEN_5873 = opcode_2 == 4'hf ? _GEN_3823 : _GEN_5359; // @[executor.scala 466:52]
  wire [7:0] _GEN_5874 = opcode_2 == 4'hf ? _GEN_3824 : _GEN_5360; // @[executor.scala 466:52]
  wire [7:0] _GEN_5875 = opcode_2 == 4'hf ? _GEN_3825 : _GEN_5361; // @[executor.scala 466:52]
  wire [7:0] _GEN_5876 = opcode_2 == 4'hf ? _GEN_3826 : _GEN_5362; // @[executor.scala 466:52]
  wire [7:0] _GEN_5877 = opcode_2 == 4'hf ? _GEN_3827 : _GEN_5363; // @[executor.scala 466:52]
  wire [7:0] _GEN_5878 = opcode_2 == 4'hf ? _GEN_3828 : _GEN_5364; // @[executor.scala 466:52]
  wire [7:0] _GEN_5879 = opcode_2 == 4'hf ? _GEN_3829 : _GEN_5365; // @[executor.scala 466:52]
  wire [7:0] _GEN_5880 = opcode_2 == 4'hf ? _GEN_3830 : _GEN_5366; // @[executor.scala 466:52]
  wire [7:0] _GEN_5881 = opcode_2 == 4'hf ? _GEN_3831 : _GEN_5367; // @[executor.scala 466:52]
  wire [7:0] _GEN_5882 = opcode_2 == 4'hf ? _GEN_3832 : _GEN_5368; // @[executor.scala 466:52]
  wire [7:0] _GEN_5883 = opcode_2 == 4'hf ? _GEN_3833 : _GEN_5369; // @[executor.scala 466:52]
  wire [7:0] _GEN_5884 = opcode_2 == 4'hf ? _GEN_3834 : _GEN_5370; // @[executor.scala 466:52]
  wire [7:0] _GEN_5885 = opcode_2 == 4'hf ? _GEN_3835 : _GEN_5371; // @[executor.scala 466:52]
  wire [7:0] _GEN_5886 = opcode_2 == 4'hf ? _GEN_3836 : _GEN_5372; // @[executor.scala 466:52]
  wire [7:0] _GEN_5887 = opcode_2 == 4'hf ? _GEN_3837 : _GEN_5373; // @[executor.scala 466:52]
  wire [7:0] _GEN_5888 = opcode_2 == 4'hf ? _GEN_3838 : _GEN_5374; // @[executor.scala 466:52]
  wire [7:0] _GEN_5889 = opcode_2 == 4'hf ? _GEN_3839 : _GEN_5375; // @[executor.scala 466:52]
  wire [7:0] _GEN_5890 = opcode_2 == 4'hf ? _GEN_3840 : _GEN_5376; // @[executor.scala 466:52]
  wire [7:0] _GEN_5891 = opcode_2 == 4'hf ? _GEN_3841 : _GEN_5377; // @[executor.scala 466:52]
  wire [7:0] _GEN_5892 = opcode_2 == 4'hf ? _GEN_3842 : _GEN_5378; // @[executor.scala 466:52]
  wire [7:0] _GEN_5893 = opcode_2 == 4'hf ? _GEN_3843 : _GEN_5379; // @[executor.scala 466:52]
  wire [7:0] _GEN_5894 = opcode_2 == 4'hf ? _GEN_3844 : _GEN_5380; // @[executor.scala 466:52]
  wire [7:0] _GEN_5895 = opcode_2 == 4'hf ? _GEN_3845 : _GEN_5381; // @[executor.scala 466:52]
  wire [7:0] _GEN_5896 = opcode_2 == 4'hf ? _GEN_3846 : _GEN_5382; // @[executor.scala 466:52]
  wire [7:0] _GEN_5897 = opcode_2 == 4'hf ? _GEN_3847 : _GEN_5383; // @[executor.scala 466:52]
  wire [7:0] _GEN_5898 = opcode_2 == 4'hf ? _GEN_3848 : _GEN_5384; // @[executor.scala 466:52]
  wire [7:0] _GEN_5899 = opcode_2 == 4'hf ? _GEN_3849 : _GEN_5385; // @[executor.scala 466:52]
  wire [7:0] _GEN_5900 = opcode_2 == 4'hf ? _GEN_3850 : _GEN_5386; // @[executor.scala 466:52]
  wire [7:0] _GEN_5901 = opcode_2 == 4'hf ? _GEN_3851 : _GEN_5387; // @[executor.scala 466:52]
  wire [7:0] _GEN_5902 = opcode_2 == 4'hf ? _GEN_3852 : _GEN_5388; // @[executor.scala 466:52]
  wire [7:0] _GEN_5903 = opcode_2 == 4'hf ? _GEN_3853 : _GEN_5389; // @[executor.scala 466:52]
  wire [7:0] _GEN_5904 = opcode_2 == 4'hf ? _GEN_3854 : _GEN_5390; // @[executor.scala 466:52]
  wire [7:0] _GEN_5905 = opcode_2 == 4'hf ? _GEN_3855 : _GEN_5391; // @[executor.scala 466:52]
  wire [7:0] _GEN_5906 = opcode_2 == 4'hf ? _GEN_3856 : _GEN_5392; // @[executor.scala 466:52]
  wire [7:0] _GEN_5907 = opcode_2 == 4'hf ? _GEN_3857 : _GEN_5393; // @[executor.scala 466:52]
  wire [7:0] _GEN_5908 = opcode_2 == 4'hf ? _GEN_3858 : _GEN_5394; // @[executor.scala 466:52]
  wire [7:0] _GEN_5909 = opcode_2 == 4'hf ? _GEN_3859 : _GEN_5395; // @[executor.scala 466:52]
  wire [7:0] _GEN_5910 = opcode_2 == 4'hf ? _GEN_3860 : _GEN_5396; // @[executor.scala 466:52]
  wire [7:0] _GEN_5911 = opcode_2 == 4'hf ? _GEN_3861 : _GEN_5397; // @[executor.scala 466:52]
  wire [7:0] _GEN_5912 = opcode_2 == 4'hf ? _GEN_3862 : _GEN_5398; // @[executor.scala 466:52]
  wire [7:0] _GEN_5913 = opcode_2 == 4'hf ? _GEN_3863 : _GEN_5399; // @[executor.scala 466:52]
  wire [7:0] _GEN_5914 = opcode_2 == 4'hf ? _GEN_3864 : _GEN_5400; // @[executor.scala 466:52]
  wire [7:0] _GEN_5915 = opcode_2 == 4'hf ? _GEN_3865 : _GEN_5401; // @[executor.scala 466:52]
  wire [7:0] _GEN_5916 = opcode_2 == 4'hf ? _GEN_3866 : _GEN_5402; // @[executor.scala 466:52]
  wire [7:0] _GEN_5917 = opcode_2 == 4'hf ? _GEN_3867 : _GEN_5403; // @[executor.scala 466:52]
  wire [7:0] _GEN_5918 = opcode_2 == 4'hf ? _GEN_3868 : _GEN_5404; // @[executor.scala 466:52]
  wire [7:0] _GEN_5919 = opcode_2 == 4'hf ? _GEN_3869 : _GEN_5405; // @[executor.scala 466:52]
  wire [7:0] _GEN_5920 = opcode_2 == 4'hf ? _GEN_3870 : _GEN_5406; // @[executor.scala 466:52]
  wire [7:0] _GEN_5921 = opcode_2 == 4'hf ? _GEN_3871 : _GEN_5407; // @[executor.scala 466:52]
  wire [7:0] _GEN_5922 = opcode_2 == 4'hf ? _GEN_3872 : _GEN_5408; // @[executor.scala 466:52]
  wire [7:0] _GEN_5923 = opcode_2 == 4'hf ? _GEN_3873 : _GEN_5409; // @[executor.scala 466:52]
  wire [7:0] _GEN_5924 = opcode_2 == 4'hf ? _GEN_3874 : _GEN_5410; // @[executor.scala 466:52]
  wire [7:0] _GEN_5925 = opcode_2 == 4'hf ? _GEN_3875 : _GEN_5411; // @[executor.scala 466:52]
  wire [7:0] _GEN_5926 = opcode_2 == 4'hf ? _GEN_3876 : _GEN_5412; // @[executor.scala 466:52]
  wire [7:0] _GEN_5927 = opcode_2 == 4'hf ? _GEN_3877 : _GEN_5413; // @[executor.scala 466:52]
  wire [7:0] _GEN_5928 = opcode_2 == 4'hf ? _GEN_3878 : _GEN_5414; // @[executor.scala 466:52]
  wire [7:0] _GEN_5929 = opcode_2 == 4'hf ? _GEN_3879 : _GEN_5415; // @[executor.scala 466:52]
  wire [7:0] _GEN_5930 = opcode_2 == 4'hf ? _GEN_3880 : _GEN_5416; // @[executor.scala 466:52]
  wire [7:0] _GEN_5931 = opcode_2 == 4'hf ? _GEN_3881 : _GEN_5417; // @[executor.scala 466:52]
  wire [7:0] _GEN_5932 = opcode_2 == 4'hf ? _GEN_3882 : _GEN_5418; // @[executor.scala 466:52]
  wire [7:0] _GEN_5933 = opcode_2 == 4'hf ? _GEN_3883 : _GEN_5419; // @[executor.scala 466:52]
  wire [7:0] _GEN_5934 = opcode_2 == 4'hf ? _GEN_3884 : _GEN_5420; // @[executor.scala 466:52]
  wire [7:0] _GEN_5935 = opcode_2 == 4'hf ? _GEN_3885 : _GEN_5421; // @[executor.scala 466:52]
  wire [7:0] _GEN_5936 = opcode_2 == 4'hf ? _GEN_3886 : _GEN_5422; // @[executor.scala 466:52]
  wire [7:0] _GEN_5937 = opcode_2 == 4'hf ? _GEN_3887 : _GEN_5423; // @[executor.scala 466:52]
  wire [7:0] _GEN_5938 = opcode_2 == 4'hf ? _GEN_3888 : _GEN_5424; // @[executor.scala 466:52]
  wire [7:0] _GEN_5939 = opcode_2 == 4'hf ? _GEN_3889 : _GEN_5425; // @[executor.scala 466:52]
  wire [7:0] _GEN_5940 = opcode_2 == 4'hf ? _GEN_3890 : _GEN_5426; // @[executor.scala 466:52]
  wire [7:0] _GEN_5941 = opcode_2 == 4'hf ? _GEN_3891 : _GEN_5427; // @[executor.scala 466:52]
  wire [7:0] _GEN_5942 = opcode_2 == 4'hf ? _GEN_3892 : _GEN_5428; // @[executor.scala 466:52]
  wire [7:0] _GEN_5943 = opcode_2 == 4'hf ? _GEN_3893 : _GEN_5429; // @[executor.scala 466:52]
  wire [7:0] _GEN_5944 = opcode_2 == 4'hf ? _GEN_3894 : _GEN_5430; // @[executor.scala 466:52]
  wire [7:0] _GEN_5945 = opcode_2 == 4'hf ? _GEN_3895 : _GEN_5431; // @[executor.scala 466:52]
  wire [7:0] _GEN_5946 = opcode_2 == 4'hf ? _GEN_3896 : _GEN_5432; // @[executor.scala 466:52]
  wire [7:0] _GEN_5947 = opcode_2 == 4'hf ? _GEN_3897 : _GEN_5433; // @[executor.scala 466:52]
  wire [7:0] _GEN_5948 = opcode_2 == 4'hf ? _GEN_3898 : _GEN_5434; // @[executor.scala 466:52]
  wire [7:0] _GEN_5949 = opcode_2 == 4'hf ? _GEN_3899 : _GEN_5435; // @[executor.scala 466:52]
  wire [7:0] _GEN_5950 = opcode_2 == 4'hf ? _GEN_3900 : _GEN_5436; // @[executor.scala 466:52]
  wire [7:0] _GEN_5951 = opcode_2 == 4'hf ? _GEN_3901 : _GEN_5437; // @[executor.scala 466:52]
  wire [7:0] _GEN_5952 = opcode_2 == 4'hf ? _GEN_3902 : _GEN_5438; // @[executor.scala 466:52]
  wire [7:0] _GEN_5953 = opcode_2 == 4'hf ? _GEN_3903 : _GEN_5439; // @[executor.scala 466:52]
  wire [7:0] _GEN_5954 = opcode_2 == 4'hf ? _GEN_3904 : _GEN_5440; // @[executor.scala 466:52]
  wire [7:0] _GEN_5955 = opcode_2 == 4'hf ? _GEN_3905 : _GEN_5441; // @[executor.scala 466:52]
  wire [7:0] _GEN_5956 = opcode_2 == 4'hf ? _GEN_3906 : _GEN_5442; // @[executor.scala 466:52]
  wire [7:0] _GEN_5957 = opcode_2 == 4'hf ? _GEN_3907 : _GEN_5443; // @[executor.scala 466:52]
  wire [7:0] _GEN_5958 = opcode_2 == 4'hf ? _GEN_3908 : _GEN_5444; // @[executor.scala 466:52]
  wire [7:0] _GEN_5959 = opcode_2 == 4'hf ? _GEN_3909 : _GEN_5445; // @[executor.scala 466:52]
  wire [7:0] _GEN_5960 = opcode_2 == 4'hf ? _GEN_3910 : _GEN_5446; // @[executor.scala 466:52]
  wire [7:0] _GEN_5961 = opcode_2 == 4'hf ? _GEN_3911 : _GEN_5447; // @[executor.scala 466:52]
  wire [7:0] _GEN_5962 = opcode_2 == 4'hf ? _GEN_3912 : _GEN_5448; // @[executor.scala 466:52]
  wire [7:0] _GEN_5963 = opcode_2 == 4'hf ? _GEN_3913 : _GEN_5449; // @[executor.scala 466:52]
  wire [7:0] _GEN_5964 = opcode_2 == 4'hf ? _GEN_3914 : _GEN_5450; // @[executor.scala 466:52]
  wire [7:0] _GEN_5965 = opcode_2 == 4'hf ? _GEN_3915 : _GEN_5451; // @[executor.scala 466:52]
  wire [7:0] _GEN_5966 = opcode_2 == 4'hf ? _GEN_3916 : _GEN_5452; // @[executor.scala 466:52]
  wire [7:0] _GEN_5967 = opcode_2 == 4'hf ? _GEN_3917 : _GEN_5453; // @[executor.scala 466:52]
  wire [7:0] _GEN_5968 = opcode_2 == 4'hf ? _GEN_3918 : _GEN_5454; // @[executor.scala 466:52]
  wire [7:0] _GEN_5969 = opcode_2 == 4'hf ? _GEN_3919 : _GEN_5455; // @[executor.scala 466:52]
  wire [7:0] _GEN_5970 = opcode_2 == 4'hf ? _GEN_3920 : _GEN_5456; // @[executor.scala 466:52]
  wire [7:0] _GEN_5971 = opcode_2 == 4'hf ? _GEN_3921 : _GEN_5457; // @[executor.scala 466:52]
  wire [7:0] _GEN_5972 = opcode_2 == 4'hf ? _GEN_3922 : _GEN_5458; // @[executor.scala 466:52]
  wire [7:0] _GEN_5973 = opcode_2 == 4'hf ? _GEN_3923 : _GEN_5459; // @[executor.scala 466:52]
  wire [7:0] _GEN_5974 = opcode_2 == 4'hf ? _GEN_3924 : _GEN_5460; // @[executor.scala 466:52]
  wire [7:0] _GEN_5975 = opcode_2 == 4'hf ? _GEN_3925 : _GEN_5461; // @[executor.scala 466:52]
  wire [7:0] _GEN_5976 = opcode_2 == 4'hf ? _GEN_3926 : _GEN_5462; // @[executor.scala 466:52]
  wire [7:0] _GEN_5977 = opcode_2 == 4'hf ? _GEN_3927 : _GEN_5463; // @[executor.scala 466:52]
  wire [7:0] _GEN_5978 = opcode_2 == 4'hf ? _GEN_3928 : _GEN_5464; // @[executor.scala 466:52]
  wire [7:0] _GEN_5979 = opcode_2 == 4'hf ? _GEN_3929 : _GEN_5465; // @[executor.scala 466:52]
  wire [7:0] _GEN_5980 = opcode_2 == 4'hf ? _GEN_3930 : _GEN_5466; // @[executor.scala 466:52]
  wire [7:0] _GEN_5981 = opcode_2 == 4'hf ? _GEN_3931 : _GEN_5467; // @[executor.scala 466:52]
  wire [7:0] _GEN_5982 = opcode_2 == 4'hf ? _GEN_3932 : _GEN_5468; // @[executor.scala 466:52]
  wire [7:0] _GEN_5983 = opcode_2 == 4'hf ? _GEN_3933 : _GEN_5469; // @[executor.scala 466:52]
  wire [7:0] _GEN_5984 = opcode_2 == 4'hf ? _GEN_3934 : _GEN_5470; // @[executor.scala 466:52]
  wire [7:0] _GEN_5985 = opcode_2 == 4'hf ? _GEN_3935 : _GEN_5471; // @[executor.scala 466:52]
  wire [7:0] _GEN_5986 = opcode_2 == 4'hf ? _GEN_3936 : _GEN_5472; // @[executor.scala 466:52]
  wire [7:0] _GEN_5987 = opcode_2 == 4'hf ? _GEN_3937 : _GEN_5473; // @[executor.scala 466:52]
  wire [7:0] _GEN_5988 = opcode_2 == 4'hf ? _GEN_3938 : _GEN_5474; // @[executor.scala 466:52]
  wire [7:0] _GEN_5989 = opcode_2 == 4'hf ? _GEN_3939 : _GEN_5475; // @[executor.scala 466:52]
  wire [7:0] _GEN_5990 = opcode_2 == 4'hf ? _GEN_3940 : _GEN_5476; // @[executor.scala 466:52]
  wire [7:0] _GEN_5991 = opcode_2 == 4'hf ? _GEN_3941 : _GEN_5477; // @[executor.scala 466:52]
  wire [7:0] _GEN_5992 = opcode_2 == 4'hf ? _GEN_3942 : _GEN_5478; // @[executor.scala 466:52]
  wire [7:0] _GEN_5993 = opcode_2 == 4'hf ? _GEN_3943 : _GEN_5479; // @[executor.scala 466:52]
  wire [7:0] _GEN_5994 = opcode_2 == 4'hf ? _GEN_3944 : _GEN_5480; // @[executor.scala 466:52]
  wire [7:0] _GEN_5995 = opcode_2 == 4'hf ? _GEN_3945 : _GEN_5481; // @[executor.scala 466:52]
  wire [7:0] _GEN_5996 = opcode_2 == 4'hf ? _GEN_3946 : _GEN_5482; // @[executor.scala 466:52]
  wire [7:0] _GEN_5997 = opcode_2 == 4'hf ? _GEN_3947 : _GEN_5483; // @[executor.scala 466:52]
  wire [7:0] _GEN_5998 = opcode_2 == 4'hf ? _GEN_3948 : _GEN_5484; // @[executor.scala 466:52]
  wire [7:0] _GEN_5999 = opcode_2 == 4'hf ? _GEN_3949 : _GEN_5485; // @[executor.scala 466:52]
  wire [7:0] _GEN_6000 = opcode_2 == 4'hf ? _GEN_3950 : _GEN_5486; // @[executor.scala 466:52]
  wire [7:0] _GEN_6001 = opcode_2 == 4'hf ? _GEN_3951 : _GEN_5487; // @[executor.scala 466:52]
  wire [7:0] _GEN_6002 = opcode_2 == 4'hf ? _GEN_3952 : _GEN_5488; // @[executor.scala 466:52]
  wire [7:0] _GEN_6003 = opcode_2 == 4'hf ? _GEN_3953 : _GEN_5489; // @[executor.scala 466:52]
  wire [7:0] _GEN_6004 = opcode_2 == 4'hf ? _GEN_3954 : _GEN_5490; // @[executor.scala 466:52]
  wire [7:0] _GEN_6005 = opcode_2 == 4'hf ? _GEN_3955 : _GEN_5491; // @[executor.scala 466:52]
  wire [7:0] _GEN_6006 = opcode_2 == 4'hf ? _GEN_3956 : _GEN_5492; // @[executor.scala 466:52]
  wire [7:0] _GEN_6007 = opcode_2 == 4'hf ? _GEN_3957 : _GEN_5493; // @[executor.scala 466:52]
  wire [7:0] _GEN_6008 = opcode_2 == 4'hf ? _GEN_3958 : _GEN_5494; // @[executor.scala 466:52]
  wire [7:0] _GEN_6009 = opcode_2 == 4'hf ? _GEN_3959 : _GEN_5495; // @[executor.scala 466:52]
  wire [7:0] _GEN_6010 = opcode_2 == 4'hf ? _GEN_3960 : _GEN_5496; // @[executor.scala 466:52]
  wire [7:0] _GEN_6011 = opcode_2 == 4'hf ? _GEN_3961 : _GEN_5497; // @[executor.scala 466:52]
  wire [7:0] _GEN_6012 = opcode_2 == 4'hf ? _GEN_3962 : _GEN_5498; // @[executor.scala 466:52]
  wire [7:0] _GEN_6013 = opcode_2 == 4'hf ? _GEN_3963 : _GEN_5499; // @[executor.scala 466:52]
  wire [7:0] _GEN_6014 = opcode_2 == 4'hf ? _GEN_3964 : _GEN_5500; // @[executor.scala 466:52]
  wire [7:0] _GEN_6015 = opcode_2 == 4'hf ? _GEN_3965 : _GEN_5501; // @[executor.scala 466:52]
  wire [7:0] _GEN_6016 = opcode_2 == 4'hf ? _GEN_3966 : _GEN_5502; // @[executor.scala 466:52]
  wire [7:0] _GEN_6017 = opcode_2 == 4'hf ? _GEN_3967 : _GEN_5503; // @[executor.scala 466:52]
  wire [7:0] _GEN_6018 = opcode_2 == 4'hf ? _GEN_3968 : _GEN_5504; // @[executor.scala 466:52]
  wire [7:0] _GEN_6019 = opcode_2 == 4'hf ? _GEN_3969 : _GEN_5505; // @[executor.scala 466:52]
  wire [7:0] _GEN_6020 = opcode_2 == 4'hf ? _GEN_3970 : _GEN_5506; // @[executor.scala 466:52]
  wire [7:0] _GEN_6021 = opcode_2 == 4'hf ? _GEN_3971 : _GEN_5507; // @[executor.scala 466:52]
  wire [7:0] _GEN_6022 = opcode_2 == 4'hf ? _GEN_3972 : _GEN_5508; // @[executor.scala 466:52]
  wire [7:0] _GEN_6023 = opcode_2 == 4'hf ? _GEN_3973 : _GEN_5509; // @[executor.scala 466:52]
  wire [7:0] _GEN_6024 = opcode_2 == 4'hf ? _GEN_3974 : _GEN_5510; // @[executor.scala 466:52]
  wire [7:0] _GEN_6025 = opcode_2 == 4'hf ? _GEN_3975 : _GEN_5511; // @[executor.scala 466:52]
  wire [7:0] _GEN_6026 = opcode_2 == 4'hf ? _GEN_3976 : _GEN_5512; // @[executor.scala 466:52]
  wire [7:0] _GEN_6027 = opcode_2 == 4'hf ? _GEN_3977 : _GEN_5513; // @[executor.scala 466:52]
  wire [7:0] _GEN_6028 = opcode_2 == 4'hf ? _GEN_3978 : _GEN_5514; // @[executor.scala 466:52]
  wire [7:0] _GEN_6029 = opcode_2 == 4'hf ? _GEN_3979 : _GEN_5515; // @[executor.scala 466:52]
  wire [7:0] _GEN_6030 = opcode_2 == 4'hf ? _GEN_3980 : _GEN_5516; // @[executor.scala 466:52]
  wire [7:0] _GEN_6031 = opcode_2 == 4'hf ? _GEN_3981 : _GEN_5517; // @[executor.scala 466:52]
  wire [7:0] _GEN_6032 = opcode_2 == 4'hf ? _GEN_3982 : _GEN_5518; // @[executor.scala 466:52]
  wire [7:0] _GEN_6033 = opcode_2 == 4'hf ? _GEN_3983 : _GEN_5519; // @[executor.scala 466:52]
  wire [7:0] _GEN_6034 = opcode_2 == 4'hf ? _GEN_3984 : _GEN_5520; // @[executor.scala 466:52]
  wire [7:0] _GEN_6035 = opcode_2 == 4'hf ? _GEN_3985 : _GEN_5521; // @[executor.scala 466:52]
  wire [7:0] _GEN_6036 = opcode_2 == 4'hf ? _GEN_3986 : _GEN_5522; // @[executor.scala 466:52]
  wire [7:0] _GEN_6037 = opcode_2 == 4'hf ? _GEN_3987 : _GEN_5523; // @[executor.scala 466:52]
  wire [7:0] _GEN_6038 = opcode_2 == 4'hf ? _GEN_3988 : _GEN_5524; // @[executor.scala 466:52]
  wire [7:0] _GEN_6039 = opcode_2 == 4'hf ? _GEN_3989 : _GEN_5525; // @[executor.scala 466:52]
  wire [7:0] _GEN_6040 = opcode_2 == 4'hf ? _GEN_3990 : _GEN_5526; // @[executor.scala 466:52]
  wire [7:0] _GEN_6041 = opcode_2 == 4'hf ? _GEN_3991 : _GEN_5527; // @[executor.scala 466:52]
  wire [7:0] _GEN_6042 = opcode_2 == 4'hf ? _GEN_3992 : _GEN_5528; // @[executor.scala 466:52]
  wire [7:0] _GEN_6043 = opcode_2 == 4'hf ? _GEN_3993 : _GEN_5529; // @[executor.scala 466:52]
  wire [7:0] _GEN_6044 = opcode_2 == 4'hf ? _GEN_3994 : _GEN_5530; // @[executor.scala 466:52]
  wire [7:0] _GEN_6045 = opcode_2 == 4'hf ? _GEN_3995 : _GEN_5531; // @[executor.scala 466:52]
  wire [7:0] _GEN_6046 = opcode_2 == 4'hf ? _GEN_3996 : _GEN_5532; // @[executor.scala 466:52]
  wire [7:0] _GEN_6047 = opcode_2 == 4'hf ? _GEN_3997 : _GEN_5533; // @[executor.scala 466:52]
  wire [7:0] _GEN_6048 = opcode_2 == 4'hf ? _GEN_3998 : _GEN_5534; // @[executor.scala 466:52]
  wire [7:0] _GEN_6049 = opcode_2 == 4'hf ? _GEN_3999 : _GEN_5535; // @[executor.scala 466:52]
  wire [7:0] _GEN_6050 = opcode_2 == 4'hf ? _GEN_4000 : _GEN_5536; // @[executor.scala 466:52]
  wire [7:0] _GEN_6051 = opcode_2 == 4'hf ? _GEN_4001 : _GEN_5537; // @[executor.scala 466:52]
  wire [7:0] _GEN_6052 = opcode_2 == 4'hf ? _GEN_4002 : _GEN_5538; // @[executor.scala 466:52]
  wire [7:0] _GEN_6053 = opcode_2 == 4'hf ? _GEN_4003 : _GEN_5539; // @[executor.scala 466:52]
  wire [7:0] _GEN_6054 = opcode_2 == 4'hf ? _GEN_4004 : _GEN_5540; // @[executor.scala 466:52]
  wire [7:0] _GEN_6055 = opcode_2 == 4'hf ? _GEN_4005 : _GEN_5541; // @[executor.scala 466:52]
  wire [7:0] _GEN_6056 = opcode_2 == 4'hf ? _GEN_4006 : _GEN_5542; // @[executor.scala 466:52]
  wire [7:0] _GEN_6057 = opcode_2 == 4'hf ? _GEN_4007 : _GEN_5543; // @[executor.scala 466:52]
  wire [7:0] _GEN_6058 = opcode_2 == 4'hf ? _GEN_4008 : _GEN_5544; // @[executor.scala 466:52]
  wire [7:0] _GEN_6059 = opcode_2 == 4'hf ? _GEN_4009 : _GEN_5545; // @[executor.scala 466:52]
  wire [7:0] _GEN_6060 = opcode_2 == 4'hf ? _GEN_4010 : _GEN_5546; // @[executor.scala 466:52]
  wire [7:0] _GEN_6061 = opcode_2 == 4'hf ? _GEN_4011 : _GEN_5547; // @[executor.scala 466:52]
  wire [7:0] _GEN_6062 = opcode_2 == 4'hf ? _GEN_4012 : _GEN_5548; // @[executor.scala 466:52]
  wire [7:0] _GEN_6063 = opcode_2 == 4'hf ? _GEN_4013 : _GEN_5549; // @[executor.scala 466:52]
  wire [7:0] _GEN_6064 = opcode_2 == 4'hf ? _GEN_4014 : _GEN_5550; // @[executor.scala 466:52]
  wire [7:0] _GEN_6065 = opcode_2 == 4'hf ? _GEN_4015 : _GEN_5551; // @[executor.scala 466:52]
  wire [7:0] _GEN_6066 = opcode_2 == 4'hf ? _GEN_4016 : _GEN_5552; // @[executor.scala 466:52]
  wire [7:0] _GEN_6067 = opcode_2 == 4'hf ? _GEN_4017 : _GEN_5553; // @[executor.scala 466:52]
  wire [7:0] _GEN_6068 = opcode_2 == 4'hf ? _GEN_4018 : _GEN_5554; // @[executor.scala 466:52]
  wire [7:0] _GEN_6069 = opcode_2 == 4'hf ? _GEN_4019 : _GEN_5555; // @[executor.scala 466:52]
  wire [7:0] _GEN_6070 = opcode_2 == 4'hf ? _GEN_4020 : _GEN_5556; // @[executor.scala 466:52]
  wire [7:0] _GEN_6071 = opcode_2 == 4'hf ? _GEN_4021 : _GEN_5557; // @[executor.scala 466:52]
  wire [7:0] _GEN_6072 = opcode_2 == 4'hf ? _GEN_4022 : _GEN_5558; // @[executor.scala 466:52]
  wire [7:0] _GEN_6073 = opcode_2 == 4'hf ? _GEN_4023 : _GEN_5559; // @[executor.scala 466:52]
  wire [7:0] _GEN_6074 = opcode_2 == 4'hf ? _GEN_4024 : _GEN_5560; // @[executor.scala 466:52]
  wire [7:0] _GEN_6075 = opcode_2 == 4'hf ? _GEN_4025 : _GEN_5561; // @[executor.scala 466:52]
  wire [7:0] _GEN_6076 = opcode_2 == 4'hf ? _GEN_4026 : _GEN_5562; // @[executor.scala 466:52]
  wire [7:0] _GEN_6077 = opcode_2 == 4'hf ? _GEN_4027 : _GEN_5563; // @[executor.scala 466:52]
  wire [7:0] _GEN_6078 = opcode_2 == 4'hf ? _GEN_4028 : _GEN_5564; // @[executor.scala 466:52]
  wire [7:0] _GEN_6079 = opcode_2 == 4'hf ? _GEN_4029 : _GEN_5565; // @[executor.scala 466:52]
  wire [7:0] _GEN_6080 = opcode_2 == 4'hf ? _GEN_4030 : _GEN_5566; // @[executor.scala 466:52]
  wire [7:0] _GEN_6081 = opcode_2 == 4'hf ? _GEN_4031 : _GEN_5567; // @[executor.scala 466:52]
  wire [7:0] _GEN_6082 = opcode_2 == 4'hf ? _GEN_4032 : _GEN_5568; // @[executor.scala 466:52]
  wire [7:0] _GEN_6083 = opcode_2 == 4'hf ? _GEN_4033 : _GEN_5569; // @[executor.scala 466:52]
  wire [7:0] _GEN_6084 = opcode_2 == 4'hf ? _GEN_4034 : _GEN_5570; // @[executor.scala 466:52]
  wire [7:0] _GEN_6085 = opcode_2 == 4'hf ? _GEN_4035 : _GEN_5571; // @[executor.scala 466:52]
  wire [7:0] _GEN_6086 = opcode_2 == 4'hf ? _GEN_4036 : _GEN_5572; // @[executor.scala 466:52]
  wire [7:0] _GEN_6087 = opcode_2 == 4'hf ? _GEN_4037 : _GEN_5573; // @[executor.scala 466:52]
  wire [7:0] _GEN_6088 = opcode_2 == 4'hf ? _GEN_4038 : _GEN_5574; // @[executor.scala 466:52]
  wire [7:0] _GEN_6089 = opcode_2 == 4'hf ? _GEN_4039 : _GEN_5575; // @[executor.scala 466:52]
  wire [7:0] _GEN_6090 = opcode_2 == 4'hf ? _GEN_4040 : _GEN_5576; // @[executor.scala 466:52]
  wire [7:0] _GEN_6091 = opcode_2 == 4'hf ? _GEN_4041 : _GEN_5577; // @[executor.scala 466:52]
  wire [7:0] _GEN_6092 = opcode_2 == 4'hf ? _GEN_4042 : _GEN_5578; // @[executor.scala 466:52]
  wire [7:0] _GEN_6093 = opcode_2 == 4'hf ? _GEN_4043 : _GEN_5579; // @[executor.scala 466:52]
  wire [7:0] _GEN_6094 = opcode_2 == 4'hf ? _GEN_4044 : _GEN_5580; // @[executor.scala 466:52]
  wire [7:0] _GEN_6095 = opcode_2 == 4'hf ? _GEN_4045 : _GEN_5581; // @[executor.scala 466:52]
  wire [7:0] _GEN_6096 = opcode_2 == 4'hf ? _GEN_4046 : _GEN_5582; // @[executor.scala 466:52]
  wire [7:0] _GEN_6097 = opcode_2 == 4'hf ? _GEN_4047 : _GEN_5583; // @[executor.scala 466:52]
  wire [7:0] _GEN_6098 = opcode_2 == 4'hf ? _GEN_4048 : _GEN_5584; // @[executor.scala 466:52]
  wire [7:0] _GEN_6099 = opcode_2 == 4'hf ? _GEN_4049 : _GEN_5585; // @[executor.scala 466:52]
  wire [7:0] _GEN_6100 = opcode_2 == 4'hf ? _GEN_4050 : _GEN_5586; // @[executor.scala 466:52]
  wire [7:0] _GEN_6101 = opcode_2 == 4'hf ? _GEN_4051 : _GEN_5587; // @[executor.scala 466:52]
  wire [7:0] _GEN_6102 = opcode_2 == 4'hf ? _GEN_4052 : _GEN_5588; // @[executor.scala 466:52]
  wire [7:0] _GEN_6103 = opcode_2 == 4'hf ? _GEN_4053 : _GEN_5589; // @[executor.scala 466:52]
  wire [7:0] _GEN_6104 = opcode_2 == 4'hf ? _GEN_4054 : _GEN_5590; // @[executor.scala 466:52]
  wire [7:0] _GEN_6105 = opcode_2 == 4'hf ? _GEN_4055 : _GEN_5591; // @[executor.scala 466:52]
  wire [7:0] _GEN_6106 = opcode_2 == 4'hf ? _GEN_4056 : _GEN_5592; // @[executor.scala 466:52]
  wire [7:0] _GEN_6107 = opcode_2 == 4'hf ? _GEN_4057 : _GEN_5593; // @[executor.scala 466:52]
  wire [7:0] _GEN_6108 = opcode_2 == 4'hf ? _GEN_4058 : _GEN_5594; // @[executor.scala 466:52]
  wire [7:0] _GEN_6109 = opcode_2 == 4'hf ? _GEN_4059 : _GEN_5595; // @[executor.scala 466:52]
  wire [7:0] _GEN_6110 = opcode_2 == 4'hf ? _GEN_4060 : _GEN_5596; // @[executor.scala 466:52]
  wire [7:0] _GEN_6111 = opcode_2 == 4'hf ? _GEN_4061 : _GEN_5597; // @[executor.scala 466:52]
  wire [7:0] _GEN_6112 = opcode_2 == 4'hf ? _GEN_4062 : _GEN_5598; // @[executor.scala 466:52]
  wire [7:0] _GEN_6113 = opcode_2 == 4'hf ? _GEN_4063 : _GEN_5599; // @[executor.scala 466:52]
  wire [7:0] _GEN_6114 = opcode_2 == 4'hf ? _GEN_4064 : _GEN_5600; // @[executor.scala 466:52]
  wire [7:0] _GEN_6115 = opcode_2 == 4'hf ? _GEN_4065 : _GEN_5601; // @[executor.scala 466:52]
  wire [7:0] _GEN_6116 = opcode_2 == 4'hf ? _GEN_4066 : _GEN_5602; // @[executor.scala 466:52]
  wire [7:0] _GEN_6117 = opcode_2 == 4'hf ? _GEN_4067 : _GEN_5603; // @[executor.scala 466:52]
  wire [7:0] _GEN_6118 = opcode_2 == 4'hf ? _GEN_4068 : _GEN_5604; // @[executor.scala 466:52]
  wire [7:0] _GEN_6119 = opcode_2 == 4'hf ? _GEN_4069 : _GEN_5605; // @[executor.scala 466:52]
  wire [7:0] _GEN_6120 = opcode_2 == 4'hf ? _GEN_4070 : _GEN_5606; // @[executor.scala 466:52]
  wire [7:0] _GEN_6121 = opcode_2 == 4'hf ? _GEN_4071 : _GEN_5607; // @[executor.scala 466:52]
  wire [7:0] _GEN_6122 = opcode_2 == 4'hf ? _GEN_4072 : _GEN_5608; // @[executor.scala 466:52]
  wire [7:0] _GEN_6123 = opcode_2 == 4'hf ? _GEN_4073 : _GEN_5609; // @[executor.scala 466:52]
  wire [7:0] _GEN_6124 = opcode_2 == 4'hf ? _GEN_4074 : _GEN_5610; // @[executor.scala 466:52]
  wire [7:0] _GEN_6125 = opcode_2 == 4'hf ? _GEN_4075 : _GEN_5611; // @[executor.scala 466:52]
  wire [7:0] _GEN_6126 = opcode_2 == 4'hf ? _GEN_4076 : _GEN_5612; // @[executor.scala 466:52]
  wire [7:0] _GEN_6127 = opcode_2 == 4'hf ? _GEN_4077 : _GEN_5613; // @[executor.scala 466:52]
  wire [7:0] _GEN_6128 = opcode_2 == 4'hf ? _GEN_4078 : _GEN_5614; // @[executor.scala 466:52]
  wire [7:0] _GEN_6129 = opcode_2 == 4'hf ? _GEN_4079 : _GEN_5615; // @[executor.scala 466:52]
  wire [7:0] _GEN_6130 = opcode_2 == 4'hf ? _GEN_4080 : _GEN_5616; // @[executor.scala 466:52]
  wire [7:0] _GEN_6131 = opcode_2 == 4'hf ? _GEN_4081 : _GEN_5617; // @[executor.scala 466:52]
  wire [7:0] _GEN_6132 = opcode_2 == 4'hf ? _GEN_4082 : _GEN_5618; // @[executor.scala 466:52]
  wire [7:0] _GEN_6133 = opcode_2 == 4'hf ? _GEN_4083 : _GEN_5619; // @[executor.scala 466:52]
  wire [7:0] _GEN_6134 = opcode_2 == 4'hf ? _GEN_4084 : _GEN_5620; // @[executor.scala 466:52]
  wire [7:0] _GEN_6135 = opcode_2 == 4'hf ? _GEN_4085 : _GEN_5621; // @[executor.scala 466:52]
  wire [7:0] _GEN_6136 = opcode_2 == 4'hf ? _GEN_4086 : _GEN_5622; // @[executor.scala 466:52]
  wire [7:0] _GEN_6137 = opcode_2 == 4'hf ? _GEN_4087 : _GEN_5623; // @[executor.scala 466:52]
  wire [7:0] _GEN_6138 = opcode_2 == 4'hf ? _GEN_4088 : _GEN_5624; // @[executor.scala 466:52]
  wire [7:0] _GEN_6139 = opcode_2 == 4'hf ? _GEN_4089 : _GEN_5625; // @[executor.scala 466:52]
  wire [7:0] _GEN_6140 = opcode_2 == 4'hf ? _GEN_4090 : _GEN_5626; // @[executor.scala 466:52]
  wire [7:0] _GEN_6141 = opcode_2 == 4'hf ? _GEN_4091 : _GEN_5627; // @[executor.scala 466:52]
  wire [7:0] _GEN_6142 = opcode_2 == 4'hf ? _GEN_4092 : _GEN_5628; // @[executor.scala 466:52]
  wire [7:0] _GEN_6143 = opcode_2 == 4'hf ? _GEN_4093 : _GEN_5629; // @[executor.scala 466:52]
  wire [7:0] _GEN_6144 = opcode_2 == 4'hf ? _GEN_4094 : _GEN_5630; // @[executor.scala 466:52]
  wire [7:0] _GEN_6145 = opcode_2 == 4'hf ? _GEN_4095 : _GEN_5631; // @[executor.scala 466:52]
  wire [7:0] _GEN_6146 = opcode_2 == 4'hf ? _GEN_4096 : _GEN_5632; // @[executor.scala 466:52]
  wire [7:0] _GEN_6147 = opcode_2 == 4'hf ? _GEN_4097 : _GEN_5633; // @[executor.scala 466:52]
  wire [7:0] _GEN_6148 = opcode_2 == 4'hf ? _GEN_4098 : _GEN_5634; // @[executor.scala 466:52]
  wire [7:0] _GEN_6149 = opcode_2 == 4'hf ? _GEN_4099 : _GEN_5635; // @[executor.scala 466:52]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_2_3 = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire [7:0] _GEN_9098 = {{2'd0}, dst_offset_3}; // @[executor.scala 473:49]
  wire [7:0] byte_1536 = field_3[7:0]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6150 = mask_3[0] ? byte_1536 : _GEN_5638; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1537 = field_3[15:8]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6151 = mask_3[1] ? byte_1537 : _GEN_5639; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1538 = field_3[23:16]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6152 = mask_3[2] ? byte_1538 : _GEN_5640; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] byte_1539 = field_3[31:24]; // @[executor.scala 475:56]
  wire [7:0] _GEN_6153 = mask_3[3] ? byte_1539 : _GEN_5641; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6154 = _GEN_9098 == 8'h0 ? _GEN_6150 : _GEN_5638; // @[executor.scala 473:84]
  wire [7:0] _GEN_6155 = _GEN_9098 == 8'h0 ? _GEN_6151 : _GEN_5639; // @[executor.scala 473:84]
  wire [7:0] _GEN_6156 = _GEN_9098 == 8'h0 ? _GEN_6152 : _GEN_5640; // @[executor.scala 473:84]
  wire [7:0] _GEN_6157 = _GEN_9098 == 8'h0 ? _GEN_6153 : _GEN_5641; // @[executor.scala 473:84]
  wire [7:0] _GEN_6158 = mask_3[0] ? byte_1536 : _GEN_5642; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6159 = mask_3[1] ? byte_1537 : _GEN_5643; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6160 = mask_3[2] ? byte_1538 : _GEN_5644; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6161 = mask_3[3] ? byte_1539 : _GEN_5645; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6162 = _GEN_9098 == 8'h1 ? _GEN_6158 : _GEN_5642; // @[executor.scala 473:84]
  wire [7:0] _GEN_6163 = _GEN_9098 == 8'h1 ? _GEN_6159 : _GEN_5643; // @[executor.scala 473:84]
  wire [7:0] _GEN_6164 = _GEN_9098 == 8'h1 ? _GEN_6160 : _GEN_5644; // @[executor.scala 473:84]
  wire [7:0] _GEN_6165 = _GEN_9098 == 8'h1 ? _GEN_6161 : _GEN_5645; // @[executor.scala 473:84]
  wire [7:0] _GEN_6166 = mask_3[0] ? byte_1536 : _GEN_5646; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6167 = mask_3[1] ? byte_1537 : _GEN_5647; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6168 = mask_3[2] ? byte_1538 : _GEN_5648; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6169 = mask_3[3] ? byte_1539 : _GEN_5649; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6170 = _GEN_9098 == 8'h2 ? _GEN_6166 : _GEN_5646; // @[executor.scala 473:84]
  wire [7:0] _GEN_6171 = _GEN_9098 == 8'h2 ? _GEN_6167 : _GEN_5647; // @[executor.scala 473:84]
  wire [7:0] _GEN_6172 = _GEN_9098 == 8'h2 ? _GEN_6168 : _GEN_5648; // @[executor.scala 473:84]
  wire [7:0] _GEN_6173 = _GEN_9098 == 8'h2 ? _GEN_6169 : _GEN_5649; // @[executor.scala 473:84]
  wire [7:0] _GEN_6174 = mask_3[0] ? byte_1536 : _GEN_5650; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6175 = mask_3[1] ? byte_1537 : _GEN_5651; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6176 = mask_3[2] ? byte_1538 : _GEN_5652; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6177 = mask_3[3] ? byte_1539 : _GEN_5653; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6178 = _GEN_9098 == 8'h3 ? _GEN_6174 : _GEN_5650; // @[executor.scala 473:84]
  wire [7:0] _GEN_6179 = _GEN_9098 == 8'h3 ? _GEN_6175 : _GEN_5651; // @[executor.scala 473:84]
  wire [7:0] _GEN_6180 = _GEN_9098 == 8'h3 ? _GEN_6176 : _GEN_5652; // @[executor.scala 473:84]
  wire [7:0] _GEN_6181 = _GEN_9098 == 8'h3 ? _GEN_6177 : _GEN_5653; // @[executor.scala 473:84]
  wire [7:0] _GEN_6182 = mask_3[0] ? byte_1536 : _GEN_5654; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6183 = mask_3[1] ? byte_1537 : _GEN_5655; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6184 = mask_3[2] ? byte_1538 : _GEN_5656; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6185 = mask_3[3] ? byte_1539 : _GEN_5657; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6186 = _GEN_9098 == 8'h4 ? _GEN_6182 : _GEN_5654; // @[executor.scala 473:84]
  wire [7:0] _GEN_6187 = _GEN_9098 == 8'h4 ? _GEN_6183 : _GEN_5655; // @[executor.scala 473:84]
  wire [7:0] _GEN_6188 = _GEN_9098 == 8'h4 ? _GEN_6184 : _GEN_5656; // @[executor.scala 473:84]
  wire [7:0] _GEN_6189 = _GEN_9098 == 8'h4 ? _GEN_6185 : _GEN_5657; // @[executor.scala 473:84]
  wire [7:0] _GEN_6190 = mask_3[0] ? byte_1536 : _GEN_5658; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6191 = mask_3[1] ? byte_1537 : _GEN_5659; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6192 = mask_3[2] ? byte_1538 : _GEN_5660; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6193 = mask_3[3] ? byte_1539 : _GEN_5661; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6194 = _GEN_9098 == 8'h5 ? _GEN_6190 : _GEN_5658; // @[executor.scala 473:84]
  wire [7:0] _GEN_6195 = _GEN_9098 == 8'h5 ? _GEN_6191 : _GEN_5659; // @[executor.scala 473:84]
  wire [7:0] _GEN_6196 = _GEN_9098 == 8'h5 ? _GEN_6192 : _GEN_5660; // @[executor.scala 473:84]
  wire [7:0] _GEN_6197 = _GEN_9098 == 8'h5 ? _GEN_6193 : _GEN_5661; // @[executor.scala 473:84]
  wire [7:0] _GEN_6198 = mask_3[0] ? byte_1536 : _GEN_5662; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6199 = mask_3[1] ? byte_1537 : _GEN_5663; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6200 = mask_3[2] ? byte_1538 : _GEN_5664; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6201 = mask_3[3] ? byte_1539 : _GEN_5665; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6202 = _GEN_9098 == 8'h6 ? _GEN_6198 : _GEN_5662; // @[executor.scala 473:84]
  wire [7:0] _GEN_6203 = _GEN_9098 == 8'h6 ? _GEN_6199 : _GEN_5663; // @[executor.scala 473:84]
  wire [7:0] _GEN_6204 = _GEN_9098 == 8'h6 ? _GEN_6200 : _GEN_5664; // @[executor.scala 473:84]
  wire [7:0] _GEN_6205 = _GEN_9098 == 8'h6 ? _GEN_6201 : _GEN_5665; // @[executor.scala 473:84]
  wire [7:0] _GEN_6206 = mask_3[0] ? byte_1536 : _GEN_5666; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6207 = mask_3[1] ? byte_1537 : _GEN_5667; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6208 = mask_3[2] ? byte_1538 : _GEN_5668; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6209 = mask_3[3] ? byte_1539 : _GEN_5669; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6210 = _GEN_9098 == 8'h7 ? _GEN_6206 : _GEN_5666; // @[executor.scala 473:84]
  wire [7:0] _GEN_6211 = _GEN_9098 == 8'h7 ? _GEN_6207 : _GEN_5667; // @[executor.scala 473:84]
  wire [7:0] _GEN_6212 = _GEN_9098 == 8'h7 ? _GEN_6208 : _GEN_5668; // @[executor.scala 473:84]
  wire [7:0] _GEN_6213 = _GEN_9098 == 8'h7 ? _GEN_6209 : _GEN_5669; // @[executor.scala 473:84]
  wire [7:0] _GEN_6214 = mask_3[0] ? byte_1536 : _GEN_5670; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6215 = mask_3[1] ? byte_1537 : _GEN_5671; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6216 = mask_3[2] ? byte_1538 : _GEN_5672; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6217 = mask_3[3] ? byte_1539 : _GEN_5673; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6218 = _GEN_9098 == 8'h8 ? _GEN_6214 : _GEN_5670; // @[executor.scala 473:84]
  wire [7:0] _GEN_6219 = _GEN_9098 == 8'h8 ? _GEN_6215 : _GEN_5671; // @[executor.scala 473:84]
  wire [7:0] _GEN_6220 = _GEN_9098 == 8'h8 ? _GEN_6216 : _GEN_5672; // @[executor.scala 473:84]
  wire [7:0] _GEN_6221 = _GEN_9098 == 8'h8 ? _GEN_6217 : _GEN_5673; // @[executor.scala 473:84]
  wire [7:0] _GEN_6222 = mask_3[0] ? byte_1536 : _GEN_5674; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6223 = mask_3[1] ? byte_1537 : _GEN_5675; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6224 = mask_3[2] ? byte_1538 : _GEN_5676; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6225 = mask_3[3] ? byte_1539 : _GEN_5677; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6226 = _GEN_9098 == 8'h9 ? _GEN_6222 : _GEN_5674; // @[executor.scala 473:84]
  wire [7:0] _GEN_6227 = _GEN_9098 == 8'h9 ? _GEN_6223 : _GEN_5675; // @[executor.scala 473:84]
  wire [7:0] _GEN_6228 = _GEN_9098 == 8'h9 ? _GEN_6224 : _GEN_5676; // @[executor.scala 473:84]
  wire [7:0] _GEN_6229 = _GEN_9098 == 8'h9 ? _GEN_6225 : _GEN_5677; // @[executor.scala 473:84]
  wire [7:0] _GEN_6230 = mask_3[0] ? byte_1536 : _GEN_5678; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6231 = mask_3[1] ? byte_1537 : _GEN_5679; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6232 = mask_3[2] ? byte_1538 : _GEN_5680; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6233 = mask_3[3] ? byte_1539 : _GEN_5681; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6234 = _GEN_9098 == 8'ha ? _GEN_6230 : _GEN_5678; // @[executor.scala 473:84]
  wire [7:0] _GEN_6235 = _GEN_9098 == 8'ha ? _GEN_6231 : _GEN_5679; // @[executor.scala 473:84]
  wire [7:0] _GEN_6236 = _GEN_9098 == 8'ha ? _GEN_6232 : _GEN_5680; // @[executor.scala 473:84]
  wire [7:0] _GEN_6237 = _GEN_9098 == 8'ha ? _GEN_6233 : _GEN_5681; // @[executor.scala 473:84]
  wire [7:0] _GEN_6238 = mask_3[0] ? byte_1536 : _GEN_5682; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6239 = mask_3[1] ? byte_1537 : _GEN_5683; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6240 = mask_3[2] ? byte_1538 : _GEN_5684; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6241 = mask_3[3] ? byte_1539 : _GEN_5685; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6242 = _GEN_9098 == 8'hb ? _GEN_6238 : _GEN_5682; // @[executor.scala 473:84]
  wire [7:0] _GEN_6243 = _GEN_9098 == 8'hb ? _GEN_6239 : _GEN_5683; // @[executor.scala 473:84]
  wire [7:0] _GEN_6244 = _GEN_9098 == 8'hb ? _GEN_6240 : _GEN_5684; // @[executor.scala 473:84]
  wire [7:0] _GEN_6245 = _GEN_9098 == 8'hb ? _GEN_6241 : _GEN_5685; // @[executor.scala 473:84]
  wire [7:0] _GEN_6246 = mask_3[0] ? byte_1536 : _GEN_5686; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6247 = mask_3[1] ? byte_1537 : _GEN_5687; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6248 = mask_3[2] ? byte_1538 : _GEN_5688; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6249 = mask_3[3] ? byte_1539 : _GEN_5689; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6250 = _GEN_9098 == 8'hc ? _GEN_6246 : _GEN_5686; // @[executor.scala 473:84]
  wire [7:0] _GEN_6251 = _GEN_9098 == 8'hc ? _GEN_6247 : _GEN_5687; // @[executor.scala 473:84]
  wire [7:0] _GEN_6252 = _GEN_9098 == 8'hc ? _GEN_6248 : _GEN_5688; // @[executor.scala 473:84]
  wire [7:0] _GEN_6253 = _GEN_9098 == 8'hc ? _GEN_6249 : _GEN_5689; // @[executor.scala 473:84]
  wire [7:0] _GEN_6254 = mask_3[0] ? byte_1536 : _GEN_5690; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6255 = mask_3[1] ? byte_1537 : _GEN_5691; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6256 = mask_3[2] ? byte_1538 : _GEN_5692; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6257 = mask_3[3] ? byte_1539 : _GEN_5693; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6258 = _GEN_9098 == 8'hd ? _GEN_6254 : _GEN_5690; // @[executor.scala 473:84]
  wire [7:0] _GEN_6259 = _GEN_9098 == 8'hd ? _GEN_6255 : _GEN_5691; // @[executor.scala 473:84]
  wire [7:0] _GEN_6260 = _GEN_9098 == 8'hd ? _GEN_6256 : _GEN_5692; // @[executor.scala 473:84]
  wire [7:0] _GEN_6261 = _GEN_9098 == 8'hd ? _GEN_6257 : _GEN_5693; // @[executor.scala 473:84]
  wire [7:0] _GEN_6262 = mask_3[0] ? byte_1536 : _GEN_5694; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6263 = mask_3[1] ? byte_1537 : _GEN_5695; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6264 = mask_3[2] ? byte_1538 : _GEN_5696; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6265 = mask_3[3] ? byte_1539 : _GEN_5697; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6266 = _GEN_9098 == 8'he ? _GEN_6262 : _GEN_5694; // @[executor.scala 473:84]
  wire [7:0] _GEN_6267 = _GEN_9098 == 8'he ? _GEN_6263 : _GEN_5695; // @[executor.scala 473:84]
  wire [7:0] _GEN_6268 = _GEN_9098 == 8'he ? _GEN_6264 : _GEN_5696; // @[executor.scala 473:84]
  wire [7:0] _GEN_6269 = _GEN_9098 == 8'he ? _GEN_6265 : _GEN_5697; // @[executor.scala 473:84]
  wire [7:0] _GEN_6270 = mask_3[0] ? byte_1536 : _GEN_5698; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6271 = mask_3[1] ? byte_1537 : _GEN_5699; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6272 = mask_3[2] ? byte_1538 : _GEN_5700; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6273 = mask_3[3] ? byte_1539 : _GEN_5701; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6274 = _GEN_9098 == 8'hf ? _GEN_6270 : _GEN_5698; // @[executor.scala 473:84]
  wire [7:0] _GEN_6275 = _GEN_9098 == 8'hf ? _GEN_6271 : _GEN_5699; // @[executor.scala 473:84]
  wire [7:0] _GEN_6276 = _GEN_9098 == 8'hf ? _GEN_6272 : _GEN_5700; // @[executor.scala 473:84]
  wire [7:0] _GEN_6277 = _GEN_9098 == 8'hf ? _GEN_6273 : _GEN_5701; // @[executor.scala 473:84]
  wire [7:0] _GEN_6278 = mask_3[0] ? byte_1536 : _GEN_5702; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6279 = mask_3[1] ? byte_1537 : _GEN_5703; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6280 = mask_3[2] ? byte_1538 : _GEN_5704; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6281 = mask_3[3] ? byte_1539 : _GEN_5705; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6282 = _GEN_9098 == 8'h10 ? _GEN_6278 : _GEN_5702; // @[executor.scala 473:84]
  wire [7:0] _GEN_6283 = _GEN_9098 == 8'h10 ? _GEN_6279 : _GEN_5703; // @[executor.scala 473:84]
  wire [7:0] _GEN_6284 = _GEN_9098 == 8'h10 ? _GEN_6280 : _GEN_5704; // @[executor.scala 473:84]
  wire [7:0] _GEN_6285 = _GEN_9098 == 8'h10 ? _GEN_6281 : _GEN_5705; // @[executor.scala 473:84]
  wire [7:0] _GEN_6286 = mask_3[0] ? byte_1536 : _GEN_5706; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6287 = mask_3[1] ? byte_1537 : _GEN_5707; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6288 = mask_3[2] ? byte_1538 : _GEN_5708; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6289 = mask_3[3] ? byte_1539 : _GEN_5709; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6290 = _GEN_9098 == 8'h11 ? _GEN_6286 : _GEN_5706; // @[executor.scala 473:84]
  wire [7:0] _GEN_6291 = _GEN_9098 == 8'h11 ? _GEN_6287 : _GEN_5707; // @[executor.scala 473:84]
  wire [7:0] _GEN_6292 = _GEN_9098 == 8'h11 ? _GEN_6288 : _GEN_5708; // @[executor.scala 473:84]
  wire [7:0] _GEN_6293 = _GEN_9098 == 8'h11 ? _GEN_6289 : _GEN_5709; // @[executor.scala 473:84]
  wire [7:0] _GEN_6294 = mask_3[0] ? byte_1536 : _GEN_5710; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6295 = mask_3[1] ? byte_1537 : _GEN_5711; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6296 = mask_3[2] ? byte_1538 : _GEN_5712; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6297 = mask_3[3] ? byte_1539 : _GEN_5713; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6298 = _GEN_9098 == 8'h12 ? _GEN_6294 : _GEN_5710; // @[executor.scala 473:84]
  wire [7:0] _GEN_6299 = _GEN_9098 == 8'h12 ? _GEN_6295 : _GEN_5711; // @[executor.scala 473:84]
  wire [7:0] _GEN_6300 = _GEN_9098 == 8'h12 ? _GEN_6296 : _GEN_5712; // @[executor.scala 473:84]
  wire [7:0] _GEN_6301 = _GEN_9098 == 8'h12 ? _GEN_6297 : _GEN_5713; // @[executor.scala 473:84]
  wire [7:0] _GEN_6302 = mask_3[0] ? byte_1536 : _GEN_5714; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6303 = mask_3[1] ? byte_1537 : _GEN_5715; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6304 = mask_3[2] ? byte_1538 : _GEN_5716; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6305 = mask_3[3] ? byte_1539 : _GEN_5717; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6306 = _GEN_9098 == 8'h13 ? _GEN_6302 : _GEN_5714; // @[executor.scala 473:84]
  wire [7:0] _GEN_6307 = _GEN_9098 == 8'h13 ? _GEN_6303 : _GEN_5715; // @[executor.scala 473:84]
  wire [7:0] _GEN_6308 = _GEN_9098 == 8'h13 ? _GEN_6304 : _GEN_5716; // @[executor.scala 473:84]
  wire [7:0] _GEN_6309 = _GEN_9098 == 8'h13 ? _GEN_6305 : _GEN_5717; // @[executor.scala 473:84]
  wire [7:0] _GEN_6310 = mask_3[0] ? byte_1536 : _GEN_5718; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6311 = mask_3[1] ? byte_1537 : _GEN_5719; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6312 = mask_3[2] ? byte_1538 : _GEN_5720; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6313 = mask_3[3] ? byte_1539 : _GEN_5721; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6314 = _GEN_9098 == 8'h14 ? _GEN_6310 : _GEN_5718; // @[executor.scala 473:84]
  wire [7:0] _GEN_6315 = _GEN_9098 == 8'h14 ? _GEN_6311 : _GEN_5719; // @[executor.scala 473:84]
  wire [7:0] _GEN_6316 = _GEN_9098 == 8'h14 ? _GEN_6312 : _GEN_5720; // @[executor.scala 473:84]
  wire [7:0] _GEN_6317 = _GEN_9098 == 8'h14 ? _GEN_6313 : _GEN_5721; // @[executor.scala 473:84]
  wire [7:0] _GEN_6318 = mask_3[0] ? byte_1536 : _GEN_5722; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6319 = mask_3[1] ? byte_1537 : _GEN_5723; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6320 = mask_3[2] ? byte_1538 : _GEN_5724; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6321 = mask_3[3] ? byte_1539 : _GEN_5725; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6322 = _GEN_9098 == 8'h15 ? _GEN_6318 : _GEN_5722; // @[executor.scala 473:84]
  wire [7:0] _GEN_6323 = _GEN_9098 == 8'h15 ? _GEN_6319 : _GEN_5723; // @[executor.scala 473:84]
  wire [7:0] _GEN_6324 = _GEN_9098 == 8'h15 ? _GEN_6320 : _GEN_5724; // @[executor.scala 473:84]
  wire [7:0] _GEN_6325 = _GEN_9098 == 8'h15 ? _GEN_6321 : _GEN_5725; // @[executor.scala 473:84]
  wire [7:0] _GEN_6326 = mask_3[0] ? byte_1536 : _GEN_5726; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6327 = mask_3[1] ? byte_1537 : _GEN_5727; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6328 = mask_3[2] ? byte_1538 : _GEN_5728; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6329 = mask_3[3] ? byte_1539 : _GEN_5729; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6330 = _GEN_9098 == 8'h16 ? _GEN_6326 : _GEN_5726; // @[executor.scala 473:84]
  wire [7:0] _GEN_6331 = _GEN_9098 == 8'h16 ? _GEN_6327 : _GEN_5727; // @[executor.scala 473:84]
  wire [7:0] _GEN_6332 = _GEN_9098 == 8'h16 ? _GEN_6328 : _GEN_5728; // @[executor.scala 473:84]
  wire [7:0] _GEN_6333 = _GEN_9098 == 8'h16 ? _GEN_6329 : _GEN_5729; // @[executor.scala 473:84]
  wire [7:0] _GEN_6334 = mask_3[0] ? byte_1536 : _GEN_5730; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6335 = mask_3[1] ? byte_1537 : _GEN_5731; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6336 = mask_3[2] ? byte_1538 : _GEN_5732; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6337 = mask_3[3] ? byte_1539 : _GEN_5733; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6338 = _GEN_9098 == 8'h17 ? _GEN_6334 : _GEN_5730; // @[executor.scala 473:84]
  wire [7:0] _GEN_6339 = _GEN_9098 == 8'h17 ? _GEN_6335 : _GEN_5731; // @[executor.scala 473:84]
  wire [7:0] _GEN_6340 = _GEN_9098 == 8'h17 ? _GEN_6336 : _GEN_5732; // @[executor.scala 473:84]
  wire [7:0] _GEN_6341 = _GEN_9098 == 8'h17 ? _GEN_6337 : _GEN_5733; // @[executor.scala 473:84]
  wire [7:0] _GEN_6342 = mask_3[0] ? byte_1536 : _GEN_5734; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6343 = mask_3[1] ? byte_1537 : _GEN_5735; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6344 = mask_3[2] ? byte_1538 : _GEN_5736; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6345 = mask_3[3] ? byte_1539 : _GEN_5737; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6346 = _GEN_9098 == 8'h18 ? _GEN_6342 : _GEN_5734; // @[executor.scala 473:84]
  wire [7:0] _GEN_6347 = _GEN_9098 == 8'h18 ? _GEN_6343 : _GEN_5735; // @[executor.scala 473:84]
  wire [7:0] _GEN_6348 = _GEN_9098 == 8'h18 ? _GEN_6344 : _GEN_5736; // @[executor.scala 473:84]
  wire [7:0] _GEN_6349 = _GEN_9098 == 8'h18 ? _GEN_6345 : _GEN_5737; // @[executor.scala 473:84]
  wire [7:0] _GEN_6350 = mask_3[0] ? byte_1536 : _GEN_5738; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6351 = mask_3[1] ? byte_1537 : _GEN_5739; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6352 = mask_3[2] ? byte_1538 : _GEN_5740; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6353 = mask_3[3] ? byte_1539 : _GEN_5741; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6354 = _GEN_9098 == 8'h19 ? _GEN_6350 : _GEN_5738; // @[executor.scala 473:84]
  wire [7:0] _GEN_6355 = _GEN_9098 == 8'h19 ? _GEN_6351 : _GEN_5739; // @[executor.scala 473:84]
  wire [7:0] _GEN_6356 = _GEN_9098 == 8'h19 ? _GEN_6352 : _GEN_5740; // @[executor.scala 473:84]
  wire [7:0] _GEN_6357 = _GEN_9098 == 8'h19 ? _GEN_6353 : _GEN_5741; // @[executor.scala 473:84]
  wire [7:0] _GEN_6358 = mask_3[0] ? byte_1536 : _GEN_5742; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6359 = mask_3[1] ? byte_1537 : _GEN_5743; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6360 = mask_3[2] ? byte_1538 : _GEN_5744; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6361 = mask_3[3] ? byte_1539 : _GEN_5745; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6362 = _GEN_9098 == 8'h1a ? _GEN_6358 : _GEN_5742; // @[executor.scala 473:84]
  wire [7:0] _GEN_6363 = _GEN_9098 == 8'h1a ? _GEN_6359 : _GEN_5743; // @[executor.scala 473:84]
  wire [7:0] _GEN_6364 = _GEN_9098 == 8'h1a ? _GEN_6360 : _GEN_5744; // @[executor.scala 473:84]
  wire [7:0] _GEN_6365 = _GEN_9098 == 8'h1a ? _GEN_6361 : _GEN_5745; // @[executor.scala 473:84]
  wire [7:0] _GEN_6366 = mask_3[0] ? byte_1536 : _GEN_5746; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6367 = mask_3[1] ? byte_1537 : _GEN_5747; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6368 = mask_3[2] ? byte_1538 : _GEN_5748; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6369 = mask_3[3] ? byte_1539 : _GEN_5749; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6370 = _GEN_9098 == 8'h1b ? _GEN_6366 : _GEN_5746; // @[executor.scala 473:84]
  wire [7:0] _GEN_6371 = _GEN_9098 == 8'h1b ? _GEN_6367 : _GEN_5747; // @[executor.scala 473:84]
  wire [7:0] _GEN_6372 = _GEN_9098 == 8'h1b ? _GEN_6368 : _GEN_5748; // @[executor.scala 473:84]
  wire [7:0] _GEN_6373 = _GEN_9098 == 8'h1b ? _GEN_6369 : _GEN_5749; // @[executor.scala 473:84]
  wire [7:0] _GEN_6374 = mask_3[0] ? byte_1536 : _GEN_5750; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6375 = mask_3[1] ? byte_1537 : _GEN_5751; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6376 = mask_3[2] ? byte_1538 : _GEN_5752; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6377 = mask_3[3] ? byte_1539 : _GEN_5753; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6378 = _GEN_9098 == 8'h1c ? _GEN_6374 : _GEN_5750; // @[executor.scala 473:84]
  wire [7:0] _GEN_6379 = _GEN_9098 == 8'h1c ? _GEN_6375 : _GEN_5751; // @[executor.scala 473:84]
  wire [7:0] _GEN_6380 = _GEN_9098 == 8'h1c ? _GEN_6376 : _GEN_5752; // @[executor.scala 473:84]
  wire [7:0] _GEN_6381 = _GEN_9098 == 8'h1c ? _GEN_6377 : _GEN_5753; // @[executor.scala 473:84]
  wire [7:0] _GEN_6382 = mask_3[0] ? byte_1536 : _GEN_5754; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6383 = mask_3[1] ? byte_1537 : _GEN_5755; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6384 = mask_3[2] ? byte_1538 : _GEN_5756; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6385 = mask_3[3] ? byte_1539 : _GEN_5757; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6386 = _GEN_9098 == 8'h1d ? _GEN_6382 : _GEN_5754; // @[executor.scala 473:84]
  wire [7:0] _GEN_6387 = _GEN_9098 == 8'h1d ? _GEN_6383 : _GEN_5755; // @[executor.scala 473:84]
  wire [7:0] _GEN_6388 = _GEN_9098 == 8'h1d ? _GEN_6384 : _GEN_5756; // @[executor.scala 473:84]
  wire [7:0] _GEN_6389 = _GEN_9098 == 8'h1d ? _GEN_6385 : _GEN_5757; // @[executor.scala 473:84]
  wire [7:0] _GEN_6390 = mask_3[0] ? byte_1536 : _GEN_5758; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6391 = mask_3[1] ? byte_1537 : _GEN_5759; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6392 = mask_3[2] ? byte_1538 : _GEN_5760; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6393 = mask_3[3] ? byte_1539 : _GEN_5761; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6394 = _GEN_9098 == 8'h1e ? _GEN_6390 : _GEN_5758; // @[executor.scala 473:84]
  wire [7:0] _GEN_6395 = _GEN_9098 == 8'h1e ? _GEN_6391 : _GEN_5759; // @[executor.scala 473:84]
  wire [7:0] _GEN_6396 = _GEN_9098 == 8'h1e ? _GEN_6392 : _GEN_5760; // @[executor.scala 473:84]
  wire [7:0] _GEN_6397 = _GEN_9098 == 8'h1e ? _GEN_6393 : _GEN_5761; // @[executor.scala 473:84]
  wire [7:0] _GEN_6398 = mask_3[0] ? byte_1536 : _GEN_5762; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6399 = mask_3[1] ? byte_1537 : _GEN_5763; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6400 = mask_3[2] ? byte_1538 : _GEN_5764; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6401 = mask_3[3] ? byte_1539 : _GEN_5765; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6402 = _GEN_9098 == 8'h1f ? _GEN_6398 : _GEN_5762; // @[executor.scala 473:84]
  wire [7:0] _GEN_6403 = _GEN_9098 == 8'h1f ? _GEN_6399 : _GEN_5763; // @[executor.scala 473:84]
  wire [7:0] _GEN_6404 = _GEN_9098 == 8'h1f ? _GEN_6400 : _GEN_5764; // @[executor.scala 473:84]
  wire [7:0] _GEN_6405 = _GEN_9098 == 8'h1f ? _GEN_6401 : _GEN_5765; // @[executor.scala 473:84]
  wire [7:0] _GEN_6406 = mask_3[0] ? byte_1536 : _GEN_5766; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6407 = mask_3[1] ? byte_1537 : _GEN_5767; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6408 = mask_3[2] ? byte_1538 : _GEN_5768; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6409 = mask_3[3] ? byte_1539 : _GEN_5769; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6410 = _GEN_9098 == 8'h20 ? _GEN_6406 : _GEN_5766; // @[executor.scala 473:84]
  wire [7:0] _GEN_6411 = _GEN_9098 == 8'h20 ? _GEN_6407 : _GEN_5767; // @[executor.scala 473:84]
  wire [7:0] _GEN_6412 = _GEN_9098 == 8'h20 ? _GEN_6408 : _GEN_5768; // @[executor.scala 473:84]
  wire [7:0] _GEN_6413 = _GEN_9098 == 8'h20 ? _GEN_6409 : _GEN_5769; // @[executor.scala 473:84]
  wire [7:0] _GEN_6414 = mask_3[0] ? byte_1536 : _GEN_5770; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6415 = mask_3[1] ? byte_1537 : _GEN_5771; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6416 = mask_3[2] ? byte_1538 : _GEN_5772; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6417 = mask_3[3] ? byte_1539 : _GEN_5773; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6418 = _GEN_9098 == 8'h21 ? _GEN_6414 : _GEN_5770; // @[executor.scala 473:84]
  wire [7:0] _GEN_6419 = _GEN_9098 == 8'h21 ? _GEN_6415 : _GEN_5771; // @[executor.scala 473:84]
  wire [7:0] _GEN_6420 = _GEN_9098 == 8'h21 ? _GEN_6416 : _GEN_5772; // @[executor.scala 473:84]
  wire [7:0] _GEN_6421 = _GEN_9098 == 8'h21 ? _GEN_6417 : _GEN_5773; // @[executor.scala 473:84]
  wire [7:0] _GEN_6422 = mask_3[0] ? byte_1536 : _GEN_5774; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6423 = mask_3[1] ? byte_1537 : _GEN_5775; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6424 = mask_3[2] ? byte_1538 : _GEN_5776; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6425 = mask_3[3] ? byte_1539 : _GEN_5777; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6426 = _GEN_9098 == 8'h22 ? _GEN_6422 : _GEN_5774; // @[executor.scala 473:84]
  wire [7:0] _GEN_6427 = _GEN_9098 == 8'h22 ? _GEN_6423 : _GEN_5775; // @[executor.scala 473:84]
  wire [7:0] _GEN_6428 = _GEN_9098 == 8'h22 ? _GEN_6424 : _GEN_5776; // @[executor.scala 473:84]
  wire [7:0] _GEN_6429 = _GEN_9098 == 8'h22 ? _GEN_6425 : _GEN_5777; // @[executor.scala 473:84]
  wire [7:0] _GEN_6430 = mask_3[0] ? byte_1536 : _GEN_5778; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6431 = mask_3[1] ? byte_1537 : _GEN_5779; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6432 = mask_3[2] ? byte_1538 : _GEN_5780; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6433 = mask_3[3] ? byte_1539 : _GEN_5781; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6434 = _GEN_9098 == 8'h23 ? _GEN_6430 : _GEN_5778; // @[executor.scala 473:84]
  wire [7:0] _GEN_6435 = _GEN_9098 == 8'h23 ? _GEN_6431 : _GEN_5779; // @[executor.scala 473:84]
  wire [7:0] _GEN_6436 = _GEN_9098 == 8'h23 ? _GEN_6432 : _GEN_5780; // @[executor.scala 473:84]
  wire [7:0] _GEN_6437 = _GEN_9098 == 8'h23 ? _GEN_6433 : _GEN_5781; // @[executor.scala 473:84]
  wire [7:0] _GEN_6438 = mask_3[0] ? byte_1536 : _GEN_5782; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6439 = mask_3[1] ? byte_1537 : _GEN_5783; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6440 = mask_3[2] ? byte_1538 : _GEN_5784; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6441 = mask_3[3] ? byte_1539 : _GEN_5785; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6442 = _GEN_9098 == 8'h24 ? _GEN_6438 : _GEN_5782; // @[executor.scala 473:84]
  wire [7:0] _GEN_6443 = _GEN_9098 == 8'h24 ? _GEN_6439 : _GEN_5783; // @[executor.scala 473:84]
  wire [7:0] _GEN_6444 = _GEN_9098 == 8'h24 ? _GEN_6440 : _GEN_5784; // @[executor.scala 473:84]
  wire [7:0] _GEN_6445 = _GEN_9098 == 8'h24 ? _GEN_6441 : _GEN_5785; // @[executor.scala 473:84]
  wire [7:0] _GEN_6446 = mask_3[0] ? byte_1536 : _GEN_5786; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6447 = mask_3[1] ? byte_1537 : _GEN_5787; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6448 = mask_3[2] ? byte_1538 : _GEN_5788; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6449 = mask_3[3] ? byte_1539 : _GEN_5789; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6450 = _GEN_9098 == 8'h25 ? _GEN_6446 : _GEN_5786; // @[executor.scala 473:84]
  wire [7:0] _GEN_6451 = _GEN_9098 == 8'h25 ? _GEN_6447 : _GEN_5787; // @[executor.scala 473:84]
  wire [7:0] _GEN_6452 = _GEN_9098 == 8'h25 ? _GEN_6448 : _GEN_5788; // @[executor.scala 473:84]
  wire [7:0] _GEN_6453 = _GEN_9098 == 8'h25 ? _GEN_6449 : _GEN_5789; // @[executor.scala 473:84]
  wire [7:0] _GEN_6454 = mask_3[0] ? byte_1536 : _GEN_5790; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6455 = mask_3[1] ? byte_1537 : _GEN_5791; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6456 = mask_3[2] ? byte_1538 : _GEN_5792; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6457 = mask_3[3] ? byte_1539 : _GEN_5793; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6458 = _GEN_9098 == 8'h26 ? _GEN_6454 : _GEN_5790; // @[executor.scala 473:84]
  wire [7:0] _GEN_6459 = _GEN_9098 == 8'h26 ? _GEN_6455 : _GEN_5791; // @[executor.scala 473:84]
  wire [7:0] _GEN_6460 = _GEN_9098 == 8'h26 ? _GEN_6456 : _GEN_5792; // @[executor.scala 473:84]
  wire [7:0] _GEN_6461 = _GEN_9098 == 8'h26 ? _GEN_6457 : _GEN_5793; // @[executor.scala 473:84]
  wire [7:0] _GEN_6462 = mask_3[0] ? byte_1536 : _GEN_5794; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6463 = mask_3[1] ? byte_1537 : _GEN_5795; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6464 = mask_3[2] ? byte_1538 : _GEN_5796; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6465 = mask_3[3] ? byte_1539 : _GEN_5797; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6466 = _GEN_9098 == 8'h27 ? _GEN_6462 : _GEN_5794; // @[executor.scala 473:84]
  wire [7:0] _GEN_6467 = _GEN_9098 == 8'h27 ? _GEN_6463 : _GEN_5795; // @[executor.scala 473:84]
  wire [7:0] _GEN_6468 = _GEN_9098 == 8'h27 ? _GEN_6464 : _GEN_5796; // @[executor.scala 473:84]
  wire [7:0] _GEN_6469 = _GEN_9098 == 8'h27 ? _GEN_6465 : _GEN_5797; // @[executor.scala 473:84]
  wire [7:0] _GEN_6470 = mask_3[0] ? byte_1536 : _GEN_5798; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6471 = mask_3[1] ? byte_1537 : _GEN_5799; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6472 = mask_3[2] ? byte_1538 : _GEN_5800; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6473 = mask_3[3] ? byte_1539 : _GEN_5801; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6474 = _GEN_9098 == 8'h28 ? _GEN_6470 : _GEN_5798; // @[executor.scala 473:84]
  wire [7:0] _GEN_6475 = _GEN_9098 == 8'h28 ? _GEN_6471 : _GEN_5799; // @[executor.scala 473:84]
  wire [7:0] _GEN_6476 = _GEN_9098 == 8'h28 ? _GEN_6472 : _GEN_5800; // @[executor.scala 473:84]
  wire [7:0] _GEN_6477 = _GEN_9098 == 8'h28 ? _GEN_6473 : _GEN_5801; // @[executor.scala 473:84]
  wire [7:0] _GEN_6478 = mask_3[0] ? byte_1536 : _GEN_5802; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6479 = mask_3[1] ? byte_1537 : _GEN_5803; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6480 = mask_3[2] ? byte_1538 : _GEN_5804; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6481 = mask_3[3] ? byte_1539 : _GEN_5805; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6482 = _GEN_9098 == 8'h29 ? _GEN_6478 : _GEN_5802; // @[executor.scala 473:84]
  wire [7:0] _GEN_6483 = _GEN_9098 == 8'h29 ? _GEN_6479 : _GEN_5803; // @[executor.scala 473:84]
  wire [7:0] _GEN_6484 = _GEN_9098 == 8'h29 ? _GEN_6480 : _GEN_5804; // @[executor.scala 473:84]
  wire [7:0] _GEN_6485 = _GEN_9098 == 8'h29 ? _GEN_6481 : _GEN_5805; // @[executor.scala 473:84]
  wire [7:0] _GEN_6486 = mask_3[0] ? byte_1536 : _GEN_5806; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6487 = mask_3[1] ? byte_1537 : _GEN_5807; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6488 = mask_3[2] ? byte_1538 : _GEN_5808; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6489 = mask_3[3] ? byte_1539 : _GEN_5809; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6490 = _GEN_9098 == 8'h2a ? _GEN_6486 : _GEN_5806; // @[executor.scala 473:84]
  wire [7:0] _GEN_6491 = _GEN_9098 == 8'h2a ? _GEN_6487 : _GEN_5807; // @[executor.scala 473:84]
  wire [7:0] _GEN_6492 = _GEN_9098 == 8'h2a ? _GEN_6488 : _GEN_5808; // @[executor.scala 473:84]
  wire [7:0] _GEN_6493 = _GEN_9098 == 8'h2a ? _GEN_6489 : _GEN_5809; // @[executor.scala 473:84]
  wire [7:0] _GEN_6494 = mask_3[0] ? byte_1536 : _GEN_5810; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6495 = mask_3[1] ? byte_1537 : _GEN_5811; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6496 = mask_3[2] ? byte_1538 : _GEN_5812; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6497 = mask_3[3] ? byte_1539 : _GEN_5813; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6498 = _GEN_9098 == 8'h2b ? _GEN_6494 : _GEN_5810; // @[executor.scala 473:84]
  wire [7:0] _GEN_6499 = _GEN_9098 == 8'h2b ? _GEN_6495 : _GEN_5811; // @[executor.scala 473:84]
  wire [7:0] _GEN_6500 = _GEN_9098 == 8'h2b ? _GEN_6496 : _GEN_5812; // @[executor.scala 473:84]
  wire [7:0] _GEN_6501 = _GEN_9098 == 8'h2b ? _GEN_6497 : _GEN_5813; // @[executor.scala 473:84]
  wire [7:0] _GEN_6502 = mask_3[0] ? byte_1536 : _GEN_5814; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6503 = mask_3[1] ? byte_1537 : _GEN_5815; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6504 = mask_3[2] ? byte_1538 : _GEN_5816; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6505 = mask_3[3] ? byte_1539 : _GEN_5817; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6506 = _GEN_9098 == 8'h2c ? _GEN_6502 : _GEN_5814; // @[executor.scala 473:84]
  wire [7:0] _GEN_6507 = _GEN_9098 == 8'h2c ? _GEN_6503 : _GEN_5815; // @[executor.scala 473:84]
  wire [7:0] _GEN_6508 = _GEN_9098 == 8'h2c ? _GEN_6504 : _GEN_5816; // @[executor.scala 473:84]
  wire [7:0] _GEN_6509 = _GEN_9098 == 8'h2c ? _GEN_6505 : _GEN_5817; // @[executor.scala 473:84]
  wire [7:0] _GEN_6510 = mask_3[0] ? byte_1536 : _GEN_5818; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6511 = mask_3[1] ? byte_1537 : _GEN_5819; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6512 = mask_3[2] ? byte_1538 : _GEN_5820; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6513 = mask_3[3] ? byte_1539 : _GEN_5821; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6514 = _GEN_9098 == 8'h2d ? _GEN_6510 : _GEN_5818; // @[executor.scala 473:84]
  wire [7:0] _GEN_6515 = _GEN_9098 == 8'h2d ? _GEN_6511 : _GEN_5819; // @[executor.scala 473:84]
  wire [7:0] _GEN_6516 = _GEN_9098 == 8'h2d ? _GEN_6512 : _GEN_5820; // @[executor.scala 473:84]
  wire [7:0] _GEN_6517 = _GEN_9098 == 8'h2d ? _GEN_6513 : _GEN_5821; // @[executor.scala 473:84]
  wire [7:0] _GEN_6518 = mask_3[0] ? byte_1536 : _GEN_5822; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6519 = mask_3[1] ? byte_1537 : _GEN_5823; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6520 = mask_3[2] ? byte_1538 : _GEN_5824; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6521 = mask_3[3] ? byte_1539 : _GEN_5825; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6522 = _GEN_9098 == 8'h2e ? _GEN_6518 : _GEN_5822; // @[executor.scala 473:84]
  wire [7:0] _GEN_6523 = _GEN_9098 == 8'h2e ? _GEN_6519 : _GEN_5823; // @[executor.scala 473:84]
  wire [7:0] _GEN_6524 = _GEN_9098 == 8'h2e ? _GEN_6520 : _GEN_5824; // @[executor.scala 473:84]
  wire [7:0] _GEN_6525 = _GEN_9098 == 8'h2e ? _GEN_6521 : _GEN_5825; // @[executor.scala 473:84]
  wire [7:0] _GEN_6526 = mask_3[0] ? byte_1536 : _GEN_5826; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6527 = mask_3[1] ? byte_1537 : _GEN_5827; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6528 = mask_3[2] ? byte_1538 : _GEN_5828; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6529 = mask_3[3] ? byte_1539 : _GEN_5829; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6530 = _GEN_9098 == 8'h2f ? _GEN_6526 : _GEN_5826; // @[executor.scala 473:84]
  wire [7:0] _GEN_6531 = _GEN_9098 == 8'h2f ? _GEN_6527 : _GEN_5827; // @[executor.scala 473:84]
  wire [7:0] _GEN_6532 = _GEN_9098 == 8'h2f ? _GEN_6528 : _GEN_5828; // @[executor.scala 473:84]
  wire [7:0] _GEN_6533 = _GEN_9098 == 8'h2f ? _GEN_6529 : _GEN_5829; // @[executor.scala 473:84]
  wire [7:0] _GEN_6534 = mask_3[0] ? byte_1536 : _GEN_5830; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6535 = mask_3[1] ? byte_1537 : _GEN_5831; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6536 = mask_3[2] ? byte_1538 : _GEN_5832; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6537 = mask_3[3] ? byte_1539 : _GEN_5833; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6538 = _GEN_9098 == 8'h30 ? _GEN_6534 : _GEN_5830; // @[executor.scala 473:84]
  wire [7:0] _GEN_6539 = _GEN_9098 == 8'h30 ? _GEN_6535 : _GEN_5831; // @[executor.scala 473:84]
  wire [7:0] _GEN_6540 = _GEN_9098 == 8'h30 ? _GEN_6536 : _GEN_5832; // @[executor.scala 473:84]
  wire [7:0] _GEN_6541 = _GEN_9098 == 8'h30 ? _GEN_6537 : _GEN_5833; // @[executor.scala 473:84]
  wire [7:0] _GEN_6542 = mask_3[0] ? byte_1536 : _GEN_5834; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6543 = mask_3[1] ? byte_1537 : _GEN_5835; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6544 = mask_3[2] ? byte_1538 : _GEN_5836; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6545 = mask_3[3] ? byte_1539 : _GEN_5837; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6546 = _GEN_9098 == 8'h31 ? _GEN_6542 : _GEN_5834; // @[executor.scala 473:84]
  wire [7:0] _GEN_6547 = _GEN_9098 == 8'h31 ? _GEN_6543 : _GEN_5835; // @[executor.scala 473:84]
  wire [7:0] _GEN_6548 = _GEN_9098 == 8'h31 ? _GEN_6544 : _GEN_5836; // @[executor.scala 473:84]
  wire [7:0] _GEN_6549 = _GEN_9098 == 8'h31 ? _GEN_6545 : _GEN_5837; // @[executor.scala 473:84]
  wire [7:0] _GEN_6550 = mask_3[0] ? byte_1536 : _GEN_5838; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6551 = mask_3[1] ? byte_1537 : _GEN_5839; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6552 = mask_3[2] ? byte_1538 : _GEN_5840; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6553 = mask_3[3] ? byte_1539 : _GEN_5841; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6554 = _GEN_9098 == 8'h32 ? _GEN_6550 : _GEN_5838; // @[executor.scala 473:84]
  wire [7:0] _GEN_6555 = _GEN_9098 == 8'h32 ? _GEN_6551 : _GEN_5839; // @[executor.scala 473:84]
  wire [7:0] _GEN_6556 = _GEN_9098 == 8'h32 ? _GEN_6552 : _GEN_5840; // @[executor.scala 473:84]
  wire [7:0] _GEN_6557 = _GEN_9098 == 8'h32 ? _GEN_6553 : _GEN_5841; // @[executor.scala 473:84]
  wire [7:0] _GEN_6558 = mask_3[0] ? byte_1536 : _GEN_5842; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6559 = mask_3[1] ? byte_1537 : _GEN_5843; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6560 = mask_3[2] ? byte_1538 : _GEN_5844; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6561 = mask_3[3] ? byte_1539 : _GEN_5845; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6562 = _GEN_9098 == 8'h33 ? _GEN_6558 : _GEN_5842; // @[executor.scala 473:84]
  wire [7:0] _GEN_6563 = _GEN_9098 == 8'h33 ? _GEN_6559 : _GEN_5843; // @[executor.scala 473:84]
  wire [7:0] _GEN_6564 = _GEN_9098 == 8'h33 ? _GEN_6560 : _GEN_5844; // @[executor.scala 473:84]
  wire [7:0] _GEN_6565 = _GEN_9098 == 8'h33 ? _GEN_6561 : _GEN_5845; // @[executor.scala 473:84]
  wire [7:0] _GEN_6566 = mask_3[0] ? byte_1536 : _GEN_5846; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6567 = mask_3[1] ? byte_1537 : _GEN_5847; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6568 = mask_3[2] ? byte_1538 : _GEN_5848; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6569 = mask_3[3] ? byte_1539 : _GEN_5849; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6570 = _GEN_9098 == 8'h34 ? _GEN_6566 : _GEN_5846; // @[executor.scala 473:84]
  wire [7:0] _GEN_6571 = _GEN_9098 == 8'h34 ? _GEN_6567 : _GEN_5847; // @[executor.scala 473:84]
  wire [7:0] _GEN_6572 = _GEN_9098 == 8'h34 ? _GEN_6568 : _GEN_5848; // @[executor.scala 473:84]
  wire [7:0] _GEN_6573 = _GEN_9098 == 8'h34 ? _GEN_6569 : _GEN_5849; // @[executor.scala 473:84]
  wire [7:0] _GEN_6574 = mask_3[0] ? byte_1536 : _GEN_5850; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6575 = mask_3[1] ? byte_1537 : _GEN_5851; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6576 = mask_3[2] ? byte_1538 : _GEN_5852; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6577 = mask_3[3] ? byte_1539 : _GEN_5853; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6578 = _GEN_9098 == 8'h35 ? _GEN_6574 : _GEN_5850; // @[executor.scala 473:84]
  wire [7:0] _GEN_6579 = _GEN_9098 == 8'h35 ? _GEN_6575 : _GEN_5851; // @[executor.scala 473:84]
  wire [7:0] _GEN_6580 = _GEN_9098 == 8'h35 ? _GEN_6576 : _GEN_5852; // @[executor.scala 473:84]
  wire [7:0] _GEN_6581 = _GEN_9098 == 8'h35 ? _GEN_6577 : _GEN_5853; // @[executor.scala 473:84]
  wire [7:0] _GEN_6582 = mask_3[0] ? byte_1536 : _GEN_5854; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6583 = mask_3[1] ? byte_1537 : _GEN_5855; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6584 = mask_3[2] ? byte_1538 : _GEN_5856; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6585 = mask_3[3] ? byte_1539 : _GEN_5857; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6586 = _GEN_9098 == 8'h36 ? _GEN_6582 : _GEN_5854; // @[executor.scala 473:84]
  wire [7:0] _GEN_6587 = _GEN_9098 == 8'h36 ? _GEN_6583 : _GEN_5855; // @[executor.scala 473:84]
  wire [7:0] _GEN_6588 = _GEN_9098 == 8'h36 ? _GEN_6584 : _GEN_5856; // @[executor.scala 473:84]
  wire [7:0] _GEN_6589 = _GEN_9098 == 8'h36 ? _GEN_6585 : _GEN_5857; // @[executor.scala 473:84]
  wire [7:0] _GEN_6590 = mask_3[0] ? byte_1536 : _GEN_5858; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6591 = mask_3[1] ? byte_1537 : _GEN_5859; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6592 = mask_3[2] ? byte_1538 : _GEN_5860; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6593 = mask_3[3] ? byte_1539 : _GEN_5861; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6594 = _GEN_9098 == 8'h37 ? _GEN_6590 : _GEN_5858; // @[executor.scala 473:84]
  wire [7:0] _GEN_6595 = _GEN_9098 == 8'h37 ? _GEN_6591 : _GEN_5859; // @[executor.scala 473:84]
  wire [7:0] _GEN_6596 = _GEN_9098 == 8'h37 ? _GEN_6592 : _GEN_5860; // @[executor.scala 473:84]
  wire [7:0] _GEN_6597 = _GEN_9098 == 8'h37 ? _GEN_6593 : _GEN_5861; // @[executor.scala 473:84]
  wire [7:0] _GEN_6598 = mask_3[0] ? byte_1536 : _GEN_5862; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6599 = mask_3[1] ? byte_1537 : _GEN_5863; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6600 = mask_3[2] ? byte_1538 : _GEN_5864; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6601 = mask_3[3] ? byte_1539 : _GEN_5865; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6602 = _GEN_9098 == 8'h38 ? _GEN_6598 : _GEN_5862; // @[executor.scala 473:84]
  wire [7:0] _GEN_6603 = _GEN_9098 == 8'h38 ? _GEN_6599 : _GEN_5863; // @[executor.scala 473:84]
  wire [7:0] _GEN_6604 = _GEN_9098 == 8'h38 ? _GEN_6600 : _GEN_5864; // @[executor.scala 473:84]
  wire [7:0] _GEN_6605 = _GEN_9098 == 8'h38 ? _GEN_6601 : _GEN_5865; // @[executor.scala 473:84]
  wire [7:0] _GEN_6606 = mask_3[0] ? byte_1536 : _GEN_5866; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6607 = mask_3[1] ? byte_1537 : _GEN_5867; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6608 = mask_3[2] ? byte_1538 : _GEN_5868; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6609 = mask_3[3] ? byte_1539 : _GEN_5869; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6610 = _GEN_9098 == 8'h39 ? _GEN_6606 : _GEN_5866; // @[executor.scala 473:84]
  wire [7:0] _GEN_6611 = _GEN_9098 == 8'h39 ? _GEN_6607 : _GEN_5867; // @[executor.scala 473:84]
  wire [7:0] _GEN_6612 = _GEN_9098 == 8'h39 ? _GEN_6608 : _GEN_5868; // @[executor.scala 473:84]
  wire [7:0] _GEN_6613 = _GEN_9098 == 8'h39 ? _GEN_6609 : _GEN_5869; // @[executor.scala 473:84]
  wire [7:0] _GEN_6614 = mask_3[0] ? byte_1536 : _GEN_5870; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6615 = mask_3[1] ? byte_1537 : _GEN_5871; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6616 = mask_3[2] ? byte_1538 : _GEN_5872; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6617 = mask_3[3] ? byte_1539 : _GEN_5873; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6618 = _GEN_9098 == 8'h3a ? _GEN_6614 : _GEN_5870; // @[executor.scala 473:84]
  wire [7:0] _GEN_6619 = _GEN_9098 == 8'h3a ? _GEN_6615 : _GEN_5871; // @[executor.scala 473:84]
  wire [7:0] _GEN_6620 = _GEN_9098 == 8'h3a ? _GEN_6616 : _GEN_5872; // @[executor.scala 473:84]
  wire [7:0] _GEN_6621 = _GEN_9098 == 8'h3a ? _GEN_6617 : _GEN_5873; // @[executor.scala 473:84]
  wire [7:0] _GEN_6622 = mask_3[0] ? byte_1536 : _GEN_5874; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6623 = mask_3[1] ? byte_1537 : _GEN_5875; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6624 = mask_3[2] ? byte_1538 : _GEN_5876; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6625 = mask_3[3] ? byte_1539 : _GEN_5877; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6626 = _GEN_9098 == 8'h3b ? _GEN_6622 : _GEN_5874; // @[executor.scala 473:84]
  wire [7:0] _GEN_6627 = _GEN_9098 == 8'h3b ? _GEN_6623 : _GEN_5875; // @[executor.scala 473:84]
  wire [7:0] _GEN_6628 = _GEN_9098 == 8'h3b ? _GEN_6624 : _GEN_5876; // @[executor.scala 473:84]
  wire [7:0] _GEN_6629 = _GEN_9098 == 8'h3b ? _GEN_6625 : _GEN_5877; // @[executor.scala 473:84]
  wire [7:0] _GEN_6630 = mask_3[0] ? byte_1536 : _GEN_5878; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6631 = mask_3[1] ? byte_1537 : _GEN_5879; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6632 = mask_3[2] ? byte_1538 : _GEN_5880; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6633 = mask_3[3] ? byte_1539 : _GEN_5881; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6634 = _GEN_9098 == 8'h3c ? _GEN_6630 : _GEN_5878; // @[executor.scala 473:84]
  wire [7:0] _GEN_6635 = _GEN_9098 == 8'h3c ? _GEN_6631 : _GEN_5879; // @[executor.scala 473:84]
  wire [7:0] _GEN_6636 = _GEN_9098 == 8'h3c ? _GEN_6632 : _GEN_5880; // @[executor.scala 473:84]
  wire [7:0] _GEN_6637 = _GEN_9098 == 8'h3c ? _GEN_6633 : _GEN_5881; // @[executor.scala 473:84]
  wire [7:0] _GEN_6638 = mask_3[0] ? byte_1536 : _GEN_5882; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6639 = mask_3[1] ? byte_1537 : _GEN_5883; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6640 = mask_3[2] ? byte_1538 : _GEN_5884; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6641 = mask_3[3] ? byte_1539 : _GEN_5885; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6642 = _GEN_9098 == 8'h3d ? _GEN_6638 : _GEN_5882; // @[executor.scala 473:84]
  wire [7:0] _GEN_6643 = _GEN_9098 == 8'h3d ? _GEN_6639 : _GEN_5883; // @[executor.scala 473:84]
  wire [7:0] _GEN_6644 = _GEN_9098 == 8'h3d ? _GEN_6640 : _GEN_5884; // @[executor.scala 473:84]
  wire [7:0] _GEN_6645 = _GEN_9098 == 8'h3d ? _GEN_6641 : _GEN_5885; // @[executor.scala 473:84]
  wire [7:0] _GEN_6646 = mask_3[0] ? byte_1536 : _GEN_5886; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6647 = mask_3[1] ? byte_1537 : _GEN_5887; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6648 = mask_3[2] ? byte_1538 : _GEN_5888; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6649 = mask_3[3] ? byte_1539 : _GEN_5889; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6650 = _GEN_9098 == 8'h3e ? _GEN_6646 : _GEN_5886; // @[executor.scala 473:84]
  wire [7:0] _GEN_6651 = _GEN_9098 == 8'h3e ? _GEN_6647 : _GEN_5887; // @[executor.scala 473:84]
  wire [7:0] _GEN_6652 = _GEN_9098 == 8'h3e ? _GEN_6648 : _GEN_5888; // @[executor.scala 473:84]
  wire [7:0] _GEN_6653 = _GEN_9098 == 8'h3e ? _GEN_6649 : _GEN_5889; // @[executor.scala 473:84]
  wire [7:0] _GEN_6654 = mask_3[0] ? byte_1536 : _GEN_5890; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6655 = mask_3[1] ? byte_1537 : _GEN_5891; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6656 = mask_3[2] ? byte_1538 : _GEN_5892; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6657 = mask_3[3] ? byte_1539 : _GEN_5893; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6658 = _GEN_9098 == 8'h3f ? _GEN_6654 : _GEN_5890; // @[executor.scala 473:84]
  wire [7:0] _GEN_6659 = _GEN_9098 == 8'h3f ? _GEN_6655 : _GEN_5891; // @[executor.scala 473:84]
  wire [7:0] _GEN_6660 = _GEN_9098 == 8'h3f ? _GEN_6656 : _GEN_5892; // @[executor.scala 473:84]
  wire [7:0] _GEN_6661 = _GEN_9098 == 8'h3f ? _GEN_6657 : _GEN_5893; // @[executor.scala 473:84]
  wire [7:0] _GEN_6662 = mask_3[0] ? byte_1536 : _GEN_5894; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6663 = mask_3[1] ? byte_1537 : _GEN_5895; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6664 = mask_3[2] ? byte_1538 : _GEN_5896; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6665 = mask_3[3] ? byte_1539 : _GEN_5897; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6666 = _GEN_9098 == 8'h40 ? _GEN_6662 : _GEN_5894; // @[executor.scala 473:84]
  wire [7:0] _GEN_6667 = _GEN_9098 == 8'h40 ? _GEN_6663 : _GEN_5895; // @[executor.scala 473:84]
  wire [7:0] _GEN_6668 = _GEN_9098 == 8'h40 ? _GEN_6664 : _GEN_5896; // @[executor.scala 473:84]
  wire [7:0] _GEN_6669 = _GEN_9098 == 8'h40 ? _GEN_6665 : _GEN_5897; // @[executor.scala 473:84]
  wire [7:0] _GEN_6670 = mask_3[0] ? byte_1536 : _GEN_5898; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6671 = mask_3[1] ? byte_1537 : _GEN_5899; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6672 = mask_3[2] ? byte_1538 : _GEN_5900; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6673 = mask_3[3] ? byte_1539 : _GEN_5901; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6674 = _GEN_9098 == 8'h41 ? _GEN_6670 : _GEN_5898; // @[executor.scala 473:84]
  wire [7:0] _GEN_6675 = _GEN_9098 == 8'h41 ? _GEN_6671 : _GEN_5899; // @[executor.scala 473:84]
  wire [7:0] _GEN_6676 = _GEN_9098 == 8'h41 ? _GEN_6672 : _GEN_5900; // @[executor.scala 473:84]
  wire [7:0] _GEN_6677 = _GEN_9098 == 8'h41 ? _GEN_6673 : _GEN_5901; // @[executor.scala 473:84]
  wire [7:0] _GEN_6678 = mask_3[0] ? byte_1536 : _GEN_5902; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6679 = mask_3[1] ? byte_1537 : _GEN_5903; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6680 = mask_3[2] ? byte_1538 : _GEN_5904; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6681 = mask_3[3] ? byte_1539 : _GEN_5905; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6682 = _GEN_9098 == 8'h42 ? _GEN_6678 : _GEN_5902; // @[executor.scala 473:84]
  wire [7:0] _GEN_6683 = _GEN_9098 == 8'h42 ? _GEN_6679 : _GEN_5903; // @[executor.scala 473:84]
  wire [7:0] _GEN_6684 = _GEN_9098 == 8'h42 ? _GEN_6680 : _GEN_5904; // @[executor.scala 473:84]
  wire [7:0] _GEN_6685 = _GEN_9098 == 8'h42 ? _GEN_6681 : _GEN_5905; // @[executor.scala 473:84]
  wire [7:0] _GEN_6686 = mask_3[0] ? byte_1536 : _GEN_5906; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6687 = mask_3[1] ? byte_1537 : _GEN_5907; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6688 = mask_3[2] ? byte_1538 : _GEN_5908; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6689 = mask_3[3] ? byte_1539 : _GEN_5909; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6690 = _GEN_9098 == 8'h43 ? _GEN_6686 : _GEN_5906; // @[executor.scala 473:84]
  wire [7:0] _GEN_6691 = _GEN_9098 == 8'h43 ? _GEN_6687 : _GEN_5907; // @[executor.scala 473:84]
  wire [7:0] _GEN_6692 = _GEN_9098 == 8'h43 ? _GEN_6688 : _GEN_5908; // @[executor.scala 473:84]
  wire [7:0] _GEN_6693 = _GEN_9098 == 8'h43 ? _GEN_6689 : _GEN_5909; // @[executor.scala 473:84]
  wire [7:0] _GEN_6694 = mask_3[0] ? byte_1536 : _GEN_5910; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6695 = mask_3[1] ? byte_1537 : _GEN_5911; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6696 = mask_3[2] ? byte_1538 : _GEN_5912; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6697 = mask_3[3] ? byte_1539 : _GEN_5913; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6698 = _GEN_9098 == 8'h44 ? _GEN_6694 : _GEN_5910; // @[executor.scala 473:84]
  wire [7:0] _GEN_6699 = _GEN_9098 == 8'h44 ? _GEN_6695 : _GEN_5911; // @[executor.scala 473:84]
  wire [7:0] _GEN_6700 = _GEN_9098 == 8'h44 ? _GEN_6696 : _GEN_5912; // @[executor.scala 473:84]
  wire [7:0] _GEN_6701 = _GEN_9098 == 8'h44 ? _GEN_6697 : _GEN_5913; // @[executor.scala 473:84]
  wire [7:0] _GEN_6702 = mask_3[0] ? byte_1536 : _GEN_5914; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6703 = mask_3[1] ? byte_1537 : _GEN_5915; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6704 = mask_3[2] ? byte_1538 : _GEN_5916; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6705 = mask_3[3] ? byte_1539 : _GEN_5917; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6706 = _GEN_9098 == 8'h45 ? _GEN_6702 : _GEN_5914; // @[executor.scala 473:84]
  wire [7:0] _GEN_6707 = _GEN_9098 == 8'h45 ? _GEN_6703 : _GEN_5915; // @[executor.scala 473:84]
  wire [7:0] _GEN_6708 = _GEN_9098 == 8'h45 ? _GEN_6704 : _GEN_5916; // @[executor.scala 473:84]
  wire [7:0] _GEN_6709 = _GEN_9098 == 8'h45 ? _GEN_6705 : _GEN_5917; // @[executor.scala 473:84]
  wire [7:0] _GEN_6710 = mask_3[0] ? byte_1536 : _GEN_5918; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6711 = mask_3[1] ? byte_1537 : _GEN_5919; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6712 = mask_3[2] ? byte_1538 : _GEN_5920; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6713 = mask_3[3] ? byte_1539 : _GEN_5921; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6714 = _GEN_9098 == 8'h46 ? _GEN_6710 : _GEN_5918; // @[executor.scala 473:84]
  wire [7:0] _GEN_6715 = _GEN_9098 == 8'h46 ? _GEN_6711 : _GEN_5919; // @[executor.scala 473:84]
  wire [7:0] _GEN_6716 = _GEN_9098 == 8'h46 ? _GEN_6712 : _GEN_5920; // @[executor.scala 473:84]
  wire [7:0] _GEN_6717 = _GEN_9098 == 8'h46 ? _GEN_6713 : _GEN_5921; // @[executor.scala 473:84]
  wire [7:0] _GEN_6718 = mask_3[0] ? byte_1536 : _GEN_5922; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6719 = mask_3[1] ? byte_1537 : _GEN_5923; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6720 = mask_3[2] ? byte_1538 : _GEN_5924; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6721 = mask_3[3] ? byte_1539 : _GEN_5925; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6722 = _GEN_9098 == 8'h47 ? _GEN_6718 : _GEN_5922; // @[executor.scala 473:84]
  wire [7:0] _GEN_6723 = _GEN_9098 == 8'h47 ? _GEN_6719 : _GEN_5923; // @[executor.scala 473:84]
  wire [7:0] _GEN_6724 = _GEN_9098 == 8'h47 ? _GEN_6720 : _GEN_5924; // @[executor.scala 473:84]
  wire [7:0] _GEN_6725 = _GEN_9098 == 8'h47 ? _GEN_6721 : _GEN_5925; // @[executor.scala 473:84]
  wire [7:0] _GEN_6726 = mask_3[0] ? byte_1536 : _GEN_5926; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6727 = mask_3[1] ? byte_1537 : _GEN_5927; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6728 = mask_3[2] ? byte_1538 : _GEN_5928; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6729 = mask_3[3] ? byte_1539 : _GEN_5929; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6730 = _GEN_9098 == 8'h48 ? _GEN_6726 : _GEN_5926; // @[executor.scala 473:84]
  wire [7:0] _GEN_6731 = _GEN_9098 == 8'h48 ? _GEN_6727 : _GEN_5927; // @[executor.scala 473:84]
  wire [7:0] _GEN_6732 = _GEN_9098 == 8'h48 ? _GEN_6728 : _GEN_5928; // @[executor.scala 473:84]
  wire [7:0] _GEN_6733 = _GEN_9098 == 8'h48 ? _GEN_6729 : _GEN_5929; // @[executor.scala 473:84]
  wire [7:0] _GEN_6734 = mask_3[0] ? byte_1536 : _GEN_5930; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6735 = mask_3[1] ? byte_1537 : _GEN_5931; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6736 = mask_3[2] ? byte_1538 : _GEN_5932; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6737 = mask_3[3] ? byte_1539 : _GEN_5933; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6738 = _GEN_9098 == 8'h49 ? _GEN_6734 : _GEN_5930; // @[executor.scala 473:84]
  wire [7:0] _GEN_6739 = _GEN_9098 == 8'h49 ? _GEN_6735 : _GEN_5931; // @[executor.scala 473:84]
  wire [7:0] _GEN_6740 = _GEN_9098 == 8'h49 ? _GEN_6736 : _GEN_5932; // @[executor.scala 473:84]
  wire [7:0] _GEN_6741 = _GEN_9098 == 8'h49 ? _GEN_6737 : _GEN_5933; // @[executor.scala 473:84]
  wire [7:0] _GEN_6742 = mask_3[0] ? byte_1536 : _GEN_5934; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6743 = mask_3[1] ? byte_1537 : _GEN_5935; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6744 = mask_3[2] ? byte_1538 : _GEN_5936; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6745 = mask_3[3] ? byte_1539 : _GEN_5937; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6746 = _GEN_9098 == 8'h4a ? _GEN_6742 : _GEN_5934; // @[executor.scala 473:84]
  wire [7:0] _GEN_6747 = _GEN_9098 == 8'h4a ? _GEN_6743 : _GEN_5935; // @[executor.scala 473:84]
  wire [7:0] _GEN_6748 = _GEN_9098 == 8'h4a ? _GEN_6744 : _GEN_5936; // @[executor.scala 473:84]
  wire [7:0] _GEN_6749 = _GEN_9098 == 8'h4a ? _GEN_6745 : _GEN_5937; // @[executor.scala 473:84]
  wire [7:0] _GEN_6750 = mask_3[0] ? byte_1536 : _GEN_5938; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6751 = mask_3[1] ? byte_1537 : _GEN_5939; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6752 = mask_3[2] ? byte_1538 : _GEN_5940; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6753 = mask_3[3] ? byte_1539 : _GEN_5941; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6754 = _GEN_9098 == 8'h4b ? _GEN_6750 : _GEN_5938; // @[executor.scala 473:84]
  wire [7:0] _GEN_6755 = _GEN_9098 == 8'h4b ? _GEN_6751 : _GEN_5939; // @[executor.scala 473:84]
  wire [7:0] _GEN_6756 = _GEN_9098 == 8'h4b ? _GEN_6752 : _GEN_5940; // @[executor.scala 473:84]
  wire [7:0] _GEN_6757 = _GEN_9098 == 8'h4b ? _GEN_6753 : _GEN_5941; // @[executor.scala 473:84]
  wire [7:0] _GEN_6758 = mask_3[0] ? byte_1536 : _GEN_5942; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6759 = mask_3[1] ? byte_1537 : _GEN_5943; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6760 = mask_3[2] ? byte_1538 : _GEN_5944; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6761 = mask_3[3] ? byte_1539 : _GEN_5945; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6762 = _GEN_9098 == 8'h4c ? _GEN_6758 : _GEN_5942; // @[executor.scala 473:84]
  wire [7:0] _GEN_6763 = _GEN_9098 == 8'h4c ? _GEN_6759 : _GEN_5943; // @[executor.scala 473:84]
  wire [7:0] _GEN_6764 = _GEN_9098 == 8'h4c ? _GEN_6760 : _GEN_5944; // @[executor.scala 473:84]
  wire [7:0] _GEN_6765 = _GEN_9098 == 8'h4c ? _GEN_6761 : _GEN_5945; // @[executor.scala 473:84]
  wire [7:0] _GEN_6766 = mask_3[0] ? byte_1536 : _GEN_5946; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6767 = mask_3[1] ? byte_1537 : _GEN_5947; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6768 = mask_3[2] ? byte_1538 : _GEN_5948; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6769 = mask_3[3] ? byte_1539 : _GEN_5949; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6770 = _GEN_9098 == 8'h4d ? _GEN_6766 : _GEN_5946; // @[executor.scala 473:84]
  wire [7:0] _GEN_6771 = _GEN_9098 == 8'h4d ? _GEN_6767 : _GEN_5947; // @[executor.scala 473:84]
  wire [7:0] _GEN_6772 = _GEN_9098 == 8'h4d ? _GEN_6768 : _GEN_5948; // @[executor.scala 473:84]
  wire [7:0] _GEN_6773 = _GEN_9098 == 8'h4d ? _GEN_6769 : _GEN_5949; // @[executor.scala 473:84]
  wire [7:0] _GEN_6774 = mask_3[0] ? byte_1536 : _GEN_5950; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6775 = mask_3[1] ? byte_1537 : _GEN_5951; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6776 = mask_3[2] ? byte_1538 : _GEN_5952; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6777 = mask_3[3] ? byte_1539 : _GEN_5953; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6778 = _GEN_9098 == 8'h4e ? _GEN_6774 : _GEN_5950; // @[executor.scala 473:84]
  wire [7:0] _GEN_6779 = _GEN_9098 == 8'h4e ? _GEN_6775 : _GEN_5951; // @[executor.scala 473:84]
  wire [7:0] _GEN_6780 = _GEN_9098 == 8'h4e ? _GEN_6776 : _GEN_5952; // @[executor.scala 473:84]
  wire [7:0] _GEN_6781 = _GEN_9098 == 8'h4e ? _GEN_6777 : _GEN_5953; // @[executor.scala 473:84]
  wire [7:0] _GEN_6782 = mask_3[0] ? byte_1536 : _GEN_5954; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6783 = mask_3[1] ? byte_1537 : _GEN_5955; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6784 = mask_3[2] ? byte_1538 : _GEN_5956; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6785 = mask_3[3] ? byte_1539 : _GEN_5957; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6786 = _GEN_9098 == 8'h4f ? _GEN_6782 : _GEN_5954; // @[executor.scala 473:84]
  wire [7:0] _GEN_6787 = _GEN_9098 == 8'h4f ? _GEN_6783 : _GEN_5955; // @[executor.scala 473:84]
  wire [7:0] _GEN_6788 = _GEN_9098 == 8'h4f ? _GEN_6784 : _GEN_5956; // @[executor.scala 473:84]
  wire [7:0] _GEN_6789 = _GEN_9098 == 8'h4f ? _GEN_6785 : _GEN_5957; // @[executor.scala 473:84]
  wire [7:0] _GEN_6790 = mask_3[0] ? byte_1536 : _GEN_5958; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6791 = mask_3[1] ? byte_1537 : _GEN_5959; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6792 = mask_3[2] ? byte_1538 : _GEN_5960; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6793 = mask_3[3] ? byte_1539 : _GEN_5961; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6794 = _GEN_9098 == 8'h50 ? _GEN_6790 : _GEN_5958; // @[executor.scala 473:84]
  wire [7:0] _GEN_6795 = _GEN_9098 == 8'h50 ? _GEN_6791 : _GEN_5959; // @[executor.scala 473:84]
  wire [7:0] _GEN_6796 = _GEN_9098 == 8'h50 ? _GEN_6792 : _GEN_5960; // @[executor.scala 473:84]
  wire [7:0] _GEN_6797 = _GEN_9098 == 8'h50 ? _GEN_6793 : _GEN_5961; // @[executor.scala 473:84]
  wire [7:0] _GEN_6798 = mask_3[0] ? byte_1536 : _GEN_5962; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6799 = mask_3[1] ? byte_1537 : _GEN_5963; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6800 = mask_3[2] ? byte_1538 : _GEN_5964; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6801 = mask_3[3] ? byte_1539 : _GEN_5965; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6802 = _GEN_9098 == 8'h51 ? _GEN_6798 : _GEN_5962; // @[executor.scala 473:84]
  wire [7:0] _GEN_6803 = _GEN_9098 == 8'h51 ? _GEN_6799 : _GEN_5963; // @[executor.scala 473:84]
  wire [7:0] _GEN_6804 = _GEN_9098 == 8'h51 ? _GEN_6800 : _GEN_5964; // @[executor.scala 473:84]
  wire [7:0] _GEN_6805 = _GEN_9098 == 8'h51 ? _GEN_6801 : _GEN_5965; // @[executor.scala 473:84]
  wire [7:0] _GEN_6806 = mask_3[0] ? byte_1536 : _GEN_5966; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6807 = mask_3[1] ? byte_1537 : _GEN_5967; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6808 = mask_3[2] ? byte_1538 : _GEN_5968; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6809 = mask_3[3] ? byte_1539 : _GEN_5969; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6810 = _GEN_9098 == 8'h52 ? _GEN_6806 : _GEN_5966; // @[executor.scala 473:84]
  wire [7:0] _GEN_6811 = _GEN_9098 == 8'h52 ? _GEN_6807 : _GEN_5967; // @[executor.scala 473:84]
  wire [7:0] _GEN_6812 = _GEN_9098 == 8'h52 ? _GEN_6808 : _GEN_5968; // @[executor.scala 473:84]
  wire [7:0] _GEN_6813 = _GEN_9098 == 8'h52 ? _GEN_6809 : _GEN_5969; // @[executor.scala 473:84]
  wire [7:0] _GEN_6814 = mask_3[0] ? byte_1536 : _GEN_5970; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6815 = mask_3[1] ? byte_1537 : _GEN_5971; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6816 = mask_3[2] ? byte_1538 : _GEN_5972; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6817 = mask_3[3] ? byte_1539 : _GEN_5973; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6818 = _GEN_9098 == 8'h53 ? _GEN_6814 : _GEN_5970; // @[executor.scala 473:84]
  wire [7:0] _GEN_6819 = _GEN_9098 == 8'h53 ? _GEN_6815 : _GEN_5971; // @[executor.scala 473:84]
  wire [7:0] _GEN_6820 = _GEN_9098 == 8'h53 ? _GEN_6816 : _GEN_5972; // @[executor.scala 473:84]
  wire [7:0] _GEN_6821 = _GEN_9098 == 8'h53 ? _GEN_6817 : _GEN_5973; // @[executor.scala 473:84]
  wire [7:0] _GEN_6822 = mask_3[0] ? byte_1536 : _GEN_5974; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6823 = mask_3[1] ? byte_1537 : _GEN_5975; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6824 = mask_3[2] ? byte_1538 : _GEN_5976; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6825 = mask_3[3] ? byte_1539 : _GEN_5977; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6826 = _GEN_9098 == 8'h54 ? _GEN_6822 : _GEN_5974; // @[executor.scala 473:84]
  wire [7:0] _GEN_6827 = _GEN_9098 == 8'h54 ? _GEN_6823 : _GEN_5975; // @[executor.scala 473:84]
  wire [7:0] _GEN_6828 = _GEN_9098 == 8'h54 ? _GEN_6824 : _GEN_5976; // @[executor.scala 473:84]
  wire [7:0] _GEN_6829 = _GEN_9098 == 8'h54 ? _GEN_6825 : _GEN_5977; // @[executor.scala 473:84]
  wire [7:0] _GEN_6830 = mask_3[0] ? byte_1536 : _GEN_5978; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6831 = mask_3[1] ? byte_1537 : _GEN_5979; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6832 = mask_3[2] ? byte_1538 : _GEN_5980; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6833 = mask_3[3] ? byte_1539 : _GEN_5981; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6834 = _GEN_9098 == 8'h55 ? _GEN_6830 : _GEN_5978; // @[executor.scala 473:84]
  wire [7:0] _GEN_6835 = _GEN_9098 == 8'h55 ? _GEN_6831 : _GEN_5979; // @[executor.scala 473:84]
  wire [7:0] _GEN_6836 = _GEN_9098 == 8'h55 ? _GEN_6832 : _GEN_5980; // @[executor.scala 473:84]
  wire [7:0] _GEN_6837 = _GEN_9098 == 8'h55 ? _GEN_6833 : _GEN_5981; // @[executor.scala 473:84]
  wire [7:0] _GEN_6838 = mask_3[0] ? byte_1536 : _GEN_5982; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6839 = mask_3[1] ? byte_1537 : _GEN_5983; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6840 = mask_3[2] ? byte_1538 : _GEN_5984; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6841 = mask_3[3] ? byte_1539 : _GEN_5985; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6842 = _GEN_9098 == 8'h56 ? _GEN_6838 : _GEN_5982; // @[executor.scala 473:84]
  wire [7:0] _GEN_6843 = _GEN_9098 == 8'h56 ? _GEN_6839 : _GEN_5983; // @[executor.scala 473:84]
  wire [7:0] _GEN_6844 = _GEN_9098 == 8'h56 ? _GEN_6840 : _GEN_5984; // @[executor.scala 473:84]
  wire [7:0] _GEN_6845 = _GEN_9098 == 8'h56 ? _GEN_6841 : _GEN_5985; // @[executor.scala 473:84]
  wire [7:0] _GEN_6846 = mask_3[0] ? byte_1536 : _GEN_5986; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6847 = mask_3[1] ? byte_1537 : _GEN_5987; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6848 = mask_3[2] ? byte_1538 : _GEN_5988; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6849 = mask_3[3] ? byte_1539 : _GEN_5989; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6850 = _GEN_9098 == 8'h57 ? _GEN_6846 : _GEN_5986; // @[executor.scala 473:84]
  wire [7:0] _GEN_6851 = _GEN_9098 == 8'h57 ? _GEN_6847 : _GEN_5987; // @[executor.scala 473:84]
  wire [7:0] _GEN_6852 = _GEN_9098 == 8'h57 ? _GEN_6848 : _GEN_5988; // @[executor.scala 473:84]
  wire [7:0] _GEN_6853 = _GEN_9098 == 8'h57 ? _GEN_6849 : _GEN_5989; // @[executor.scala 473:84]
  wire [7:0] _GEN_6854 = mask_3[0] ? byte_1536 : _GEN_5990; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6855 = mask_3[1] ? byte_1537 : _GEN_5991; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6856 = mask_3[2] ? byte_1538 : _GEN_5992; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6857 = mask_3[3] ? byte_1539 : _GEN_5993; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6858 = _GEN_9098 == 8'h58 ? _GEN_6854 : _GEN_5990; // @[executor.scala 473:84]
  wire [7:0] _GEN_6859 = _GEN_9098 == 8'h58 ? _GEN_6855 : _GEN_5991; // @[executor.scala 473:84]
  wire [7:0] _GEN_6860 = _GEN_9098 == 8'h58 ? _GEN_6856 : _GEN_5992; // @[executor.scala 473:84]
  wire [7:0] _GEN_6861 = _GEN_9098 == 8'h58 ? _GEN_6857 : _GEN_5993; // @[executor.scala 473:84]
  wire [7:0] _GEN_6862 = mask_3[0] ? byte_1536 : _GEN_5994; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6863 = mask_3[1] ? byte_1537 : _GEN_5995; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6864 = mask_3[2] ? byte_1538 : _GEN_5996; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6865 = mask_3[3] ? byte_1539 : _GEN_5997; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6866 = _GEN_9098 == 8'h59 ? _GEN_6862 : _GEN_5994; // @[executor.scala 473:84]
  wire [7:0] _GEN_6867 = _GEN_9098 == 8'h59 ? _GEN_6863 : _GEN_5995; // @[executor.scala 473:84]
  wire [7:0] _GEN_6868 = _GEN_9098 == 8'h59 ? _GEN_6864 : _GEN_5996; // @[executor.scala 473:84]
  wire [7:0] _GEN_6869 = _GEN_9098 == 8'h59 ? _GEN_6865 : _GEN_5997; // @[executor.scala 473:84]
  wire [7:0] _GEN_6870 = mask_3[0] ? byte_1536 : _GEN_5998; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6871 = mask_3[1] ? byte_1537 : _GEN_5999; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6872 = mask_3[2] ? byte_1538 : _GEN_6000; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6873 = mask_3[3] ? byte_1539 : _GEN_6001; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6874 = _GEN_9098 == 8'h5a ? _GEN_6870 : _GEN_5998; // @[executor.scala 473:84]
  wire [7:0] _GEN_6875 = _GEN_9098 == 8'h5a ? _GEN_6871 : _GEN_5999; // @[executor.scala 473:84]
  wire [7:0] _GEN_6876 = _GEN_9098 == 8'h5a ? _GEN_6872 : _GEN_6000; // @[executor.scala 473:84]
  wire [7:0] _GEN_6877 = _GEN_9098 == 8'h5a ? _GEN_6873 : _GEN_6001; // @[executor.scala 473:84]
  wire [7:0] _GEN_6878 = mask_3[0] ? byte_1536 : _GEN_6002; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6879 = mask_3[1] ? byte_1537 : _GEN_6003; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6880 = mask_3[2] ? byte_1538 : _GEN_6004; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6881 = mask_3[3] ? byte_1539 : _GEN_6005; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6882 = _GEN_9098 == 8'h5b ? _GEN_6878 : _GEN_6002; // @[executor.scala 473:84]
  wire [7:0] _GEN_6883 = _GEN_9098 == 8'h5b ? _GEN_6879 : _GEN_6003; // @[executor.scala 473:84]
  wire [7:0] _GEN_6884 = _GEN_9098 == 8'h5b ? _GEN_6880 : _GEN_6004; // @[executor.scala 473:84]
  wire [7:0] _GEN_6885 = _GEN_9098 == 8'h5b ? _GEN_6881 : _GEN_6005; // @[executor.scala 473:84]
  wire [7:0] _GEN_6886 = mask_3[0] ? byte_1536 : _GEN_6006; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6887 = mask_3[1] ? byte_1537 : _GEN_6007; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6888 = mask_3[2] ? byte_1538 : _GEN_6008; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6889 = mask_3[3] ? byte_1539 : _GEN_6009; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6890 = _GEN_9098 == 8'h5c ? _GEN_6886 : _GEN_6006; // @[executor.scala 473:84]
  wire [7:0] _GEN_6891 = _GEN_9098 == 8'h5c ? _GEN_6887 : _GEN_6007; // @[executor.scala 473:84]
  wire [7:0] _GEN_6892 = _GEN_9098 == 8'h5c ? _GEN_6888 : _GEN_6008; // @[executor.scala 473:84]
  wire [7:0] _GEN_6893 = _GEN_9098 == 8'h5c ? _GEN_6889 : _GEN_6009; // @[executor.scala 473:84]
  wire [7:0] _GEN_6894 = mask_3[0] ? byte_1536 : _GEN_6010; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6895 = mask_3[1] ? byte_1537 : _GEN_6011; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6896 = mask_3[2] ? byte_1538 : _GEN_6012; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6897 = mask_3[3] ? byte_1539 : _GEN_6013; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6898 = _GEN_9098 == 8'h5d ? _GEN_6894 : _GEN_6010; // @[executor.scala 473:84]
  wire [7:0] _GEN_6899 = _GEN_9098 == 8'h5d ? _GEN_6895 : _GEN_6011; // @[executor.scala 473:84]
  wire [7:0] _GEN_6900 = _GEN_9098 == 8'h5d ? _GEN_6896 : _GEN_6012; // @[executor.scala 473:84]
  wire [7:0] _GEN_6901 = _GEN_9098 == 8'h5d ? _GEN_6897 : _GEN_6013; // @[executor.scala 473:84]
  wire [7:0] _GEN_6902 = mask_3[0] ? byte_1536 : _GEN_6014; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6903 = mask_3[1] ? byte_1537 : _GEN_6015; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6904 = mask_3[2] ? byte_1538 : _GEN_6016; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6905 = mask_3[3] ? byte_1539 : _GEN_6017; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6906 = _GEN_9098 == 8'h5e ? _GEN_6902 : _GEN_6014; // @[executor.scala 473:84]
  wire [7:0] _GEN_6907 = _GEN_9098 == 8'h5e ? _GEN_6903 : _GEN_6015; // @[executor.scala 473:84]
  wire [7:0] _GEN_6908 = _GEN_9098 == 8'h5e ? _GEN_6904 : _GEN_6016; // @[executor.scala 473:84]
  wire [7:0] _GEN_6909 = _GEN_9098 == 8'h5e ? _GEN_6905 : _GEN_6017; // @[executor.scala 473:84]
  wire [7:0] _GEN_6910 = mask_3[0] ? byte_1536 : _GEN_6018; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6911 = mask_3[1] ? byte_1537 : _GEN_6019; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6912 = mask_3[2] ? byte_1538 : _GEN_6020; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6913 = mask_3[3] ? byte_1539 : _GEN_6021; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6914 = _GEN_9098 == 8'h5f ? _GEN_6910 : _GEN_6018; // @[executor.scala 473:84]
  wire [7:0] _GEN_6915 = _GEN_9098 == 8'h5f ? _GEN_6911 : _GEN_6019; // @[executor.scala 473:84]
  wire [7:0] _GEN_6916 = _GEN_9098 == 8'h5f ? _GEN_6912 : _GEN_6020; // @[executor.scala 473:84]
  wire [7:0] _GEN_6917 = _GEN_9098 == 8'h5f ? _GEN_6913 : _GEN_6021; // @[executor.scala 473:84]
  wire [7:0] _GEN_6918 = mask_3[0] ? byte_1536 : _GEN_6022; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6919 = mask_3[1] ? byte_1537 : _GEN_6023; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6920 = mask_3[2] ? byte_1538 : _GEN_6024; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6921 = mask_3[3] ? byte_1539 : _GEN_6025; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6922 = _GEN_9098 == 8'h60 ? _GEN_6918 : _GEN_6022; // @[executor.scala 473:84]
  wire [7:0] _GEN_6923 = _GEN_9098 == 8'h60 ? _GEN_6919 : _GEN_6023; // @[executor.scala 473:84]
  wire [7:0] _GEN_6924 = _GEN_9098 == 8'h60 ? _GEN_6920 : _GEN_6024; // @[executor.scala 473:84]
  wire [7:0] _GEN_6925 = _GEN_9098 == 8'h60 ? _GEN_6921 : _GEN_6025; // @[executor.scala 473:84]
  wire [7:0] _GEN_6926 = mask_3[0] ? byte_1536 : _GEN_6026; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6927 = mask_3[1] ? byte_1537 : _GEN_6027; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6928 = mask_3[2] ? byte_1538 : _GEN_6028; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6929 = mask_3[3] ? byte_1539 : _GEN_6029; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6930 = _GEN_9098 == 8'h61 ? _GEN_6926 : _GEN_6026; // @[executor.scala 473:84]
  wire [7:0] _GEN_6931 = _GEN_9098 == 8'h61 ? _GEN_6927 : _GEN_6027; // @[executor.scala 473:84]
  wire [7:0] _GEN_6932 = _GEN_9098 == 8'h61 ? _GEN_6928 : _GEN_6028; // @[executor.scala 473:84]
  wire [7:0] _GEN_6933 = _GEN_9098 == 8'h61 ? _GEN_6929 : _GEN_6029; // @[executor.scala 473:84]
  wire [7:0] _GEN_6934 = mask_3[0] ? byte_1536 : _GEN_6030; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6935 = mask_3[1] ? byte_1537 : _GEN_6031; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6936 = mask_3[2] ? byte_1538 : _GEN_6032; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6937 = mask_3[3] ? byte_1539 : _GEN_6033; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6938 = _GEN_9098 == 8'h62 ? _GEN_6934 : _GEN_6030; // @[executor.scala 473:84]
  wire [7:0] _GEN_6939 = _GEN_9098 == 8'h62 ? _GEN_6935 : _GEN_6031; // @[executor.scala 473:84]
  wire [7:0] _GEN_6940 = _GEN_9098 == 8'h62 ? _GEN_6936 : _GEN_6032; // @[executor.scala 473:84]
  wire [7:0] _GEN_6941 = _GEN_9098 == 8'h62 ? _GEN_6937 : _GEN_6033; // @[executor.scala 473:84]
  wire [7:0] _GEN_6942 = mask_3[0] ? byte_1536 : _GEN_6034; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6943 = mask_3[1] ? byte_1537 : _GEN_6035; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6944 = mask_3[2] ? byte_1538 : _GEN_6036; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6945 = mask_3[3] ? byte_1539 : _GEN_6037; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6946 = _GEN_9098 == 8'h63 ? _GEN_6942 : _GEN_6034; // @[executor.scala 473:84]
  wire [7:0] _GEN_6947 = _GEN_9098 == 8'h63 ? _GEN_6943 : _GEN_6035; // @[executor.scala 473:84]
  wire [7:0] _GEN_6948 = _GEN_9098 == 8'h63 ? _GEN_6944 : _GEN_6036; // @[executor.scala 473:84]
  wire [7:0] _GEN_6949 = _GEN_9098 == 8'h63 ? _GEN_6945 : _GEN_6037; // @[executor.scala 473:84]
  wire [7:0] _GEN_6950 = mask_3[0] ? byte_1536 : _GEN_6038; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6951 = mask_3[1] ? byte_1537 : _GEN_6039; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6952 = mask_3[2] ? byte_1538 : _GEN_6040; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6953 = mask_3[3] ? byte_1539 : _GEN_6041; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6954 = _GEN_9098 == 8'h64 ? _GEN_6950 : _GEN_6038; // @[executor.scala 473:84]
  wire [7:0] _GEN_6955 = _GEN_9098 == 8'h64 ? _GEN_6951 : _GEN_6039; // @[executor.scala 473:84]
  wire [7:0] _GEN_6956 = _GEN_9098 == 8'h64 ? _GEN_6952 : _GEN_6040; // @[executor.scala 473:84]
  wire [7:0] _GEN_6957 = _GEN_9098 == 8'h64 ? _GEN_6953 : _GEN_6041; // @[executor.scala 473:84]
  wire [7:0] _GEN_6958 = mask_3[0] ? byte_1536 : _GEN_6042; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6959 = mask_3[1] ? byte_1537 : _GEN_6043; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6960 = mask_3[2] ? byte_1538 : _GEN_6044; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6961 = mask_3[3] ? byte_1539 : _GEN_6045; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6962 = _GEN_9098 == 8'h65 ? _GEN_6958 : _GEN_6042; // @[executor.scala 473:84]
  wire [7:0] _GEN_6963 = _GEN_9098 == 8'h65 ? _GEN_6959 : _GEN_6043; // @[executor.scala 473:84]
  wire [7:0] _GEN_6964 = _GEN_9098 == 8'h65 ? _GEN_6960 : _GEN_6044; // @[executor.scala 473:84]
  wire [7:0] _GEN_6965 = _GEN_9098 == 8'h65 ? _GEN_6961 : _GEN_6045; // @[executor.scala 473:84]
  wire [7:0] _GEN_6966 = mask_3[0] ? byte_1536 : _GEN_6046; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6967 = mask_3[1] ? byte_1537 : _GEN_6047; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6968 = mask_3[2] ? byte_1538 : _GEN_6048; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6969 = mask_3[3] ? byte_1539 : _GEN_6049; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6970 = _GEN_9098 == 8'h66 ? _GEN_6966 : _GEN_6046; // @[executor.scala 473:84]
  wire [7:0] _GEN_6971 = _GEN_9098 == 8'h66 ? _GEN_6967 : _GEN_6047; // @[executor.scala 473:84]
  wire [7:0] _GEN_6972 = _GEN_9098 == 8'h66 ? _GEN_6968 : _GEN_6048; // @[executor.scala 473:84]
  wire [7:0] _GEN_6973 = _GEN_9098 == 8'h66 ? _GEN_6969 : _GEN_6049; // @[executor.scala 473:84]
  wire [7:0] _GEN_6974 = mask_3[0] ? byte_1536 : _GEN_6050; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6975 = mask_3[1] ? byte_1537 : _GEN_6051; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6976 = mask_3[2] ? byte_1538 : _GEN_6052; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6977 = mask_3[3] ? byte_1539 : _GEN_6053; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6978 = _GEN_9098 == 8'h67 ? _GEN_6974 : _GEN_6050; // @[executor.scala 473:84]
  wire [7:0] _GEN_6979 = _GEN_9098 == 8'h67 ? _GEN_6975 : _GEN_6051; // @[executor.scala 473:84]
  wire [7:0] _GEN_6980 = _GEN_9098 == 8'h67 ? _GEN_6976 : _GEN_6052; // @[executor.scala 473:84]
  wire [7:0] _GEN_6981 = _GEN_9098 == 8'h67 ? _GEN_6977 : _GEN_6053; // @[executor.scala 473:84]
  wire [7:0] _GEN_6982 = mask_3[0] ? byte_1536 : _GEN_6054; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6983 = mask_3[1] ? byte_1537 : _GEN_6055; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6984 = mask_3[2] ? byte_1538 : _GEN_6056; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6985 = mask_3[3] ? byte_1539 : _GEN_6057; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6986 = _GEN_9098 == 8'h68 ? _GEN_6982 : _GEN_6054; // @[executor.scala 473:84]
  wire [7:0] _GEN_6987 = _GEN_9098 == 8'h68 ? _GEN_6983 : _GEN_6055; // @[executor.scala 473:84]
  wire [7:0] _GEN_6988 = _GEN_9098 == 8'h68 ? _GEN_6984 : _GEN_6056; // @[executor.scala 473:84]
  wire [7:0] _GEN_6989 = _GEN_9098 == 8'h68 ? _GEN_6985 : _GEN_6057; // @[executor.scala 473:84]
  wire [7:0] _GEN_6990 = mask_3[0] ? byte_1536 : _GEN_6058; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6991 = mask_3[1] ? byte_1537 : _GEN_6059; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6992 = mask_3[2] ? byte_1538 : _GEN_6060; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6993 = mask_3[3] ? byte_1539 : _GEN_6061; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6994 = _GEN_9098 == 8'h69 ? _GEN_6990 : _GEN_6058; // @[executor.scala 473:84]
  wire [7:0] _GEN_6995 = _GEN_9098 == 8'h69 ? _GEN_6991 : _GEN_6059; // @[executor.scala 473:84]
  wire [7:0] _GEN_6996 = _GEN_9098 == 8'h69 ? _GEN_6992 : _GEN_6060; // @[executor.scala 473:84]
  wire [7:0] _GEN_6997 = _GEN_9098 == 8'h69 ? _GEN_6993 : _GEN_6061; // @[executor.scala 473:84]
  wire [7:0] _GEN_6998 = mask_3[0] ? byte_1536 : _GEN_6062; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_6999 = mask_3[1] ? byte_1537 : _GEN_6063; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7000 = mask_3[2] ? byte_1538 : _GEN_6064; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7001 = mask_3[3] ? byte_1539 : _GEN_6065; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7002 = _GEN_9098 == 8'h6a ? _GEN_6998 : _GEN_6062; // @[executor.scala 473:84]
  wire [7:0] _GEN_7003 = _GEN_9098 == 8'h6a ? _GEN_6999 : _GEN_6063; // @[executor.scala 473:84]
  wire [7:0] _GEN_7004 = _GEN_9098 == 8'h6a ? _GEN_7000 : _GEN_6064; // @[executor.scala 473:84]
  wire [7:0] _GEN_7005 = _GEN_9098 == 8'h6a ? _GEN_7001 : _GEN_6065; // @[executor.scala 473:84]
  wire [7:0] _GEN_7006 = mask_3[0] ? byte_1536 : _GEN_6066; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7007 = mask_3[1] ? byte_1537 : _GEN_6067; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7008 = mask_3[2] ? byte_1538 : _GEN_6068; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7009 = mask_3[3] ? byte_1539 : _GEN_6069; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7010 = _GEN_9098 == 8'h6b ? _GEN_7006 : _GEN_6066; // @[executor.scala 473:84]
  wire [7:0] _GEN_7011 = _GEN_9098 == 8'h6b ? _GEN_7007 : _GEN_6067; // @[executor.scala 473:84]
  wire [7:0] _GEN_7012 = _GEN_9098 == 8'h6b ? _GEN_7008 : _GEN_6068; // @[executor.scala 473:84]
  wire [7:0] _GEN_7013 = _GEN_9098 == 8'h6b ? _GEN_7009 : _GEN_6069; // @[executor.scala 473:84]
  wire [7:0] _GEN_7014 = mask_3[0] ? byte_1536 : _GEN_6070; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7015 = mask_3[1] ? byte_1537 : _GEN_6071; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7016 = mask_3[2] ? byte_1538 : _GEN_6072; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7017 = mask_3[3] ? byte_1539 : _GEN_6073; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7018 = _GEN_9098 == 8'h6c ? _GEN_7014 : _GEN_6070; // @[executor.scala 473:84]
  wire [7:0] _GEN_7019 = _GEN_9098 == 8'h6c ? _GEN_7015 : _GEN_6071; // @[executor.scala 473:84]
  wire [7:0] _GEN_7020 = _GEN_9098 == 8'h6c ? _GEN_7016 : _GEN_6072; // @[executor.scala 473:84]
  wire [7:0] _GEN_7021 = _GEN_9098 == 8'h6c ? _GEN_7017 : _GEN_6073; // @[executor.scala 473:84]
  wire [7:0] _GEN_7022 = mask_3[0] ? byte_1536 : _GEN_6074; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7023 = mask_3[1] ? byte_1537 : _GEN_6075; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7024 = mask_3[2] ? byte_1538 : _GEN_6076; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7025 = mask_3[3] ? byte_1539 : _GEN_6077; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7026 = _GEN_9098 == 8'h6d ? _GEN_7022 : _GEN_6074; // @[executor.scala 473:84]
  wire [7:0] _GEN_7027 = _GEN_9098 == 8'h6d ? _GEN_7023 : _GEN_6075; // @[executor.scala 473:84]
  wire [7:0] _GEN_7028 = _GEN_9098 == 8'h6d ? _GEN_7024 : _GEN_6076; // @[executor.scala 473:84]
  wire [7:0] _GEN_7029 = _GEN_9098 == 8'h6d ? _GEN_7025 : _GEN_6077; // @[executor.scala 473:84]
  wire [7:0] _GEN_7030 = mask_3[0] ? byte_1536 : _GEN_6078; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7031 = mask_3[1] ? byte_1537 : _GEN_6079; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7032 = mask_3[2] ? byte_1538 : _GEN_6080; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7033 = mask_3[3] ? byte_1539 : _GEN_6081; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7034 = _GEN_9098 == 8'h6e ? _GEN_7030 : _GEN_6078; // @[executor.scala 473:84]
  wire [7:0] _GEN_7035 = _GEN_9098 == 8'h6e ? _GEN_7031 : _GEN_6079; // @[executor.scala 473:84]
  wire [7:0] _GEN_7036 = _GEN_9098 == 8'h6e ? _GEN_7032 : _GEN_6080; // @[executor.scala 473:84]
  wire [7:0] _GEN_7037 = _GEN_9098 == 8'h6e ? _GEN_7033 : _GEN_6081; // @[executor.scala 473:84]
  wire [7:0] _GEN_7038 = mask_3[0] ? byte_1536 : _GEN_6082; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7039 = mask_3[1] ? byte_1537 : _GEN_6083; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7040 = mask_3[2] ? byte_1538 : _GEN_6084; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7041 = mask_3[3] ? byte_1539 : _GEN_6085; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7042 = _GEN_9098 == 8'h6f ? _GEN_7038 : _GEN_6082; // @[executor.scala 473:84]
  wire [7:0] _GEN_7043 = _GEN_9098 == 8'h6f ? _GEN_7039 : _GEN_6083; // @[executor.scala 473:84]
  wire [7:0] _GEN_7044 = _GEN_9098 == 8'h6f ? _GEN_7040 : _GEN_6084; // @[executor.scala 473:84]
  wire [7:0] _GEN_7045 = _GEN_9098 == 8'h6f ? _GEN_7041 : _GEN_6085; // @[executor.scala 473:84]
  wire [7:0] _GEN_7046 = mask_3[0] ? byte_1536 : _GEN_6086; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7047 = mask_3[1] ? byte_1537 : _GEN_6087; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7048 = mask_3[2] ? byte_1538 : _GEN_6088; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7049 = mask_3[3] ? byte_1539 : _GEN_6089; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7050 = _GEN_9098 == 8'h70 ? _GEN_7046 : _GEN_6086; // @[executor.scala 473:84]
  wire [7:0] _GEN_7051 = _GEN_9098 == 8'h70 ? _GEN_7047 : _GEN_6087; // @[executor.scala 473:84]
  wire [7:0] _GEN_7052 = _GEN_9098 == 8'h70 ? _GEN_7048 : _GEN_6088; // @[executor.scala 473:84]
  wire [7:0] _GEN_7053 = _GEN_9098 == 8'h70 ? _GEN_7049 : _GEN_6089; // @[executor.scala 473:84]
  wire [7:0] _GEN_7054 = mask_3[0] ? byte_1536 : _GEN_6090; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7055 = mask_3[1] ? byte_1537 : _GEN_6091; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7056 = mask_3[2] ? byte_1538 : _GEN_6092; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7057 = mask_3[3] ? byte_1539 : _GEN_6093; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7058 = _GEN_9098 == 8'h71 ? _GEN_7054 : _GEN_6090; // @[executor.scala 473:84]
  wire [7:0] _GEN_7059 = _GEN_9098 == 8'h71 ? _GEN_7055 : _GEN_6091; // @[executor.scala 473:84]
  wire [7:0] _GEN_7060 = _GEN_9098 == 8'h71 ? _GEN_7056 : _GEN_6092; // @[executor.scala 473:84]
  wire [7:0] _GEN_7061 = _GEN_9098 == 8'h71 ? _GEN_7057 : _GEN_6093; // @[executor.scala 473:84]
  wire [7:0] _GEN_7062 = mask_3[0] ? byte_1536 : _GEN_6094; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7063 = mask_3[1] ? byte_1537 : _GEN_6095; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7064 = mask_3[2] ? byte_1538 : _GEN_6096; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7065 = mask_3[3] ? byte_1539 : _GEN_6097; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7066 = _GEN_9098 == 8'h72 ? _GEN_7062 : _GEN_6094; // @[executor.scala 473:84]
  wire [7:0] _GEN_7067 = _GEN_9098 == 8'h72 ? _GEN_7063 : _GEN_6095; // @[executor.scala 473:84]
  wire [7:0] _GEN_7068 = _GEN_9098 == 8'h72 ? _GEN_7064 : _GEN_6096; // @[executor.scala 473:84]
  wire [7:0] _GEN_7069 = _GEN_9098 == 8'h72 ? _GEN_7065 : _GEN_6097; // @[executor.scala 473:84]
  wire [7:0] _GEN_7070 = mask_3[0] ? byte_1536 : _GEN_6098; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7071 = mask_3[1] ? byte_1537 : _GEN_6099; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7072 = mask_3[2] ? byte_1538 : _GEN_6100; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7073 = mask_3[3] ? byte_1539 : _GEN_6101; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7074 = _GEN_9098 == 8'h73 ? _GEN_7070 : _GEN_6098; // @[executor.scala 473:84]
  wire [7:0] _GEN_7075 = _GEN_9098 == 8'h73 ? _GEN_7071 : _GEN_6099; // @[executor.scala 473:84]
  wire [7:0] _GEN_7076 = _GEN_9098 == 8'h73 ? _GEN_7072 : _GEN_6100; // @[executor.scala 473:84]
  wire [7:0] _GEN_7077 = _GEN_9098 == 8'h73 ? _GEN_7073 : _GEN_6101; // @[executor.scala 473:84]
  wire [7:0] _GEN_7078 = mask_3[0] ? byte_1536 : _GEN_6102; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7079 = mask_3[1] ? byte_1537 : _GEN_6103; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7080 = mask_3[2] ? byte_1538 : _GEN_6104; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7081 = mask_3[3] ? byte_1539 : _GEN_6105; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7082 = _GEN_9098 == 8'h74 ? _GEN_7078 : _GEN_6102; // @[executor.scala 473:84]
  wire [7:0] _GEN_7083 = _GEN_9098 == 8'h74 ? _GEN_7079 : _GEN_6103; // @[executor.scala 473:84]
  wire [7:0] _GEN_7084 = _GEN_9098 == 8'h74 ? _GEN_7080 : _GEN_6104; // @[executor.scala 473:84]
  wire [7:0] _GEN_7085 = _GEN_9098 == 8'h74 ? _GEN_7081 : _GEN_6105; // @[executor.scala 473:84]
  wire [7:0] _GEN_7086 = mask_3[0] ? byte_1536 : _GEN_6106; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7087 = mask_3[1] ? byte_1537 : _GEN_6107; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7088 = mask_3[2] ? byte_1538 : _GEN_6108; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7089 = mask_3[3] ? byte_1539 : _GEN_6109; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7090 = _GEN_9098 == 8'h75 ? _GEN_7086 : _GEN_6106; // @[executor.scala 473:84]
  wire [7:0] _GEN_7091 = _GEN_9098 == 8'h75 ? _GEN_7087 : _GEN_6107; // @[executor.scala 473:84]
  wire [7:0] _GEN_7092 = _GEN_9098 == 8'h75 ? _GEN_7088 : _GEN_6108; // @[executor.scala 473:84]
  wire [7:0] _GEN_7093 = _GEN_9098 == 8'h75 ? _GEN_7089 : _GEN_6109; // @[executor.scala 473:84]
  wire [7:0] _GEN_7094 = mask_3[0] ? byte_1536 : _GEN_6110; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7095 = mask_3[1] ? byte_1537 : _GEN_6111; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7096 = mask_3[2] ? byte_1538 : _GEN_6112; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7097 = mask_3[3] ? byte_1539 : _GEN_6113; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7098 = _GEN_9098 == 8'h76 ? _GEN_7094 : _GEN_6110; // @[executor.scala 473:84]
  wire [7:0] _GEN_7099 = _GEN_9098 == 8'h76 ? _GEN_7095 : _GEN_6111; // @[executor.scala 473:84]
  wire [7:0] _GEN_7100 = _GEN_9098 == 8'h76 ? _GEN_7096 : _GEN_6112; // @[executor.scala 473:84]
  wire [7:0] _GEN_7101 = _GEN_9098 == 8'h76 ? _GEN_7097 : _GEN_6113; // @[executor.scala 473:84]
  wire [7:0] _GEN_7102 = mask_3[0] ? byte_1536 : _GEN_6114; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7103 = mask_3[1] ? byte_1537 : _GEN_6115; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7104 = mask_3[2] ? byte_1538 : _GEN_6116; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7105 = mask_3[3] ? byte_1539 : _GEN_6117; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7106 = _GEN_9098 == 8'h77 ? _GEN_7102 : _GEN_6114; // @[executor.scala 473:84]
  wire [7:0] _GEN_7107 = _GEN_9098 == 8'h77 ? _GEN_7103 : _GEN_6115; // @[executor.scala 473:84]
  wire [7:0] _GEN_7108 = _GEN_9098 == 8'h77 ? _GEN_7104 : _GEN_6116; // @[executor.scala 473:84]
  wire [7:0] _GEN_7109 = _GEN_9098 == 8'h77 ? _GEN_7105 : _GEN_6117; // @[executor.scala 473:84]
  wire [7:0] _GEN_7110 = mask_3[0] ? byte_1536 : _GEN_6118; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7111 = mask_3[1] ? byte_1537 : _GEN_6119; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7112 = mask_3[2] ? byte_1538 : _GEN_6120; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7113 = mask_3[3] ? byte_1539 : _GEN_6121; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7114 = _GEN_9098 == 8'h78 ? _GEN_7110 : _GEN_6118; // @[executor.scala 473:84]
  wire [7:0] _GEN_7115 = _GEN_9098 == 8'h78 ? _GEN_7111 : _GEN_6119; // @[executor.scala 473:84]
  wire [7:0] _GEN_7116 = _GEN_9098 == 8'h78 ? _GEN_7112 : _GEN_6120; // @[executor.scala 473:84]
  wire [7:0] _GEN_7117 = _GEN_9098 == 8'h78 ? _GEN_7113 : _GEN_6121; // @[executor.scala 473:84]
  wire [7:0] _GEN_7118 = mask_3[0] ? byte_1536 : _GEN_6122; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7119 = mask_3[1] ? byte_1537 : _GEN_6123; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7120 = mask_3[2] ? byte_1538 : _GEN_6124; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7121 = mask_3[3] ? byte_1539 : _GEN_6125; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7122 = _GEN_9098 == 8'h79 ? _GEN_7118 : _GEN_6122; // @[executor.scala 473:84]
  wire [7:0] _GEN_7123 = _GEN_9098 == 8'h79 ? _GEN_7119 : _GEN_6123; // @[executor.scala 473:84]
  wire [7:0] _GEN_7124 = _GEN_9098 == 8'h79 ? _GEN_7120 : _GEN_6124; // @[executor.scala 473:84]
  wire [7:0] _GEN_7125 = _GEN_9098 == 8'h79 ? _GEN_7121 : _GEN_6125; // @[executor.scala 473:84]
  wire [7:0] _GEN_7126 = mask_3[0] ? byte_1536 : _GEN_6126; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7127 = mask_3[1] ? byte_1537 : _GEN_6127; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7128 = mask_3[2] ? byte_1538 : _GEN_6128; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7129 = mask_3[3] ? byte_1539 : _GEN_6129; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7130 = _GEN_9098 == 8'h7a ? _GEN_7126 : _GEN_6126; // @[executor.scala 473:84]
  wire [7:0] _GEN_7131 = _GEN_9098 == 8'h7a ? _GEN_7127 : _GEN_6127; // @[executor.scala 473:84]
  wire [7:0] _GEN_7132 = _GEN_9098 == 8'h7a ? _GEN_7128 : _GEN_6128; // @[executor.scala 473:84]
  wire [7:0] _GEN_7133 = _GEN_9098 == 8'h7a ? _GEN_7129 : _GEN_6129; // @[executor.scala 473:84]
  wire [7:0] _GEN_7134 = mask_3[0] ? byte_1536 : _GEN_6130; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7135 = mask_3[1] ? byte_1537 : _GEN_6131; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7136 = mask_3[2] ? byte_1538 : _GEN_6132; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7137 = mask_3[3] ? byte_1539 : _GEN_6133; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7138 = _GEN_9098 == 8'h7b ? _GEN_7134 : _GEN_6130; // @[executor.scala 473:84]
  wire [7:0] _GEN_7139 = _GEN_9098 == 8'h7b ? _GEN_7135 : _GEN_6131; // @[executor.scala 473:84]
  wire [7:0] _GEN_7140 = _GEN_9098 == 8'h7b ? _GEN_7136 : _GEN_6132; // @[executor.scala 473:84]
  wire [7:0] _GEN_7141 = _GEN_9098 == 8'h7b ? _GEN_7137 : _GEN_6133; // @[executor.scala 473:84]
  wire [7:0] _GEN_7142 = mask_3[0] ? byte_1536 : _GEN_6134; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7143 = mask_3[1] ? byte_1537 : _GEN_6135; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7144 = mask_3[2] ? byte_1538 : _GEN_6136; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7145 = mask_3[3] ? byte_1539 : _GEN_6137; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7146 = _GEN_9098 == 8'h7c ? _GEN_7142 : _GEN_6134; // @[executor.scala 473:84]
  wire [7:0] _GEN_7147 = _GEN_9098 == 8'h7c ? _GEN_7143 : _GEN_6135; // @[executor.scala 473:84]
  wire [7:0] _GEN_7148 = _GEN_9098 == 8'h7c ? _GEN_7144 : _GEN_6136; // @[executor.scala 473:84]
  wire [7:0] _GEN_7149 = _GEN_9098 == 8'h7c ? _GEN_7145 : _GEN_6137; // @[executor.scala 473:84]
  wire [7:0] _GEN_7150 = mask_3[0] ? byte_1536 : _GEN_6138; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7151 = mask_3[1] ? byte_1537 : _GEN_6139; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7152 = mask_3[2] ? byte_1538 : _GEN_6140; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7153 = mask_3[3] ? byte_1539 : _GEN_6141; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7154 = _GEN_9098 == 8'h7d ? _GEN_7150 : _GEN_6138; // @[executor.scala 473:84]
  wire [7:0] _GEN_7155 = _GEN_9098 == 8'h7d ? _GEN_7151 : _GEN_6139; // @[executor.scala 473:84]
  wire [7:0] _GEN_7156 = _GEN_9098 == 8'h7d ? _GEN_7152 : _GEN_6140; // @[executor.scala 473:84]
  wire [7:0] _GEN_7157 = _GEN_9098 == 8'h7d ? _GEN_7153 : _GEN_6141; // @[executor.scala 473:84]
  wire [7:0] _GEN_7158 = mask_3[0] ? byte_1536 : _GEN_6142; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7159 = mask_3[1] ? byte_1537 : _GEN_6143; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7160 = mask_3[2] ? byte_1538 : _GEN_6144; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7161 = mask_3[3] ? byte_1539 : _GEN_6145; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7162 = _GEN_9098 == 8'h7e ? _GEN_7158 : _GEN_6142; // @[executor.scala 473:84]
  wire [7:0] _GEN_7163 = _GEN_9098 == 8'h7e ? _GEN_7159 : _GEN_6143; // @[executor.scala 473:84]
  wire [7:0] _GEN_7164 = _GEN_9098 == 8'h7e ? _GEN_7160 : _GEN_6144; // @[executor.scala 473:84]
  wire [7:0] _GEN_7165 = _GEN_9098 == 8'h7e ? _GEN_7161 : _GEN_6145; // @[executor.scala 473:84]
  wire [7:0] _GEN_7166 = mask_3[0] ? byte_1536 : _GEN_6146; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7167 = mask_3[1] ? byte_1537 : _GEN_6147; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7168 = mask_3[2] ? byte_1538 : _GEN_6148; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7169 = mask_3[3] ? byte_1539 : _GEN_6149; // @[executor.scala 476:55 executor.scala 477:71]
  wire [7:0] _GEN_7170 = _GEN_9098 == 8'h7f ? _GEN_7166 : _GEN_6146; // @[executor.scala 473:84]
  wire [7:0] _GEN_7171 = _GEN_9098 == 8'h7f ? _GEN_7167 : _GEN_6147; // @[executor.scala 473:84]
  wire [7:0] _GEN_7172 = _GEN_9098 == 8'h7f ? _GEN_7168 : _GEN_6148; // @[executor.scala 473:84]
  wire [7:0] _GEN_7173 = _GEN_9098 == 8'h7f ? _GEN_7169 : _GEN_6149; // @[executor.scala 473:84]
  wire [7:0] _GEN_7174 = opcode_3 != 4'h0 ? _GEN_6154 : _GEN_5638; // @[executor.scala 470:55]
  wire [7:0] _GEN_7175 = opcode_3 != 4'h0 ? _GEN_6155 : _GEN_5639; // @[executor.scala 470:55]
  wire [7:0] _GEN_7176 = opcode_3 != 4'h0 ? _GEN_6156 : _GEN_5640; // @[executor.scala 470:55]
  wire [7:0] _GEN_7177 = opcode_3 != 4'h0 ? _GEN_6157 : _GEN_5641; // @[executor.scala 470:55]
  wire [7:0] _GEN_7178 = opcode_3 != 4'h0 ? _GEN_6162 : _GEN_5642; // @[executor.scala 470:55]
  wire [7:0] _GEN_7179 = opcode_3 != 4'h0 ? _GEN_6163 : _GEN_5643; // @[executor.scala 470:55]
  wire [7:0] _GEN_7180 = opcode_3 != 4'h0 ? _GEN_6164 : _GEN_5644; // @[executor.scala 470:55]
  wire [7:0] _GEN_7181 = opcode_3 != 4'h0 ? _GEN_6165 : _GEN_5645; // @[executor.scala 470:55]
  wire [7:0] _GEN_7182 = opcode_3 != 4'h0 ? _GEN_6170 : _GEN_5646; // @[executor.scala 470:55]
  wire [7:0] _GEN_7183 = opcode_3 != 4'h0 ? _GEN_6171 : _GEN_5647; // @[executor.scala 470:55]
  wire [7:0] _GEN_7184 = opcode_3 != 4'h0 ? _GEN_6172 : _GEN_5648; // @[executor.scala 470:55]
  wire [7:0] _GEN_7185 = opcode_3 != 4'h0 ? _GEN_6173 : _GEN_5649; // @[executor.scala 470:55]
  wire [7:0] _GEN_7186 = opcode_3 != 4'h0 ? _GEN_6178 : _GEN_5650; // @[executor.scala 470:55]
  wire [7:0] _GEN_7187 = opcode_3 != 4'h0 ? _GEN_6179 : _GEN_5651; // @[executor.scala 470:55]
  wire [7:0] _GEN_7188 = opcode_3 != 4'h0 ? _GEN_6180 : _GEN_5652; // @[executor.scala 470:55]
  wire [7:0] _GEN_7189 = opcode_3 != 4'h0 ? _GEN_6181 : _GEN_5653; // @[executor.scala 470:55]
  wire [7:0] _GEN_7190 = opcode_3 != 4'h0 ? _GEN_6186 : _GEN_5654; // @[executor.scala 470:55]
  wire [7:0] _GEN_7191 = opcode_3 != 4'h0 ? _GEN_6187 : _GEN_5655; // @[executor.scala 470:55]
  wire [7:0] _GEN_7192 = opcode_3 != 4'h0 ? _GEN_6188 : _GEN_5656; // @[executor.scala 470:55]
  wire [7:0] _GEN_7193 = opcode_3 != 4'h0 ? _GEN_6189 : _GEN_5657; // @[executor.scala 470:55]
  wire [7:0] _GEN_7194 = opcode_3 != 4'h0 ? _GEN_6194 : _GEN_5658; // @[executor.scala 470:55]
  wire [7:0] _GEN_7195 = opcode_3 != 4'h0 ? _GEN_6195 : _GEN_5659; // @[executor.scala 470:55]
  wire [7:0] _GEN_7196 = opcode_3 != 4'h0 ? _GEN_6196 : _GEN_5660; // @[executor.scala 470:55]
  wire [7:0] _GEN_7197 = opcode_3 != 4'h0 ? _GEN_6197 : _GEN_5661; // @[executor.scala 470:55]
  wire [7:0] _GEN_7198 = opcode_3 != 4'h0 ? _GEN_6202 : _GEN_5662; // @[executor.scala 470:55]
  wire [7:0] _GEN_7199 = opcode_3 != 4'h0 ? _GEN_6203 : _GEN_5663; // @[executor.scala 470:55]
  wire [7:0] _GEN_7200 = opcode_3 != 4'h0 ? _GEN_6204 : _GEN_5664; // @[executor.scala 470:55]
  wire [7:0] _GEN_7201 = opcode_3 != 4'h0 ? _GEN_6205 : _GEN_5665; // @[executor.scala 470:55]
  wire [7:0] _GEN_7202 = opcode_3 != 4'h0 ? _GEN_6210 : _GEN_5666; // @[executor.scala 470:55]
  wire [7:0] _GEN_7203 = opcode_3 != 4'h0 ? _GEN_6211 : _GEN_5667; // @[executor.scala 470:55]
  wire [7:0] _GEN_7204 = opcode_3 != 4'h0 ? _GEN_6212 : _GEN_5668; // @[executor.scala 470:55]
  wire [7:0] _GEN_7205 = opcode_3 != 4'h0 ? _GEN_6213 : _GEN_5669; // @[executor.scala 470:55]
  wire [7:0] _GEN_7206 = opcode_3 != 4'h0 ? _GEN_6218 : _GEN_5670; // @[executor.scala 470:55]
  wire [7:0] _GEN_7207 = opcode_3 != 4'h0 ? _GEN_6219 : _GEN_5671; // @[executor.scala 470:55]
  wire [7:0] _GEN_7208 = opcode_3 != 4'h0 ? _GEN_6220 : _GEN_5672; // @[executor.scala 470:55]
  wire [7:0] _GEN_7209 = opcode_3 != 4'h0 ? _GEN_6221 : _GEN_5673; // @[executor.scala 470:55]
  wire [7:0] _GEN_7210 = opcode_3 != 4'h0 ? _GEN_6226 : _GEN_5674; // @[executor.scala 470:55]
  wire [7:0] _GEN_7211 = opcode_3 != 4'h0 ? _GEN_6227 : _GEN_5675; // @[executor.scala 470:55]
  wire [7:0] _GEN_7212 = opcode_3 != 4'h0 ? _GEN_6228 : _GEN_5676; // @[executor.scala 470:55]
  wire [7:0] _GEN_7213 = opcode_3 != 4'h0 ? _GEN_6229 : _GEN_5677; // @[executor.scala 470:55]
  wire [7:0] _GEN_7214 = opcode_3 != 4'h0 ? _GEN_6234 : _GEN_5678; // @[executor.scala 470:55]
  wire [7:0] _GEN_7215 = opcode_3 != 4'h0 ? _GEN_6235 : _GEN_5679; // @[executor.scala 470:55]
  wire [7:0] _GEN_7216 = opcode_3 != 4'h0 ? _GEN_6236 : _GEN_5680; // @[executor.scala 470:55]
  wire [7:0] _GEN_7217 = opcode_3 != 4'h0 ? _GEN_6237 : _GEN_5681; // @[executor.scala 470:55]
  wire [7:0] _GEN_7218 = opcode_3 != 4'h0 ? _GEN_6242 : _GEN_5682; // @[executor.scala 470:55]
  wire [7:0] _GEN_7219 = opcode_3 != 4'h0 ? _GEN_6243 : _GEN_5683; // @[executor.scala 470:55]
  wire [7:0] _GEN_7220 = opcode_3 != 4'h0 ? _GEN_6244 : _GEN_5684; // @[executor.scala 470:55]
  wire [7:0] _GEN_7221 = opcode_3 != 4'h0 ? _GEN_6245 : _GEN_5685; // @[executor.scala 470:55]
  wire [7:0] _GEN_7222 = opcode_3 != 4'h0 ? _GEN_6250 : _GEN_5686; // @[executor.scala 470:55]
  wire [7:0] _GEN_7223 = opcode_3 != 4'h0 ? _GEN_6251 : _GEN_5687; // @[executor.scala 470:55]
  wire [7:0] _GEN_7224 = opcode_3 != 4'h0 ? _GEN_6252 : _GEN_5688; // @[executor.scala 470:55]
  wire [7:0] _GEN_7225 = opcode_3 != 4'h0 ? _GEN_6253 : _GEN_5689; // @[executor.scala 470:55]
  wire [7:0] _GEN_7226 = opcode_3 != 4'h0 ? _GEN_6258 : _GEN_5690; // @[executor.scala 470:55]
  wire [7:0] _GEN_7227 = opcode_3 != 4'h0 ? _GEN_6259 : _GEN_5691; // @[executor.scala 470:55]
  wire [7:0] _GEN_7228 = opcode_3 != 4'h0 ? _GEN_6260 : _GEN_5692; // @[executor.scala 470:55]
  wire [7:0] _GEN_7229 = opcode_3 != 4'h0 ? _GEN_6261 : _GEN_5693; // @[executor.scala 470:55]
  wire [7:0] _GEN_7230 = opcode_3 != 4'h0 ? _GEN_6266 : _GEN_5694; // @[executor.scala 470:55]
  wire [7:0] _GEN_7231 = opcode_3 != 4'h0 ? _GEN_6267 : _GEN_5695; // @[executor.scala 470:55]
  wire [7:0] _GEN_7232 = opcode_3 != 4'h0 ? _GEN_6268 : _GEN_5696; // @[executor.scala 470:55]
  wire [7:0] _GEN_7233 = opcode_3 != 4'h0 ? _GEN_6269 : _GEN_5697; // @[executor.scala 470:55]
  wire [7:0] _GEN_7234 = opcode_3 != 4'h0 ? _GEN_6274 : _GEN_5698; // @[executor.scala 470:55]
  wire [7:0] _GEN_7235 = opcode_3 != 4'h0 ? _GEN_6275 : _GEN_5699; // @[executor.scala 470:55]
  wire [7:0] _GEN_7236 = opcode_3 != 4'h0 ? _GEN_6276 : _GEN_5700; // @[executor.scala 470:55]
  wire [7:0] _GEN_7237 = opcode_3 != 4'h0 ? _GEN_6277 : _GEN_5701; // @[executor.scala 470:55]
  wire [7:0] _GEN_7238 = opcode_3 != 4'h0 ? _GEN_6282 : _GEN_5702; // @[executor.scala 470:55]
  wire [7:0] _GEN_7239 = opcode_3 != 4'h0 ? _GEN_6283 : _GEN_5703; // @[executor.scala 470:55]
  wire [7:0] _GEN_7240 = opcode_3 != 4'h0 ? _GEN_6284 : _GEN_5704; // @[executor.scala 470:55]
  wire [7:0] _GEN_7241 = opcode_3 != 4'h0 ? _GEN_6285 : _GEN_5705; // @[executor.scala 470:55]
  wire [7:0] _GEN_7242 = opcode_3 != 4'h0 ? _GEN_6290 : _GEN_5706; // @[executor.scala 470:55]
  wire [7:0] _GEN_7243 = opcode_3 != 4'h0 ? _GEN_6291 : _GEN_5707; // @[executor.scala 470:55]
  wire [7:0] _GEN_7244 = opcode_3 != 4'h0 ? _GEN_6292 : _GEN_5708; // @[executor.scala 470:55]
  wire [7:0] _GEN_7245 = opcode_3 != 4'h0 ? _GEN_6293 : _GEN_5709; // @[executor.scala 470:55]
  wire [7:0] _GEN_7246 = opcode_3 != 4'h0 ? _GEN_6298 : _GEN_5710; // @[executor.scala 470:55]
  wire [7:0] _GEN_7247 = opcode_3 != 4'h0 ? _GEN_6299 : _GEN_5711; // @[executor.scala 470:55]
  wire [7:0] _GEN_7248 = opcode_3 != 4'h0 ? _GEN_6300 : _GEN_5712; // @[executor.scala 470:55]
  wire [7:0] _GEN_7249 = opcode_3 != 4'h0 ? _GEN_6301 : _GEN_5713; // @[executor.scala 470:55]
  wire [7:0] _GEN_7250 = opcode_3 != 4'h0 ? _GEN_6306 : _GEN_5714; // @[executor.scala 470:55]
  wire [7:0] _GEN_7251 = opcode_3 != 4'h0 ? _GEN_6307 : _GEN_5715; // @[executor.scala 470:55]
  wire [7:0] _GEN_7252 = opcode_3 != 4'h0 ? _GEN_6308 : _GEN_5716; // @[executor.scala 470:55]
  wire [7:0] _GEN_7253 = opcode_3 != 4'h0 ? _GEN_6309 : _GEN_5717; // @[executor.scala 470:55]
  wire [7:0] _GEN_7254 = opcode_3 != 4'h0 ? _GEN_6314 : _GEN_5718; // @[executor.scala 470:55]
  wire [7:0] _GEN_7255 = opcode_3 != 4'h0 ? _GEN_6315 : _GEN_5719; // @[executor.scala 470:55]
  wire [7:0] _GEN_7256 = opcode_3 != 4'h0 ? _GEN_6316 : _GEN_5720; // @[executor.scala 470:55]
  wire [7:0] _GEN_7257 = opcode_3 != 4'h0 ? _GEN_6317 : _GEN_5721; // @[executor.scala 470:55]
  wire [7:0] _GEN_7258 = opcode_3 != 4'h0 ? _GEN_6322 : _GEN_5722; // @[executor.scala 470:55]
  wire [7:0] _GEN_7259 = opcode_3 != 4'h0 ? _GEN_6323 : _GEN_5723; // @[executor.scala 470:55]
  wire [7:0] _GEN_7260 = opcode_3 != 4'h0 ? _GEN_6324 : _GEN_5724; // @[executor.scala 470:55]
  wire [7:0] _GEN_7261 = opcode_3 != 4'h0 ? _GEN_6325 : _GEN_5725; // @[executor.scala 470:55]
  wire [7:0] _GEN_7262 = opcode_3 != 4'h0 ? _GEN_6330 : _GEN_5726; // @[executor.scala 470:55]
  wire [7:0] _GEN_7263 = opcode_3 != 4'h0 ? _GEN_6331 : _GEN_5727; // @[executor.scala 470:55]
  wire [7:0] _GEN_7264 = opcode_3 != 4'h0 ? _GEN_6332 : _GEN_5728; // @[executor.scala 470:55]
  wire [7:0] _GEN_7265 = opcode_3 != 4'h0 ? _GEN_6333 : _GEN_5729; // @[executor.scala 470:55]
  wire [7:0] _GEN_7266 = opcode_3 != 4'h0 ? _GEN_6338 : _GEN_5730; // @[executor.scala 470:55]
  wire [7:0] _GEN_7267 = opcode_3 != 4'h0 ? _GEN_6339 : _GEN_5731; // @[executor.scala 470:55]
  wire [7:0] _GEN_7268 = opcode_3 != 4'h0 ? _GEN_6340 : _GEN_5732; // @[executor.scala 470:55]
  wire [7:0] _GEN_7269 = opcode_3 != 4'h0 ? _GEN_6341 : _GEN_5733; // @[executor.scala 470:55]
  wire [7:0] _GEN_7270 = opcode_3 != 4'h0 ? _GEN_6346 : _GEN_5734; // @[executor.scala 470:55]
  wire [7:0] _GEN_7271 = opcode_3 != 4'h0 ? _GEN_6347 : _GEN_5735; // @[executor.scala 470:55]
  wire [7:0] _GEN_7272 = opcode_3 != 4'h0 ? _GEN_6348 : _GEN_5736; // @[executor.scala 470:55]
  wire [7:0] _GEN_7273 = opcode_3 != 4'h0 ? _GEN_6349 : _GEN_5737; // @[executor.scala 470:55]
  wire [7:0] _GEN_7274 = opcode_3 != 4'h0 ? _GEN_6354 : _GEN_5738; // @[executor.scala 470:55]
  wire [7:0] _GEN_7275 = opcode_3 != 4'h0 ? _GEN_6355 : _GEN_5739; // @[executor.scala 470:55]
  wire [7:0] _GEN_7276 = opcode_3 != 4'h0 ? _GEN_6356 : _GEN_5740; // @[executor.scala 470:55]
  wire [7:0] _GEN_7277 = opcode_3 != 4'h0 ? _GEN_6357 : _GEN_5741; // @[executor.scala 470:55]
  wire [7:0] _GEN_7278 = opcode_3 != 4'h0 ? _GEN_6362 : _GEN_5742; // @[executor.scala 470:55]
  wire [7:0] _GEN_7279 = opcode_3 != 4'h0 ? _GEN_6363 : _GEN_5743; // @[executor.scala 470:55]
  wire [7:0] _GEN_7280 = opcode_3 != 4'h0 ? _GEN_6364 : _GEN_5744; // @[executor.scala 470:55]
  wire [7:0] _GEN_7281 = opcode_3 != 4'h0 ? _GEN_6365 : _GEN_5745; // @[executor.scala 470:55]
  wire [7:0] _GEN_7282 = opcode_3 != 4'h0 ? _GEN_6370 : _GEN_5746; // @[executor.scala 470:55]
  wire [7:0] _GEN_7283 = opcode_3 != 4'h0 ? _GEN_6371 : _GEN_5747; // @[executor.scala 470:55]
  wire [7:0] _GEN_7284 = opcode_3 != 4'h0 ? _GEN_6372 : _GEN_5748; // @[executor.scala 470:55]
  wire [7:0] _GEN_7285 = opcode_3 != 4'h0 ? _GEN_6373 : _GEN_5749; // @[executor.scala 470:55]
  wire [7:0] _GEN_7286 = opcode_3 != 4'h0 ? _GEN_6378 : _GEN_5750; // @[executor.scala 470:55]
  wire [7:0] _GEN_7287 = opcode_3 != 4'h0 ? _GEN_6379 : _GEN_5751; // @[executor.scala 470:55]
  wire [7:0] _GEN_7288 = opcode_3 != 4'h0 ? _GEN_6380 : _GEN_5752; // @[executor.scala 470:55]
  wire [7:0] _GEN_7289 = opcode_3 != 4'h0 ? _GEN_6381 : _GEN_5753; // @[executor.scala 470:55]
  wire [7:0] _GEN_7290 = opcode_3 != 4'h0 ? _GEN_6386 : _GEN_5754; // @[executor.scala 470:55]
  wire [7:0] _GEN_7291 = opcode_3 != 4'h0 ? _GEN_6387 : _GEN_5755; // @[executor.scala 470:55]
  wire [7:0] _GEN_7292 = opcode_3 != 4'h0 ? _GEN_6388 : _GEN_5756; // @[executor.scala 470:55]
  wire [7:0] _GEN_7293 = opcode_3 != 4'h0 ? _GEN_6389 : _GEN_5757; // @[executor.scala 470:55]
  wire [7:0] _GEN_7294 = opcode_3 != 4'h0 ? _GEN_6394 : _GEN_5758; // @[executor.scala 470:55]
  wire [7:0] _GEN_7295 = opcode_3 != 4'h0 ? _GEN_6395 : _GEN_5759; // @[executor.scala 470:55]
  wire [7:0] _GEN_7296 = opcode_3 != 4'h0 ? _GEN_6396 : _GEN_5760; // @[executor.scala 470:55]
  wire [7:0] _GEN_7297 = opcode_3 != 4'h0 ? _GEN_6397 : _GEN_5761; // @[executor.scala 470:55]
  wire [7:0] _GEN_7298 = opcode_3 != 4'h0 ? _GEN_6402 : _GEN_5762; // @[executor.scala 470:55]
  wire [7:0] _GEN_7299 = opcode_3 != 4'h0 ? _GEN_6403 : _GEN_5763; // @[executor.scala 470:55]
  wire [7:0] _GEN_7300 = opcode_3 != 4'h0 ? _GEN_6404 : _GEN_5764; // @[executor.scala 470:55]
  wire [7:0] _GEN_7301 = opcode_3 != 4'h0 ? _GEN_6405 : _GEN_5765; // @[executor.scala 470:55]
  wire [7:0] _GEN_7302 = opcode_3 != 4'h0 ? _GEN_6410 : _GEN_5766; // @[executor.scala 470:55]
  wire [7:0] _GEN_7303 = opcode_3 != 4'h0 ? _GEN_6411 : _GEN_5767; // @[executor.scala 470:55]
  wire [7:0] _GEN_7304 = opcode_3 != 4'h0 ? _GEN_6412 : _GEN_5768; // @[executor.scala 470:55]
  wire [7:0] _GEN_7305 = opcode_3 != 4'h0 ? _GEN_6413 : _GEN_5769; // @[executor.scala 470:55]
  wire [7:0] _GEN_7306 = opcode_3 != 4'h0 ? _GEN_6418 : _GEN_5770; // @[executor.scala 470:55]
  wire [7:0] _GEN_7307 = opcode_3 != 4'h0 ? _GEN_6419 : _GEN_5771; // @[executor.scala 470:55]
  wire [7:0] _GEN_7308 = opcode_3 != 4'h0 ? _GEN_6420 : _GEN_5772; // @[executor.scala 470:55]
  wire [7:0] _GEN_7309 = opcode_3 != 4'h0 ? _GEN_6421 : _GEN_5773; // @[executor.scala 470:55]
  wire [7:0] _GEN_7310 = opcode_3 != 4'h0 ? _GEN_6426 : _GEN_5774; // @[executor.scala 470:55]
  wire [7:0] _GEN_7311 = opcode_3 != 4'h0 ? _GEN_6427 : _GEN_5775; // @[executor.scala 470:55]
  wire [7:0] _GEN_7312 = opcode_3 != 4'h0 ? _GEN_6428 : _GEN_5776; // @[executor.scala 470:55]
  wire [7:0] _GEN_7313 = opcode_3 != 4'h0 ? _GEN_6429 : _GEN_5777; // @[executor.scala 470:55]
  wire [7:0] _GEN_7314 = opcode_3 != 4'h0 ? _GEN_6434 : _GEN_5778; // @[executor.scala 470:55]
  wire [7:0] _GEN_7315 = opcode_3 != 4'h0 ? _GEN_6435 : _GEN_5779; // @[executor.scala 470:55]
  wire [7:0] _GEN_7316 = opcode_3 != 4'h0 ? _GEN_6436 : _GEN_5780; // @[executor.scala 470:55]
  wire [7:0] _GEN_7317 = opcode_3 != 4'h0 ? _GEN_6437 : _GEN_5781; // @[executor.scala 470:55]
  wire [7:0] _GEN_7318 = opcode_3 != 4'h0 ? _GEN_6442 : _GEN_5782; // @[executor.scala 470:55]
  wire [7:0] _GEN_7319 = opcode_3 != 4'h0 ? _GEN_6443 : _GEN_5783; // @[executor.scala 470:55]
  wire [7:0] _GEN_7320 = opcode_3 != 4'h0 ? _GEN_6444 : _GEN_5784; // @[executor.scala 470:55]
  wire [7:0] _GEN_7321 = opcode_3 != 4'h0 ? _GEN_6445 : _GEN_5785; // @[executor.scala 470:55]
  wire [7:0] _GEN_7322 = opcode_3 != 4'h0 ? _GEN_6450 : _GEN_5786; // @[executor.scala 470:55]
  wire [7:0] _GEN_7323 = opcode_3 != 4'h0 ? _GEN_6451 : _GEN_5787; // @[executor.scala 470:55]
  wire [7:0] _GEN_7324 = opcode_3 != 4'h0 ? _GEN_6452 : _GEN_5788; // @[executor.scala 470:55]
  wire [7:0] _GEN_7325 = opcode_3 != 4'h0 ? _GEN_6453 : _GEN_5789; // @[executor.scala 470:55]
  wire [7:0] _GEN_7326 = opcode_3 != 4'h0 ? _GEN_6458 : _GEN_5790; // @[executor.scala 470:55]
  wire [7:0] _GEN_7327 = opcode_3 != 4'h0 ? _GEN_6459 : _GEN_5791; // @[executor.scala 470:55]
  wire [7:0] _GEN_7328 = opcode_3 != 4'h0 ? _GEN_6460 : _GEN_5792; // @[executor.scala 470:55]
  wire [7:0] _GEN_7329 = opcode_3 != 4'h0 ? _GEN_6461 : _GEN_5793; // @[executor.scala 470:55]
  wire [7:0] _GEN_7330 = opcode_3 != 4'h0 ? _GEN_6466 : _GEN_5794; // @[executor.scala 470:55]
  wire [7:0] _GEN_7331 = opcode_3 != 4'h0 ? _GEN_6467 : _GEN_5795; // @[executor.scala 470:55]
  wire [7:0] _GEN_7332 = opcode_3 != 4'h0 ? _GEN_6468 : _GEN_5796; // @[executor.scala 470:55]
  wire [7:0] _GEN_7333 = opcode_3 != 4'h0 ? _GEN_6469 : _GEN_5797; // @[executor.scala 470:55]
  wire [7:0] _GEN_7334 = opcode_3 != 4'h0 ? _GEN_6474 : _GEN_5798; // @[executor.scala 470:55]
  wire [7:0] _GEN_7335 = opcode_3 != 4'h0 ? _GEN_6475 : _GEN_5799; // @[executor.scala 470:55]
  wire [7:0] _GEN_7336 = opcode_3 != 4'h0 ? _GEN_6476 : _GEN_5800; // @[executor.scala 470:55]
  wire [7:0] _GEN_7337 = opcode_3 != 4'h0 ? _GEN_6477 : _GEN_5801; // @[executor.scala 470:55]
  wire [7:0] _GEN_7338 = opcode_3 != 4'h0 ? _GEN_6482 : _GEN_5802; // @[executor.scala 470:55]
  wire [7:0] _GEN_7339 = opcode_3 != 4'h0 ? _GEN_6483 : _GEN_5803; // @[executor.scala 470:55]
  wire [7:0] _GEN_7340 = opcode_3 != 4'h0 ? _GEN_6484 : _GEN_5804; // @[executor.scala 470:55]
  wire [7:0] _GEN_7341 = opcode_3 != 4'h0 ? _GEN_6485 : _GEN_5805; // @[executor.scala 470:55]
  wire [7:0] _GEN_7342 = opcode_3 != 4'h0 ? _GEN_6490 : _GEN_5806; // @[executor.scala 470:55]
  wire [7:0] _GEN_7343 = opcode_3 != 4'h0 ? _GEN_6491 : _GEN_5807; // @[executor.scala 470:55]
  wire [7:0] _GEN_7344 = opcode_3 != 4'h0 ? _GEN_6492 : _GEN_5808; // @[executor.scala 470:55]
  wire [7:0] _GEN_7345 = opcode_3 != 4'h0 ? _GEN_6493 : _GEN_5809; // @[executor.scala 470:55]
  wire [7:0] _GEN_7346 = opcode_3 != 4'h0 ? _GEN_6498 : _GEN_5810; // @[executor.scala 470:55]
  wire [7:0] _GEN_7347 = opcode_3 != 4'h0 ? _GEN_6499 : _GEN_5811; // @[executor.scala 470:55]
  wire [7:0] _GEN_7348 = opcode_3 != 4'h0 ? _GEN_6500 : _GEN_5812; // @[executor.scala 470:55]
  wire [7:0] _GEN_7349 = opcode_3 != 4'h0 ? _GEN_6501 : _GEN_5813; // @[executor.scala 470:55]
  wire [7:0] _GEN_7350 = opcode_3 != 4'h0 ? _GEN_6506 : _GEN_5814; // @[executor.scala 470:55]
  wire [7:0] _GEN_7351 = opcode_3 != 4'h0 ? _GEN_6507 : _GEN_5815; // @[executor.scala 470:55]
  wire [7:0] _GEN_7352 = opcode_3 != 4'h0 ? _GEN_6508 : _GEN_5816; // @[executor.scala 470:55]
  wire [7:0] _GEN_7353 = opcode_3 != 4'h0 ? _GEN_6509 : _GEN_5817; // @[executor.scala 470:55]
  wire [7:0] _GEN_7354 = opcode_3 != 4'h0 ? _GEN_6514 : _GEN_5818; // @[executor.scala 470:55]
  wire [7:0] _GEN_7355 = opcode_3 != 4'h0 ? _GEN_6515 : _GEN_5819; // @[executor.scala 470:55]
  wire [7:0] _GEN_7356 = opcode_3 != 4'h0 ? _GEN_6516 : _GEN_5820; // @[executor.scala 470:55]
  wire [7:0] _GEN_7357 = opcode_3 != 4'h0 ? _GEN_6517 : _GEN_5821; // @[executor.scala 470:55]
  wire [7:0] _GEN_7358 = opcode_3 != 4'h0 ? _GEN_6522 : _GEN_5822; // @[executor.scala 470:55]
  wire [7:0] _GEN_7359 = opcode_3 != 4'h0 ? _GEN_6523 : _GEN_5823; // @[executor.scala 470:55]
  wire [7:0] _GEN_7360 = opcode_3 != 4'h0 ? _GEN_6524 : _GEN_5824; // @[executor.scala 470:55]
  wire [7:0] _GEN_7361 = opcode_3 != 4'h0 ? _GEN_6525 : _GEN_5825; // @[executor.scala 470:55]
  wire [7:0] _GEN_7362 = opcode_3 != 4'h0 ? _GEN_6530 : _GEN_5826; // @[executor.scala 470:55]
  wire [7:0] _GEN_7363 = opcode_3 != 4'h0 ? _GEN_6531 : _GEN_5827; // @[executor.scala 470:55]
  wire [7:0] _GEN_7364 = opcode_3 != 4'h0 ? _GEN_6532 : _GEN_5828; // @[executor.scala 470:55]
  wire [7:0] _GEN_7365 = opcode_3 != 4'h0 ? _GEN_6533 : _GEN_5829; // @[executor.scala 470:55]
  wire [7:0] _GEN_7366 = opcode_3 != 4'h0 ? _GEN_6538 : _GEN_5830; // @[executor.scala 470:55]
  wire [7:0] _GEN_7367 = opcode_3 != 4'h0 ? _GEN_6539 : _GEN_5831; // @[executor.scala 470:55]
  wire [7:0] _GEN_7368 = opcode_3 != 4'h0 ? _GEN_6540 : _GEN_5832; // @[executor.scala 470:55]
  wire [7:0] _GEN_7369 = opcode_3 != 4'h0 ? _GEN_6541 : _GEN_5833; // @[executor.scala 470:55]
  wire [7:0] _GEN_7370 = opcode_3 != 4'h0 ? _GEN_6546 : _GEN_5834; // @[executor.scala 470:55]
  wire [7:0] _GEN_7371 = opcode_3 != 4'h0 ? _GEN_6547 : _GEN_5835; // @[executor.scala 470:55]
  wire [7:0] _GEN_7372 = opcode_3 != 4'h0 ? _GEN_6548 : _GEN_5836; // @[executor.scala 470:55]
  wire [7:0] _GEN_7373 = opcode_3 != 4'h0 ? _GEN_6549 : _GEN_5837; // @[executor.scala 470:55]
  wire [7:0] _GEN_7374 = opcode_3 != 4'h0 ? _GEN_6554 : _GEN_5838; // @[executor.scala 470:55]
  wire [7:0] _GEN_7375 = opcode_3 != 4'h0 ? _GEN_6555 : _GEN_5839; // @[executor.scala 470:55]
  wire [7:0] _GEN_7376 = opcode_3 != 4'h0 ? _GEN_6556 : _GEN_5840; // @[executor.scala 470:55]
  wire [7:0] _GEN_7377 = opcode_3 != 4'h0 ? _GEN_6557 : _GEN_5841; // @[executor.scala 470:55]
  wire [7:0] _GEN_7378 = opcode_3 != 4'h0 ? _GEN_6562 : _GEN_5842; // @[executor.scala 470:55]
  wire [7:0] _GEN_7379 = opcode_3 != 4'h0 ? _GEN_6563 : _GEN_5843; // @[executor.scala 470:55]
  wire [7:0] _GEN_7380 = opcode_3 != 4'h0 ? _GEN_6564 : _GEN_5844; // @[executor.scala 470:55]
  wire [7:0] _GEN_7381 = opcode_3 != 4'h0 ? _GEN_6565 : _GEN_5845; // @[executor.scala 470:55]
  wire [7:0] _GEN_7382 = opcode_3 != 4'h0 ? _GEN_6570 : _GEN_5846; // @[executor.scala 470:55]
  wire [7:0] _GEN_7383 = opcode_3 != 4'h0 ? _GEN_6571 : _GEN_5847; // @[executor.scala 470:55]
  wire [7:0] _GEN_7384 = opcode_3 != 4'h0 ? _GEN_6572 : _GEN_5848; // @[executor.scala 470:55]
  wire [7:0] _GEN_7385 = opcode_3 != 4'h0 ? _GEN_6573 : _GEN_5849; // @[executor.scala 470:55]
  wire [7:0] _GEN_7386 = opcode_3 != 4'h0 ? _GEN_6578 : _GEN_5850; // @[executor.scala 470:55]
  wire [7:0] _GEN_7387 = opcode_3 != 4'h0 ? _GEN_6579 : _GEN_5851; // @[executor.scala 470:55]
  wire [7:0] _GEN_7388 = opcode_3 != 4'h0 ? _GEN_6580 : _GEN_5852; // @[executor.scala 470:55]
  wire [7:0] _GEN_7389 = opcode_3 != 4'h0 ? _GEN_6581 : _GEN_5853; // @[executor.scala 470:55]
  wire [7:0] _GEN_7390 = opcode_3 != 4'h0 ? _GEN_6586 : _GEN_5854; // @[executor.scala 470:55]
  wire [7:0] _GEN_7391 = opcode_3 != 4'h0 ? _GEN_6587 : _GEN_5855; // @[executor.scala 470:55]
  wire [7:0] _GEN_7392 = opcode_3 != 4'h0 ? _GEN_6588 : _GEN_5856; // @[executor.scala 470:55]
  wire [7:0] _GEN_7393 = opcode_3 != 4'h0 ? _GEN_6589 : _GEN_5857; // @[executor.scala 470:55]
  wire [7:0] _GEN_7394 = opcode_3 != 4'h0 ? _GEN_6594 : _GEN_5858; // @[executor.scala 470:55]
  wire [7:0] _GEN_7395 = opcode_3 != 4'h0 ? _GEN_6595 : _GEN_5859; // @[executor.scala 470:55]
  wire [7:0] _GEN_7396 = opcode_3 != 4'h0 ? _GEN_6596 : _GEN_5860; // @[executor.scala 470:55]
  wire [7:0] _GEN_7397 = opcode_3 != 4'h0 ? _GEN_6597 : _GEN_5861; // @[executor.scala 470:55]
  wire [7:0] _GEN_7398 = opcode_3 != 4'h0 ? _GEN_6602 : _GEN_5862; // @[executor.scala 470:55]
  wire [7:0] _GEN_7399 = opcode_3 != 4'h0 ? _GEN_6603 : _GEN_5863; // @[executor.scala 470:55]
  wire [7:0] _GEN_7400 = opcode_3 != 4'h0 ? _GEN_6604 : _GEN_5864; // @[executor.scala 470:55]
  wire [7:0] _GEN_7401 = opcode_3 != 4'h0 ? _GEN_6605 : _GEN_5865; // @[executor.scala 470:55]
  wire [7:0] _GEN_7402 = opcode_3 != 4'h0 ? _GEN_6610 : _GEN_5866; // @[executor.scala 470:55]
  wire [7:0] _GEN_7403 = opcode_3 != 4'h0 ? _GEN_6611 : _GEN_5867; // @[executor.scala 470:55]
  wire [7:0] _GEN_7404 = opcode_3 != 4'h0 ? _GEN_6612 : _GEN_5868; // @[executor.scala 470:55]
  wire [7:0] _GEN_7405 = opcode_3 != 4'h0 ? _GEN_6613 : _GEN_5869; // @[executor.scala 470:55]
  wire [7:0] _GEN_7406 = opcode_3 != 4'h0 ? _GEN_6618 : _GEN_5870; // @[executor.scala 470:55]
  wire [7:0] _GEN_7407 = opcode_3 != 4'h0 ? _GEN_6619 : _GEN_5871; // @[executor.scala 470:55]
  wire [7:0] _GEN_7408 = opcode_3 != 4'h0 ? _GEN_6620 : _GEN_5872; // @[executor.scala 470:55]
  wire [7:0] _GEN_7409 = opcode_3 != 4'h0 ? _GEN_6621 : _GEN_5873; // @[executor.scala 470:55]
  wire [7:0] _GEN_7410 = opcode_3 != 4'h0 ? _GEN_6626 : _GEN_5874; // @[executor.scala 470:55]
  wire [7:0] _GEN_7411 = opcode_3 != 4'h0 ? _GEN_6627 : _GEN_5875; // @[executor.scala 470:55]
  wire [7:0] _GEN_7412 = opcode_3 != 4'h0 ? _GEN_6628 : _GEN_5876; // @[executor.scala 470:55]
  wire [7:0] _GEN_7413 = opcode_3 != 4'h0 ? _GEN_6629 : _GEN_5877; // @[executor.scala 470:55]
  wire [7:0] _GEN_7414 = opcode_3 != 4'h0 ? _GEN_6634 : _GEN_5878; // @[executor.scala 470:55]
  wire [7:0] _GEN_7415 = opcode_3 != 4'h0 ? _GEN_6635 : _GEN_5879; // @[executor.scala 470:55]
  wire [7:0] _GEN_7416 = opcode_3 != 4'h0 ? _GEN_6636 : _GEN_5880; // @[executor.scala 470:55]
  wire [7:0] _GEN_7417 = opcode_3 != 4'h0 ? _GEN_6637 : _GEN_5881; // @[executor.scala 470:55]
  wire [7:0] _GEN_7418 = opcode_3 != 4'h0 ? _GEN_6642 : _GEN_5882; // @[executor.scala 470:55]
  wire [7:0] _GEN_7419 = opcode_3 != 4'h0 ? _GEN_6643 : _GEN_5883; // @[executor.scala 470:55]
  wire [7:0] _GEN_7420 = opcode_3 != 4'h0 ? _GEN_6644 : _GEN_5884; // @[executor.scala 470:55]
  wire [7:0] _GEN_7421 = opcode_3 != 4'h0 ? _GEN_6645 : _GEN_5885; // @[executor.scala 470:55]
  wire [7:0] _GEN_7422 = opcode_3 != 4'h0 ? _GEN_6650 : _GEN_5886; // @[executor.scala 470:55]
  wire [7:0] _GEN_7423 = opcode_3 != 4'h0 ? _GEN_6651 : _GEN_5887; // @[executor.scala 470:55]
  wire [7:0] _GEN_7424 = opcode_3 != 4'h0 ? _GEN_6652 : _GEN_5888; // @[executor.scala 470:55]
  wire [7:0] _GEN_7425 = opcode_3 != 4'h0 ? _GEN_6653 : _GEN_5889; // @[executor.scala 470:55]
  wire [7:0] _GEN_7426 = opcode_3 != 4'h0 ? _GEN_6658 : _GEN_5890; // @[executor.scala 470:55]
  wire [7:0] _GEN_7427 = opcode_3 != 4'h0 ? _GEN_6659 : _GEN_5891; // @[executor.scala 470:55]
  wire [7:0] _GEN_7428 = opcode_3 != 4'h0 ? _GEN_6660 : _GEN_5892; // @[executor.scala 470:55]
  wire [7:0] _GEN_7429 = opcode_3 != 4'h0 ? _GEN_6661 : _GEN_5893; // @[executor.scala 470:55]
  wire [7:0] _GEN_7430 = opcode_3 != 4'h0 ? _GEN_6666 : _GEN_5894; // @[executor.scala 470:55]
  wire [7:0] _GEN_7431 = opcode_3 != 4'h0 ? _GEN_6667 : _GEN_5895; // @[executor.scala 470:55]
  wire [7:0] _GEN_7432 = opcode_3 != 4'h0 ? _GEN_6668 : _GEN_5896; // @[executor.scala 470:55]
  wire [7:0] _GEN_7433 = opcode_3 != 4'h0 ? _GEN_6669 : _GEN_5897; // @[executor.scala 470:55]
  wire [7:0] _GEN_7434 = opcode_3 != 4'h0 ? _GEN_6674 : _GEN_5898; // @[executor.scala 470:55]
  wire [7:0] _GEN_7435 = opcode_3 != 4'h0 ? _GEN_6675 : _GEN_5899; // @[executor.scala 470:55]
  wire [7:0] _GEN_7436 = opcode_3 != 4'h0 ? _GEN_6676 : _GEN_5900; // @[executor.scala 470:55]
  wire [7:0] _GEN_7437 = opcode_3 != 4'h0 ? _GEN_6677 : _GEN_5901; // @[executor.scala 470:55]
  wire [7:0] _GEN_7438 = opcode_3 != 4'h0 ? _GEN_6682 : _GEN_5902; // @[executor.scala 470:55]
  wire [7:0] _GEN_7439 = opcode_3 != 4'h0 ? _GEN_6683 : _GEN_5903; // @[executor.scala 470:55]
  wire [7:0] _GEN_7440 = opcode_3 != 4'h0 ? _GEN_6684 : _GEN_5904; // @[executor.scala 470:55]
  wire [7:0] _GEN_7441 = opcode_3 != 4'h0 ? _GEN_6685 : _GEN_5905; // @[executor.scala 470:55]
  wire [7:0] _GEN_7442 = opcode_3 != 4'h0 ? _GEN_6690 : _GEN_5906; // @[executor.scala 470:55]
  wire [7:0] _GEN_7443 = opcode_3 != 4'h0 ? _GEN_6691 : _GEN_5907; // @[executor.scala 470:55]
  wire [7:0] _GEN_7444 = opcode_3 != 4'h0 ? _GEN_6692 : _GEN_5908; // @[executor.scala 470:55]
  wire [7:0] _GEN_7445 = opcode_3 != 4'h0 ? _GEN_6693 : _GEN_5909; // @[executor.scala 470:55]
  wire [7:0] _GEN_7446 = opcode_3 != 4'h0 ? _GEN_6698 : _GEN_5910; // @[executor.scala 470:55]
  wire [7:0] _GEN_7447 = opcode_3 != 4'h0 ? _GEN_6699 : _GEN_5911; // @[executor.scala 470:55]
  wire [7:0] _GEN_7448 = opcode_3 != 4'h0 ? _GEN_6700 : _GEN_5912; // @[executor.scala 470:55]
  wire [7:0] _GEN_7449 = opcode_3 != 4'h0 ? _GEN_6701 : _GEN_5913; // @[executor.scala 470:55]
  wire [7:0] _GEN_7450 = opcode_3 != 4'h0 ? _GEN_6706 : _GEN_5914; // @[executor.scala 470:55]
  wire [7:0] _GEN_7451 = opcode_3 != 4'h0 ? _GEN_6707 : _GEN_5915; // @[executor.scala 470:55]
  wire [7:0] _GEN_7452 = opcode_3 != 4'h0 ? _GEN_6708 : _GEN_5916; // @[executor.scala 470:55]
  wire [7:0] _GEN_7453 = opcode_3 != 4'h0 ? _GEN_6709 : _GEN_5917; // @[executor.scala 470:55]
  wire [7:0] _GEN_7454 = opcode_3 != 4'h0 ? _GEN_6714 : _GEN_5918; // @[executor.scala 470:55]
  wire [7:0] _GEN_7455 = opcode_3 != 4'h0 ? _GEN_6715 : _GEN_5919; // @[executor.scala 470:55]
  wire [7:0] _GEN_7456 = opcode_3 != 4'h0 ? _GEN_6716 : _GEN_5920; // @[executor.scala 470:55]
  wire [7:0] _GEN_7457 = opcode_3 != 4'h0 ? _GEN_6717 : _GEN_5921; // @[executor.scala 470:55]
  wire [7:0] _GEN_7458 = opcode_3 != 4'h0 ? _GEN_6722 : _GEN_5922; // @[executor.scala 470:55]
  wire [7:0] _GEN_7459 = opcode_3 != 4'h0 ? _GEN_6723 : _GEN_5923; // @[executor.scala 470:55]
  wire [7:0] _GEN_7460 = opcode_3 != 4'h0 ? _GEN_6724 : _GEN_5924; // @[executor.scala 470:55]
  wire [7:0] _GEN_7461 = opcode_3 != 4'h0 ? _GEN_6725 : _GEN_5925; // @[executor.scala 470:55]
  wire [7:0] _GEN_7462 = opcode_3 != 4'h0 ? _GEN_6730 : _GEN_5926; // @[executor.scala 470:55]
  wire [7:0] _GEN_7463 = opcode_3 != 4'h0 ? _GEN_6731 : _GEN_5927; // @[executor.scala 470:55]
  wire [7:0] _GEN_7464 = opcode_3 != 4'h0 ? _GEN_6732 : _GEN_5928; // @[executor.scala 470:55]
  wire [7:0] _GEN_7465 = opcode_3 != 4'h0 ? _GEN_6733 : _GEN_5929; // @[executor.scala 470:55]
  wire [7:0] _GEN_7466 = opcode_3 != 4'h0 ? _GEN_6738 : _GEN_5930; // @[executor.scala 470:55]
  wire [7:0] _GEN_7467 = opcode_3 != 4'h0 ? _GEN_6739 : _GEN_5931; // @[executor.scala 470:55]
  wire [7:0] _GEN_7468 = opcode_3 != 4'h0 ? _GEN_6740 : _GEN_5932; // @[executor.scala 470:55]
  wire [7:0] _GEN_7469 = opcode_3 != 4'h0 ? _GEN_6741 : _GEN_5933; // @[executor.scala 470:55]
  wire [7:0] _GEN_7470 = opcode_3 != 4'h0 ? _GEN_6746 : _GEN_5934; // @[executor.scala 470:55]
  wire [7:0] _GEN_7471 = opcode_3 != 4'h0 ? _GEN_6747 : _GEN_5935; // @[executor.scala 470:55]
  wire [7:0] _GEN_7472 = opcode_3 != 4'h0 ? _GEN_6748 : _GEN_5936; // @[executor.scala 470:55]
  wire [7:0] _GEN_7473 = opcode_3 != 4'h0 ? _GEN_6749 : _GEN_5937; // @[executor.scala 470:55]
  wire [7:0] _GEN_7474 = opcode_3 != 4'h0 ? _GEN_6754 : _GEN_5938; // @[executor.scala 470:55]
  wire [7:0] _GEN_7475 = opcode_3 != 4'h0 ? _GEN_6755 : _GEN_5939; // @[executor.scala 470:55]
  wire [7:0] _GEN_7476 = opcode_3 != 4'h0 ? _GEN_6756 : _GEN_5940; // @[executor.scala 470:55]
  wire [7:0] _GEN_7477 = opcode_3 != 4'h0 ? _GEN_6757 : _GEN_5941; // @[executor.scala 470:55]
  wire [7:0] _GEN_7478 = opcode_3 != 4'h0 ? _GEN_6762 : _GEN_5942; // @[executor.scala 470:55]
  wire [7:0] _GEN_7479 = opcode_3 != 4'h0 ? _GEN_6763 : _GEN_5943; // @[executor.scala 470:55]
  wire [7:0] _GEN_7480 = opcode_3 != 4'h0 ? _GEN_6764 : _GEN_5944; // @[executor.scala 470:55]
  wire [7:0] _GEN_7481 = opcode_3 != 4'h0 ? _GEN_6765 : _GEN_5945; // @[executor.scala 470:55]
  wire [7:0] _GEN_7482 = opcode_3 != 4'h0 ? _GEN_6770 : _GEN_5946; // @[executor.scala 470:55]
  wire [7:0] _GEN_7483 = opcode_3 != 4'h0 ? _GEN_6771 : _GEN_5947; // @[executor.scala 470:55]
  wire [7:0] _GEN_7484 = opcode_3 != 4'h0 ? _GEN_6772 : _GEN_5948; // @[executor.scala 470:55]
  wire [7:0] _GEN_7485 = opcode_3 != 4'h0 ? _GEN_6773 : _GEN_5949; // @[executor.scala 470:55]
  wire [7:0] _GEN_7486 = opcode_3 != 4'h0 ? _GEN_6778 : _GEN_5950; // @[executor.scala 470:55]
  wire [7:0] _GEN_7487 = opcode_3 != 4'h0 ? _GEN_6779 : _GEN_5951; // @[executor.scala 470:55]
  wire [7:0] _GEN_7488 = opcode_3 != 4'h0 ? _GEN_6780 : _GEN_5952; // @[executor.scala 470:55]
  wire [7:0] _GEN_7489 = opcode_3 != 4'h0 ? _GEN_6781 : _GEN_5953; // @[executor.scala 470:55]
  wire [7:0] _GEN_7490 = opcode_3 != 4'h0 ? _GEN_6786 : _GEN_5954; // @[executor.scala 470:55]
  wire [7:0] _GEN_7491 = opcode_3 != 4'h0 ? _GEN_6787 : _GEN_5955; // @[executor.scala 470:55]
  wire [7:0] _GEN_7492 = opcode_3 != 4'h0 ? _GEN_6788 : _GEN_5956; // @[executor.scala 470:55]
  wire [7:0] _GEN_7493 = opcode_3 != 4'h0 ? _GEN_6789 : _GEN_5957; // @[executor.scala 470:55]
  wire [7:0] _GEN_7494 = opcode_3 != 4'h0 ? _GEN_6794 : _GEN_5958; // @[executor.scala 470:55]
  wire [7:0] _GEN_7495 = opcode_3 != 4'h0 ? _GEN_6795 : _GEN_5959; // @[executor.scala 470:55]
  wire [7:0] _GEN_7496 = opcode_3 != 4'h0 ? _GEN_6796 : _GEN_5960; // @[executor.scala 470:55]
  wire [7:0] _GEN_7497 = opcode_3 != 4'h0 ? _GEN_6797 : _GEN_5961; // @[executor.scala 470:55]
  wire [7:0] _GEN_7498 = opcode_3 != 4'h0 ? _GEN_6802 : _GEN_5962; // @[executor.scala 470:55]
  wire [7:0] _GEN_7499 = opcode_3 != 4'h0 ? _GEN_6803 : _GEN_5963; // @[executor.scala 470:55]
  wire [7:0] _GEN_7500 = opcode_3 != 4'h0 ? _GEN_6804 : _GEN_5964; // @[executor.scala 470:55]
  wire [7:0] _GEN_7501 = opcode_3 != 4'h0 ? _GEN_6805 : _GEN_5965; // @[executor.scala 470:55]
  wire [7:0] _GEN_7502 = opcode_3 != 4'h0 ? _GEN_6810 : _GEN_5966; // @[executor.scala 470:55]
  wire [7:0] _GEN_7503 = opcode_3 != 4'h0 ? _GEN_6811 : _GEN_5967; // @[executor.scala 470:55]
  wire [7:0] _GEN_7504 = opcode_3 != 4'h0 ? _GEN_6812 : _GEN_5968; // @[executor.scala 470:55]
  wire [7:0] _GEN_7505 = opcode_3 != 4'h0 ? _GEN_6813 : _GEN_5969; // @[executor.scala 470:55]
  wire [7:0] _GEN_7506 = opcode_3 != 4'h0 ? _GEN_6818 : _GEN_5970; // @[executor.scala 470:55]
  wire [7:0] _GEN_7507 = opcode_3 != 4'h0 ? _GEN_6819 : _GEN_5971; // @[executor.scala 470:55]
  wire [7:0] _GEN_7508 = opcode_3 != 4'h0 ? _GEN_6820 : _GEN_5972; // @[executor.scala 470:55]
  wire [7:0] _GEN_7509 = opcode_3 != 4'h0 ? _GEN_6821 : _GEN_5973; // @[executor.scala 470:55]
  wire [7:0] _GEN_7510 = opcode_3 != 4'h0 ? _GEN_6826 : _GEN_5974; // @[executor.scala 470:55]
  wire [7:0] _GEN_7511 = opcode_3 != 4'h0 ? _GEN_6827 : _GEN_5975; // @[executor.scala 470:55]
  wire [7:0] _GEN_7512 = opcode_3 != 4'h0 ? _GEN_6828 : _GEN_5976; // @[executor.scala 470:55]
  wire [7:0] _GEN_7513 = opcode_3 != 4'h0 ? _GEN_6829 : _GEN_5977; // @[executor.scala 470:55]
  wire [7:0] _GEN_7514 = opcode_3 != 4'h0 ? _GEN_6834 : _GEN_5978; // @[executor.scala 470:55]
  wire [7:0] _GEN_7515 = opcode_3 != 4'h0 ? _GEN_6835 : _GEN_5979; // @[executor.scala 470:55]
  wire [7:0] _GEN_7516 = opcode_3 != 4'h0 ? _GEN_6836 : _GEN_5980; // @[executor.scala 470:55]
  wire [7:0] _GEN_7517 = opcode_3 != 4'h0 ? _GEN_6837 : _GEN_5981; // @[executor.scala 470:55]
  wire [7:0] _GEN_7518 = opcode_3 != 4'h0 ? _GEN_6842 : _GEN_5982; // @[executor.scala 470:55]
  wire [7:0] _GEN_7519 = opcode_3 != 4'h0 ? _GEN_6843 : _GEN_5983; // @[executor.scala 470:55]
  wire [7:0] _GEN_7520 = opcode_3 != 4'h0 ? _GEN_6844 : _GEN_5984; // @[executor.scala 470:55]
  wire [7:0] _GEN_7521 = opcode_3 != 4'h0 ? _GEN_6845 : _GEN_5985; // @[executor.scala 470:55]
  wire [7:0] _GEN_7522 = opcode_3 != 4'h0 ? _GEN_6850 : _GEN_5986; // @[executor.scala 470:55]
  wire [7:0] _GEN_7523 = opcode_3 != 4'h0 ? _GEN_6851 : _GEN_5987; // @[executor.scala 470:55]
  wire [7:0] _GEN_7524 = opcode_3 != 4'h0 ? _GEN_6852 : _GEN_5988; // @[executor.scala 470:55]
  wire [7:0] _GEN_7525 = opcode_3 != 4'h0 ? _GEN_6853 : _GEN_5989; // @[executor.scala 470:55]
  wire [7:0] _GEN_7526 = opcode_3 != 4'h0 ? _GEN_6858 : _GEN_5990; // @[executor.scala 470:55]
  wire [7:0] _GEN_7527 = opcode_3 != 4'h0 ? _GEN_6859 : _GEN_5991; // @[executor.scala 470:55]
  wire [7:0] _GEN_7528 = opcode_3 != 4'h0 ? _GEN_6860 : _GEN_5992; // @[executor.scala 470:55]
  wire [7:0] _GEN_7529 = opcode_3 != 4'h0 ? _GEN_6861 : _GEN_5993; // @[executor.scala 470:55]
  wire [7:0] _GEN_7530 = opcode_3 != 4'h0 ? _GEN_6866 : _GEN_5994; // @[executor.scala 470:55]
  wire [7:0] _GEN_7531 = opcode_3 != 4'h0 ? _GEN_6867 : _GEN_5995; // @[executor.scala 470:55]
  wire [7:0] _GEN_7532 = opcode_3 != 4'h0 ? _GEN_6868 : _GEN_5996; // @[executor.scala 470:55]
  wire [7:0] _GEN_7533 = opcode_3 != 4'h0 ? _GEN_6869 : _GEN_5997; // @[executor.scala 470:55]
  wire [7:0] _GEN_7534 = opcode_3 != 4'h0 ? _GEN_6874 : _GEN_5998; // @[executor.scala 470:55]
  wire [7:0] _GEN_7535 = opcode_3 != 4'h0 ? _GEN_6875 : _GEN_5999; // @[executor.scala 470:55]
  wire [7:0] _GEN_7536 = opcode_3 != 4'h0 ? _GEN_6876 : _GEN_6000; // @[executor.scala 470:55]
  wire [7:0] _GEN_7537 = opcode_3 != 4'h0 ? _GEN_6877 : _GEN_6001; // @[executor.scala 470:55]
  wire [7:0] _GEN_7538 = opcode_3 != 4'h0 ? _GEN_6882 : _GEN_6002; // @[executor.scala 470:55]
  wire [7:0] _GEN_7539 = opcode_3 != 4'h0 ? _GEN_6883 : _GEN_6003; // @[executor.scala 470:55]
  wire [7:0] _GEN_7540 = opcode_3 != 4'h0 ? _GEN_6884 : _GEN_6004; // @[executor.scala 470:55]
  wire [7:0] _GEN_7541 = opcode_3 != 4'h0 ? _GEN_6885 : _GEN_6005; // @[executor.scala 470:55]
  wire [7:0] _GEN_7542 = opcode_3 != 4'h0 ? _GEN_6890 : _GEN_6006; // @[executor.scala 470:55]
  wire [7:0] _GEN_7543 = opcode_3 != 4'h0 ? _GEN_6891 : _GEN_6007; // @[executor.scala 470:55]
  wire [7:0] _GEN_7544 = opcode_3 != 4'h0 ? _GEN_6892 : _GEN_6008; // @[executor.scala 470:55]
  wire [7:0] _GEN_7545 = opcode_3 != 4'h0 ? _GEN_6893 : _GEN_6009; // @[executor.scala 470:55]
  wire [7:0] _GEN_7546 = opcode_3 != 4'h0 ? _GEN_6898 : _GEN_6010; // @[executor.scala 470:55]
  wire [7:0] _GEN_7547 = opcode_3 != 4'h0 ? _GEN_6899 : _GEN_6011; // @[executor.scala 470:55]
  wire [7:0] _GEN_7548 = opcode_3 != 4'h0 ? _GEN_6900 : _GEN_6012; // @[executor.scala 470:55]
  wire [7:0] _GEN_7549 = opcode_3 != 4'h0 ? _GEN_6901 : _GEN_6013; // @[executor.scala 470:55]
  wire [7:0] _GEN_7550 = opcode_3 != 4'h0 ? _GEN_6906 : _GEN_6014; // @[executor.scala 470:55]
  wire [7:0] _GEN_7551 = opcode_3 != 4'h0 ? _GEN_6907 : _GEN_6015; // @[executor.scala 470:55]
  wire [7:0] _GEN_7552 = opcode_3 != 4'h0 ? _GEN_6908 : _GEN_6016; // @[executor.scala 470:55]
  wire [7:0] _GEN_7553 = opcode_3 != 4'h0 ? _GEN_6909 : _GEN_6017; // @[executor.scala 470:55]
  wire [7:0] _GEN_7554 = opcode_3 != 4'h0 ? _GEN_6914 : _GEN_6018; // @[executor.scala 470:55]
  wire [7:0] _GEN_7555 = opcode_3 != 4'h0 ? _GEN_6915 : _GEN_6019; // @[executor.scala 470:55]
  wire [7:0] _GEN_7556 = opcode_3 != 4'h0 ? _GEN_6916 : _GEN_6020; // @[executor.scala 470:55]
  wire [7:0] _GEN_7557 = opcode_3 != 4'h0 ? _GEN_6917 : _GEN_6021; // @[executor.scala 470:55]
  wire [7:0] _GEN_7558 = opcode_3 != 4'h0 ? _GEN_6922 : _GEN_6022; // @[executor.scala 470:55]
  wire [7:0] _GEN_7559 = opcode_3 != 4'h0 ? _GEN_6923 : _GEN_6023; // @[executor.scala 470:55]
  wire [7:0] _GEN_7560 = opcode_3 != 4'h0 ? _GEN_6924 : _GEN_6024; // @[executor.scala 470:55]
  wire [7:0] _GEN_7561 = opcode_3 != 4'h0 ? _GEN_6925 : _GEN_6025; // @[executor.scala 470:55]
  wire [7:0] _GEN_7562 = opcode_3 != 4'h0 ? _GEN_6930 : _GEN_6026; // @[executor.scala 470:55]
  wire [7:0] _GEN_7563 = opcode_3 != 4'h0 ? _GEN_6931 : _GEN_6027; // @[executor.scala 470:55]
  wire [7:0] _GEN_7564 = opcode_3 != 4'h0 ? _GEN_6932 : _GEN_6028; // @[executor.scala 470:55]
  wire [7:0] _GEN_7565 = opcode_3 != 4'h0 ? _GEN_6933 : _GEN_6029; // @[executor.scala 470:55]
  wire [7:0] _GEN_7566 = opcode_3 != 4'h0 ? _GEN_6938 : _GEN_6030; // @[executor.scala 470:55]
  wire [7:0] _GEN_7567 = opcode_3 != 4'h0 ? _GEN_6939 : _GEN_6031; // @[executor.scala 470:55]
  wire [7:0] _GEN_7568 = opcode_3 != 4'h0 ? _GEN_6940 : _GEN_6032; // @[executor.scala 470:55]
  wire [7:0] _GEN_7569 = opcode_3 != 4'h0 ? _GEN_6941 : _GEN_6033; // @[executor.scala 470:55]
  wire [7:0] _GEN_7570 = opcode_3 != 4'h0 ? _GEN_6946 : _GEN_6034; // @[executor.scala 470:55]
  wire [7:0] _GEN_7571 = opcode_3 != 4'h0 ? _GEN_6947 : _GEN_6035; // @[executor.scala 470:55]
  wire [7:0] _GEN_7572 = opcode_3 != 4'h0 ? _GEN_6948 : _GEN_6036; // @[executor.scala 470:55]
  wire [7:0] _GEN_7573 = opcode_3 != 4'h0 ? _GEN_6949 : _GEN_6037; // @[executor.scala 470:55]
  wire [7:0] _GEN_7574 = opcode_3 != 4'h0 ? _GEN_6954 : _GEN_6038; // @[executor.scala 470:55]
  wire [7:0] _GEN_7575 = opcode_3 != 4'h0 ? _GEN_6955 : _GEN_6039; // @[executor.scala 470:55]
  wire [7:0] _GEN_7576 = opcode_3 != 4'h0 ? _GEN_6956 : _GEN_6040; // @[executor.scala 470:55]
  wire [7:0] _GEN_7577 = opcode_3 != 4'h0 ? _GEN_6957 : _GEN_6041; // @[executor.scala 470:55]
  wire [7:0] _GEN_7578 = opcode_3 != 4'h0 ? _GEN_6962 : _GEN_6042; // @[executor.scala 470:55]
  wire [7:0] _GEN_7579 = opcode_3 != 4'h0 ? _GEN_6963 : _GEN_6043; // @[executor.scala 470:55]
  wire [7:0] _GEN_7580 = opcode_3 != 4'h0 ? _GEN_6964 : _GEN_6044; // @[executor.scala 470:55]
  wire [7:0] _GEN_7581 = opcode_3 != 4'h0 ? _GEN_6965 : _GEN_6045; // @[executor.scala 470:55]
  wire [7:0] _GEN_7582 = opcode_3 != 4'h0 ? _GEN_6970 : _GEN_6046; // @[executor.scala 470:55]
  wire [7:0] _GEN_7583 = opcode_3 != 4'h0 ? _GEN_6971 : _GEN_6047; // @[executor.scala 470:55]
  wire [7:0] _GEN_7584 = opcode_3 != 4'h0 ? _GEN_6972 : _GEN_6048; // @[executor.scala 470:55]
  wire [7:0] _GEN_7585 = opcode_3 != 4'h0 ? _GEN_6973 : _GEN_6049; // @[executor.scala 470:55]
  wire [7:0] _GEN_7586 = opcode_3 != 4'h0 ? _GEN_6978 : _GEN_6050; // @[executor.scala 470:55]
  wire [7:0] _GEN_7587 = opcode_3 != 4'h0 ? _GEN_6979 : _GEN_6051; // @[executor.scala 470:55]
  wire [7:0] _GEN_7588 = opcode_3 != 4'h0 ? _GEN_6980 : _GEN_6052; // @[executor.scala 470:55]
  wire [7:0] _GEN_7589 = opcode_3 != 4'h0 ? _GEN_6981 : _GEN_6053; // @[executor.scala 470:55]
  wire [7:0] _GEN_7590 = opcode_3 != 4'h0 ? _GEN_6986 : _GEN_6054; // @[executor.scala 470:55]
  wire [7:0] _GEN_7591 = opcode_3 != 4'h0 ? _GEN_6987 : _GEN_6055; // @[executor.scala 470:55]
  wire [7:0] _GEN_7592 = opcode_3 != 4'h0 ? _GEN_6988 : _GEN_6056; // @[executor.scala 470:55]
  wire [7:0] _GEN_7593 = opcode_3 != 4'h0 ? _GEN_6989 : _GEN_6057; // @[executor.scala 470:55]
  wire [7:0] _GEN_7594 = opcode_3 != 4'h0 ? _GEN_6994 : _GEN_6058; // @[executor.scala 470:55]
  wire [7:0] _GEN_7595 = opcode_3 != 4'h0 ? _GEN_6995 : _GEN_6059; // @[executor.scala 470:55]
  wire [7:0] _GEN_7596 = opcode_3 != 4'h0 ? _GEN_6996 : _GEN_6060; // @[executor.scala 470:55]
  wire [7:0] _GEN_7597 = opcode_3 != 4'h0 ? _GEN_6997 : _GEN_6061; // @[executor.scala 470:55]
  wire [7:0] _GEN_7598 = opcode_3 != 4'h0 ? _GEN_7002 : _GEN_6062; // @[executor.scala 470:55]
  wire [7:0] _GEN_7599 = opcode_3 != 4'h0 ? _GEN_7003 : _GEN_6063; // @[executor.scala 470:55]
  wire [7:0] _GEN_7600 = opcode_3 != 4'h0 ? _GEN_7004 : _GEN_6064; // @[executor.scala 470:55]
  wire [7:0] _GEN_7601 = opcode_3 != 4'h0 ? _GEN_7005 : _GEN_6065; // @[executor.scala 470:55]
  wire [7:0] _GEN_7602 = opcode_3 != 4'h0 ? _GEN_7010 : _GEN_6066; // @[executor.scala 470:55]
  wire [7:0] _GEN_7603 = opcode_3 != 4'h0 ? _GEN_7011 : _GEN_6067; // @[executor.scala 470:55]
  wire [7:0] _GEN_7604 = opcode_3 != 4'h0 ? _GEN_7012 : _GEN_6068; // @[executor.scala 470:55]
  wire [7:0] _GEN_7605 = opcode_3 != 4'h0 ? _GEN_7013 : _GEN_6069; // @[executor.scala 470:55]
  wire [7:0] _GEN_7606 = opcode_3 != 4'h0 ? _GEN_7018 : _GEN_6070; // @[executor.scala 470:55]
  wire [7:0] _GEN_7607 = opcode_3 != 4'h0 ? _GEN_7019 : _GEN_6071; // @[executor.scala 470:55]
  wire [7:0] _GEN_7608 = opcode_3 != 4'h0 ? _GEN_7020 : _GEN_6072; // @[executor.scala 470:55]
  wire [7:0] _GEN_7609 = opcode_3 != 4'h0 ? _GEN_7021 : _GEN_6073; // @[executor.scala 470:55]
  wire [7:0] _GEN_7610 = opcode_3 != 4'h0 ? _GEN_7026 : _GEN_6074; // @[executor.scala 470:55]
  wire [7:0] _GEN_7611 = opcode_3 != 4'h0 ? _GEN_7027 : _GEN_6075; // @[executor.scala 470:55]
  wire [7:0] _GEN_7612 = opcode_3 != 4'h0 ? _GEN_7028 : _GEN_6076; // @[executor.scala 470:55]
  wire [7:0] _GEN_7613 = opcode_3 != 4'h0 ? _GEN_7029 : _GEN_6077; // @[executor.scala 470:55]
  wire [7:0] _GEN_7614 = opcode_3 != 4'h0 ? _GEN_7034 : _GEN_6078; // @[executor.scala 470:55]
  wire [7:0] _GEN_7615 = opcode_3 != 4'h0 ? _GEN_7035 : _GEN_6079; // @[executor.scala 470:55]
  wire [7:0] _GEN_7616 = opcode_3 != 4'h0 ? _GEN_7036 : _GEN_6080; // @[executor.scala 470:55]
  wire [7:0] _GEN_7617 = opcode_3 != 4'h0 ? _GEN_7037 : _GEN_6081; // @[executor.scala 470:55]
  wire [7:0] _GEN_7618 = opcode_3 != 4'h0 ? _GEN_7042 : _GEN_6082; // @[executor.scala 470:55]
  wire [7:0] _GEN_7619 = opcode_3 != 4'h0 ? _GEN_7043 : _GEN_6083; // @[executor.scala 470:55]
  wire [7:0] _GEN_7620 = opcode_3 != 4'h0 ? _GEN_7044 : _GEN_6084; // @[executor.scala 470:55]
  wire [7:0] _GEN_7621 = opcode_3 != 4'h0 ? _GEN_7045 : _GEN_6085; // @[executor.scala 470:55]
  wire [7:0] _GEN_7622 = opcode_3 != 4'h0 ? _GEN_7050 : _GEN_6086; // @[executor.scala 470:55]
  wire [7:0] _GEN_7623 = opcode_3 != 4'h0 ? _GEN_7051 : _GEN_6087; // @[executor.scala 470:55]
  wire [7:0] _GEN_7624 = opcode_3 != 4'h0 ? _GEN_7052 : _GEN_6088; // @[executor.scala 470:55]
  wire [7:0] _GEN_7625 = opcode_3 != 4'h0 ? _GEN_7053 : _GEN_6089; // @[executor.scala 470:55]
  wire [7:0] _GEN_7626 = opcode_3 != 4'h0 ? _GEN_7058 : _GEN_6090; // @[executor.scala 470:55]
  wire [7:0] _GEN_7627 = opcode_3 != 4'h0 ? _GEN_7059 : _GEN_6091; // @[executor.scala 470:55]
  wire [7:0] _GEN_7628 = opcode_3 != 4'h0 ? _GEN_7060 : _GEN_6092; // @[executor.scala 470:55]
  wire [7:0] _GEN_7629 = opcode_3 != 4'h0 ? _GEN_7061 : _GEN_6093; // @[executor.scala 470:55]
  wire [7:0] _GEN_7630 = opcode_3 != 4'h0 ? _GEN_7066 : _GEN_6094; // @[executor.scala 470:55]
  wire [7:0] _GEN_7631 = opcode_3 != 4'h0 ? _GEN_7067 : _GEN_6095; // @[executor.scala 470:55]
  wire [7:0] _GEN_7632 = opcode_3 != 4'h0 ? _GEN_7068 : _GEN_6096; // @[executor.scala 470:55]
  wire [7:0] _GEN_7633 = opcode_3 != 4'h0 ? _GEN_7069 : _GEN_6097; // @[executor.scala 470:55]
  wire [7:0] _GEN_7634 = opcode_3 != 4'h0 ? _GEN_7074 : _GEN_6098; // @[executor.scala 470:55]
  wire [7:0] _GEN_7635 = opcode_3 != 4'h0 ? _GEN_7075 : _GEN_6099; // @[executor.scala 470:55]
  wire [7:0] _GEN_7636 = opcode_3 != 4'h0 ? _GEN_7076 : _GEN_6100; // @[executor.scala 470:55]
  wire [7:0] _GEN_7637 = opcode_3 != 4'h0 ? _GEN_7077 : _GEN_6101; // @[executor.scala 470:55]
  wire [7:0] _GEN_7638 = opcode_3 != 4'h0 ? _GEN_7082 : _GEN_6102; // @[executor.scala 470:55]
  wire [7:0] _GEN_7639 = opcode_3 != 4'h0 ? _GEN_7083 : _GEN_6103; // @[executor.scala 470:55]
  wire [7:0] _GEN_7640 = opcode_3 != 4'h0 ? _GEN_7084 : _GEN_6104; // @[executor.scala 470:55]
  wire [7:0] _GEN_7641 = opcode_3 != 4'h0 ? _GEN_7085 : _GEN_6105; // @[executor.scala 470:55]
  wire [7:0] _GEN_7642 = opcode_3 != 4'h0 ? _GEN_7090 : _GEN_6106; // @[executor.scala 470:55]
  wire [7:0] _GEN_7643 = opcode_3 != 4'h0 ? _GEN_7091 : _GEN_6107; // @[executor.scala 470:55]
  wire [7:0] _GEN_7644 = opcode_3 != 4'h0 ? _GEN_7092 : _GEN_6108; // @[executor.scala 470:55]
  wire [7:0] _GEN_7645 = opcode_3 != 4'h0 ? _GEN_7093 : _GEN_6109; // @[executor.scala 470:55]
  wire [7:0] _GEN_7646 = opcode_3 != 4'h0 ? _GEN_7098 : _GEN_6110; // @[executor.scala 470:55]
  wire [7:0] _GEN_7647 = opcode_3 != 4'h0 ? _GEN_7099 : _GEN_6111; // @[executor.scala 470:55]
  wire [7:0] _GEN_7648 = opcode_3 != 4'h0 ? _GEN_7100 : _GEN_6112; // @[executor.scala 470:55]
  wire [7:0] _GEN_7649 = opcode_3 != 4'h0 ? _GEN_7101 : _GEN_6113; // @[executor.scala 470:55]
  wire [7:0] _GEN_7650 = opcode_3 != 4'h0 ? _GEN_7106 : _GEN_6114; // @[executor.scala 470:55]
  wire [7:0] _GEN_7651 = opcode_3 != 4'h0 ? _GEN_7107 : _GEN_6115; // @[executor.scala 470:55]
  wire [7:0] _GEN_7652 = opcode_3 != 4'h0 ? _GEN_7108 : _GEN_6116; // @[executor.scala 470:55]
  wire [7:0] _GEN_7653 = opcode_3 != 4'h0 ? _GEN_7109 : _GEN_6117; // @[executor.scala 470:55]
  wire [7:0] _GEN_7654 = opcode_3 != 4'h0 ? _GEN_7114 : _GEN_6118; // @[executor.scala 470:55]
  wire [7:0] _GEN_7655 = opcode_3 != 4'h0 ? _GEN_7115 : _GEN_6119; // @[executor.scala 470:55]
  wire [7:0] _GEN_7656 = opcode_3 != 4'h0 ? _GEN_7116 : _GEN_6120; // @[executor.scala 470:55]
  wire [7:0] _GEN_7657 = opcode_3 != 4'h0 ? _GEN_7117 : _GEN_6121; // @[executor.scala 470:55]
  wire [7:0] _GEN_7658 = opcode_3 != 4'h0 ? _GEN_7122 : _GEN_6122; // @[executor.scala 470:55]
  wire [7:0] _GEN_7659 = opcode_3 != 4'h0 ? _GEN_7123 : _GEN_6123; // @[executor.scala 470:55]
  wire [7:0] _GEN_7660 = opcode_3 != 4'h0 ? _GEN_7124 : _GEN_6124; // @[executor.scala 470:55]
  wire [7:0] _GEN_7661 = opcode_3 != 4'h0 ? _GEN_7125 : _GEN_6125; // @[executor.scala 470:55]
  wire [7:0] _GEN_7662 = opcode_3 != 4'h0 ? _GEN_7130 : _GEN_6126; // @[executor.scala 470:55]
  wire [7:0] _GEN_7663 = opcode_3 != 4'h0 ? _GEN_7131 : _GEN_6127; // @[executor.scala 470:55]
  wire [7:0] _GEN_7664 = opcode_3 != 4'h0 ? _GEN_7132 : _GEN_6128; // @[executor.scala 470:55]
  wire [7:0] _GEN_7665 = opcode_3 != 4'h0 ? _GEN_7133 : _GEN_6129; // @[executor.scala 470:55]
  wire [7:0] _GEN_7666 = opcode_3 != 4'h0 ? _GEN_7138 : _GEN_6130; // @[executor.scala 470:55]
  wire [7:0] _GEN_7667 = opcode_3 != 4'h0 ? _GEN_7139 : _GEN_6131; // @[executor.scala 470:55]
  wire [7:0] _GEN_7668 = opcode_3 != 4'h0 ? _GEN_7140 : _GEN_6132; // @[executor.scala 470:55]
  wire [7:0] _GEN_7669 = opcode_3 != 4'h0 ? _GEN_7141 : _GEN_6133; // @[executor.scala 470:55]
  wire [7:0] _GEN_7670 = opcode_3 != 4'h0 ? _GEN_7146 : _GEN_6134; // @[executor.scala 470:55]
  wire [7:0] _GEN_7671 = opcode_3 != 4'h0 ? _GEN_7147 : _GEN_6135; // @[executor.scala 470:55]
  wire [7:0] _GEN_7672 = opcode_3 != 4'h0 ? _GEN_7148 : _GEN_6136; // @[executor.scala 470:55]
  wire [7:0] _GEN_7673 = opcode_3 != 4'h0 ? _GEN_7149 : _GEN_6137; // @[executor.scala 470:55]
  wire [7:0] _GEN_7674 = opcode_3 != 4'h0 ? _GEN_7154 : _GEN_6138; // @[executor.scala 470:55]
  wire [7:0] _GEN_7675 = opcode_3 != 4'h0 ? _GEN_7155 : _GEN_6139; // @[executor.scala 470:55]
  wire [7:0] _GEN_7676 = opcode_3 != 4'h0 ? _GEN_7156 : _GEN_6140; // @[executor.scala 470:55]
  wire [7:0] _GEN_7677 = opcode_3 != 4'h0 ? _GEN_7157 : _GEN_6141; // @[executor.scala 470:55]
  wire [7:0] _GEN_7678 = opcode_3 != 4'h0 ? _GEN_7162 : _GEN_6142; // @[executor.scala 470:55]
  wire [7:0] _GEN_7679 = opcode_3 != 4'h0 ? _GEN_7163 : _GEN_6143; // @[executor.scala 470:55]
  wire [7:0] _GEN_7680 = opcode_3 != 4'h0 ? _GEN_7164 : _GEN_6144; // @[executor.scala 470:55]
  wire [7:0] _GEN_7681 = opcode_3 != 4'h0 ? _GEN_7165 : _GEN_6145; // @[executor.scala 470:55]
  wire [7:0] _GEN_7682 = opcode_3 != 4'h0 ? _GEN_7170 : _GEN_6146; // @[executor.scala 470:55]
  wire [7:0] _GEN_7683 = opcode_3 != 4'h0 ? _GEN_7171 : _GEN_6147; // @[executor.scala 470:55]
  wire [7:0] _GEN_7684 = opcode_3 != 4'h0 ? _GEN_7172 : _GEN_6148; // @[executor.scala 470:55]
  wire [7:0] _GEN_7685 = opcode_3 != 4'h0 ? _GEN_7173 : _GEN_6149; // @[executor.scala 470:55]
  wire [3:0] _GEN_7686 = opcode_3 == 4'hf ? parameter_2_3[13:10] : _GEN_5636; // @[executor.scala 466:52 executor.scala 467:55]
  wire  _GEN_7687 = opcode_3 == 4'hf ? parameter_2_3[0] : _GEN_5637; // @[executor.scala 466:52 executor.scala 468:55]
  wire [7:0] _GEN_7688 = opcode_3 == 4'hf ? _GEN_5638 : _GEN_7174; // @[executor.scala 466:52]
  wire [7:0] _GEN_7689 = opcode_3 == 4'hf ? _GEN_5639 : _GEN_7175; // @[executor.scala 466:52]
  wire [7:0] _GEN_7690 = opcode_3 == 4'hf ? _GEN_5640 : _GEN_7176; // @[executor.scala 466:52]
  wire [7:0] _GEN_7691 = opcode_3 == 4'hf ? _GEN_5641 : _GEN_7177; // @[executor.scala 466:52]
  wire [7:0] _GEN_7692 = opcode_3 == 4'hf ? _GEN_5642 : _GEN_7178; // @[executor.scala 466:52]
  wire [7:0] _GEN_7693 = opcode_3 == 4'hf ? _GEN_5643 : _GEN_7179; // @[executor.scala 466:52]
  wire [7:0] _GEN_7694 = opcode_3 == 4'hf ? _GEN_5644 : _GEN_7180; // @[executor.scala 466:52]
  wire [7:0] _GEN_7695 = opcode_3 == 4'hf ? _GEN_5645 : _GEN_7181; // @[executor.scala 466:52]
  wire [7:0] _GEN_7696 = opcode_3 == 4'hf ? _GEN_5646 : _GEN_7182; // @[executor.scala 466:52]
  wire [7:0] _GEN_7697 = opcode_3 == 4'hf ? _GEN_5647 : _GEN_7183; // @[executor.scala 466:52]
  wire [7:0] _GEN_7698 = opcode_3 == 4'hf ? _GEN_5648 : _GEN_7184; // @[executor.scala 466:52]
  wire [7:0] _GEN_7699 = opcode_3 == 4'hf ? _GEN_5649 : _GEN_7185; // @[executor.scala 466:52]
  wire [7:0] _GEN_7700 = opcode_3 == 4'hf ? _GEN_5650 : _GEN_7186; // @[executor.scala 466:52]
  wire [7:0] _GEN_7701 = opcode_3 == 4'hf ? _GEN_5651 : _GEN_7187; // @[executor.scala 466:52]
  wire [7:0] _GEN_7702 = opcode_3 == 4'hf ? _GEN_5652 : _GEN_7188; // @[executor.scala 466:52]
  wire [7:0] _GEN_7703 = opcode_3 == 4'hf ? _GEN_5653 : _GEN_7189; // @[executor.scala 466:52]
  wire [7:0] _GEN_7704 = opcode_3 == 4'hf ? _GEN_5654 : _GEN_7190; // @[executor.scala 466:52]
  wire [7:0] _GEN_7705 = opcode_3 == 4'hf ? _GEN_5655 : _GEN_7191; // @[executor.scala 466:52]
  wire [7:0] _GEN_7706 = opcode_3 == 4'hf ? _GEN_5656 : _GEN_7192; // @[executor.scala 466:52]
  wire [7:0] _GEN_7707 = opcode_3 == 4'hf ? _GEN_5657 : _GEN_7193; // @[executor.scala 466:52]
  wire [7:0] _GEN_7708 = opcode_3 == 4'hf ? _GEN_5658 : _GEN_7194; // @[executor.scala 466:52]
  wire [7:0] _GEN_7709 = opcode_3 == 4'hf ? _GEN_5659 : _GEN_7195; // @[executor.scala 466:52]
  wire [7:0] _GEN_7710 = opcode_3 == 4'hf ? _GEN_5660 : _GEN_7196; // @[executor.scala 466:52]
  wire [7:0] _GEN_7711 = opcode_3 == 4'hf ? _GEN_5661 : _GEN_7197; // @[executor.scala 466:52]
  wire [7:0] _GEN_7712 = opcode_3 == 4'hf ? _GEN_5662 : _GEN_7198; // @[executor.scala 466:52]
  wire [7:0] _GEN_7713 = opcode_3 == 4'hf ? _GEN_5663 : _GEN_7199; // @[executor.scala 466:52]
  wire [7:0] _GEN_7714 = opcode_3 == 4'hf ? _GEN_5664 : _GEN_7200; // @[executor.scala 466:52]
  wire [7:0] _GEN_7715 = opcode_3 == 4'hf ? _GEN_5665 : _GEN_7201; // @[executor.scala 466:52]
  wire [7:0] _GEN_7716 = opcode_3 == 4'hf ? _GEN_5666 : _GEN_7202; // @[executor.scala 466:52]
  wire [7:0] _GEN_7717 = opcode_3 == 4'hf ? _GEN_5667 : _GEN_7203; // @[executor.scala 466:52]
  wire [7:0] _GEN_7718 = opcode_3 == 4'hf ? _GEN_5668 : _GEN_7204; // @[executor.scala 466:52]
  wire [7:0] _GEN_7719 = opcode_3 == 4'hf ? _GEN_5669 : _GEN_7205; // @[executor.scala 466:52]
  wire [7:0] _GEN_7720 = opcode_3 == 4'hf ? _GEN_5670 : _GEN_7206; // @[executor.scala 466:52]
  wire [7:0] _GEN_7721 = opcode_3 == 4'hf ? _GEN_5671 : _GEN_7207; // @[executor.scala 466:52]
  wire [7:0] _GEN_7722 = opcode_3 == 4'hf ? _GEN_5672 : _GEN_7208; // @[executor.scala 466:52]
  wire [7:0] _GEN_7723 = opcode_3 == 4'hf ? _GEN_5673 : _GEN_7209; // @[executor.scala 466:52]
  wire [7:0] _GEN_7724 = opcode_3 == 4'hf ? _GEN_5674 : _GEN_7210; // @[executor.scala 466:52]
  wire [7:0] _GEN_7725 = opcode_3 == 4'hf ? _GEN_5675 : _GEN_7211; // @[executor.scala 466:52]
  wire [7:0] _GEN_7726 = opcode_3 == 4'hf ? _GEN_5676 : _GEN_7212; // @[executor.scala 466:52]
  wire [7:0] _GEN_7727 = opcode_3 == 4'hf ? _GEN_5677 : _GEN_7213; // @[executor.scala 466:52]
  wire [7:0] _GEN_7728 = opcode_3 == 4'hf ? _GEN_5678 : _GEN_7214; // @[executor.scala 466:52]
  wire [7:0] _GEN_7729 = opcode_3 == 4'hf ? _GEN_5679 : _GEN_7215; // @[executor.scala 466:52]
  wire [7:0] _GEN_7730 = opcode_3 == 4'hf ? _GEN_5680 : _GEN_7216; // @[executor.scala 466:52]
  wire [7:0] _GEN_7731 = opcode_3 == 4'hf ? _GEN_5681 : _GEN_7217; // @[executor.scala 466:52]
  wire [7:0] _GEN_7732 = opcode_3 == 4'hf ? _GEN_5682 : _GEN_7218; // @[executor.scala 466:52]
  wire [7:0] _GEN_7733 = opcode_3 == 4'hf ? _GEN_5683 : _GEN_7219; // @[executor.scala 466:52]
  wire [7:0] _GEN_7734 = opcode_3 == 4'hf ? _GEN_5684 : _GEN_7220; // @[executor.scala 466:52]
  wire [7:0] _GEN_7735 = opcode_3 == 4'hf ? _GEN_5685 : _GEN_7221; // @[executor.scala 466:52]
  wire [7:0] _GEN_7736 = opcode_3 == 4'hf ? _GEN_5686 : _GEN_7222; // @[executor.scala 466:52]
  wire [7:0] _GEN_7737 = opcode_3 == 4'hf ? _GEN_5687 : _GEN_7223; // @[executor.scala 466:52]
  wire [7:0] _GEN_7738 = opcode_3 == 4'hf ? _GEN_5688 : _GEN_7224; // @[executor.scala 466:52]
  wire [7:0] _GEN_7739 = opcode_3 == 4'hf ? _GEN_5689 : _GEN_7225; // @[executor.scala 466:52]
  wire [7:0] _GEN_7740 = opcode_3 == 4'hf ? _GEN_5690 : _GEN_7226; // @[executor.scala 466:52]
  wire [7:0] _GEN_7741 = opcode_3 == 4'hf ? _GEN_5691 : _GEN_7227; // @[executor.scala 466:52]
  wire [7:0] _GEN_7742 = opcode_3 == 4'hf ? _GEN_5692 : _GEN_7228; // @[executor.scala 466:52]
  wire [7:0] _GEN_7743 = opcode_3 == 4'hf ? _GEN_5693 : _GEN_7229; // @[executor.scala 466:52]
  wire [7:0] _GEN_7744 = opcode_3 == 4'hf ? _GEN_5694 : _GEN_7230; // @[executor.scala 466:52]
  wire [7:0] _GEN_7745 = opcode_3 == 4'hf ? _GEN_5695 : _GEN_7231; // @[executor.scala 466:52]
  wire [7:0] _GEN_7746 = opcode_3 == 4'hf ? _GEN_5696 : _GEN_7232; // @[executor.scala 466:52]
  wire [7:0] _GEN_7747 = opcode_3 == 4'hf ? _GEN_5697 : _GEN_7233; // @[executor.scala 466:52]
  wire [7:0] _GEN_7748 = opcode_3 == 4'hf ? _GEN_5698 : _GEN_7234; // @[executor.scala 466:52]
  wire [7:0] _GEN_7749 = opcode_3 == 4'hf ? _GEN_5699 : _GEN_7235; // @[executor.scala 466:52]
  wire [7:0] _GEN_7750 = opcode_3 == 4'hf ? _GEN_5700 : _GEN_7236; // @[executor.scala 466:52]
  wire [7:0] _GEN_7751 = opcode_3 == 4'hf ? _GEN_5701 : _GEN_7237; // @[executor.scala 466:52]
  wire [7:0] _GEN_7752 = opcode_3 == 4'hf ? _GEN_5702 : _GEN_7238; // @[executor.scala 466:52]
  wire [7:0] _GEN_7753 = opcode_3 == 4'hf ? _GEN_5703 : _GEN_7239; // @[executor.scala 466:52]
  wire [7:0] _GEN_7754 = opcode_3 == 4'hf ? _GEN_5704 : _GEN_7240; // @[executor.scala 466:52]
  wire [7:0] _GEN_7755 = opcode_3 == 4'hf ? _GEN_5705 : _GEN_7241; // @[executor.scala 466:52]
  wire [7:0] _GEN_7756 = opcode_3 == 4'hf ? _GEN_5706 : _GEN_7242; // @[executor.scala 466:52]
  wire [7:0] _GEN_7757 = opcode_3 == 4'hf ? _GEN_5707 : _GEN_7243; // @[executor.scala 466:52]
  wire [7:0] _GEN_7758 = opcode_3 == 4'hf ? _GEN_5708 : _GEN_7244; // @[executor.scala 466:52]
  wire [7:0] _GEN_7759 = opcode_3 == 4'hf ? _GEN_5709 : _GEN_7245; // @[executor.scala 466:52]
  wire [7:0] _GEN_7760 = opcode_3 == 4'hf ? _GEN_5710 : _GEN_7246; // @[executor.scala 466:52]
  wire [7:0] _GEN_7761 = opcode_3 == 4'hf ? _GEN_5711 : _GEN_7247; // @[executor.scala 466:52]
  wire [7:0] _GEN_7762 = opcode_3 == 4'hf ? _GEN_5712 : _GEN_7248; // @[executor.scala 466:52]
  wire [7:0] _GEN_7763 = opcode_3 == 4'hf ? _GEN_5713 : _GEN_7249; // @[executor.scala 466:52]
  wire [7:0] _GEN_7764 = opcode_3 == 4'hf ? _GEN_5714 : _GEN_7250; // @[executor.scala 466:52]
  wire [7:0] _GEN_7765 = opcode_3 == 4'hf ? _GEN_5715 : _GEN_7251; // @[executor.scala 466:52]
  wire [7:0] _GEN_7766 = opcode_3 == 4'hf ? _GEN_5716 : _GEN_7252; // @[executor.scala 466:52]
  wire [7:0] _GEN_7767 = opcode_3 == 4'hf ? _GEN_5717 : _GEN_7253; // @[executor.scala 466:52]
  wire [7:0] _GEN_7768 = opcode_3 == 4'hf ? _GEN_5718 : _GEN_7254; // @[executor.scala 466:52]
  wire [7:0] _GEN_7769 = opcode_3 == 4'hf ? _GEN_5719 : _GEN_7255; // @[executor.scala 466:52]
  wire [7:0] _GEN_7770 = opcode_3 == 4'hf ? _GEN_5720 : _GEN_7256; // @[executor.scala 466:52]
  wire [7:0] _GEN_7771 = opcode_3 == 4'hf ? _GEN_5721 : _GEN_7257; // @[executor.scala 466:52]
  wire [7:0] _GEN_7772 = opcode_3 == 4'hf ? _GEN_5722 : _GEN_7258; // @[executor.scala 466:52]
  wire [7:0] _GEN_7773 = opcode_3 == 4'hf ? _GEN_5723 : _GEN_7259; // @[executor.scala 466:52]
  wire [7:0] _GEN_7774 = opcode_3 == 4'hf ? _GEN_5724 : _GEN_7260; // @[executor.scala 466:52]
  wire [7:0] _GEN_7775 = opcode_3 == 4'hf ? _GEN_5725 : _GEN_7261; // @[executor.scala 466:52]
  wire [7:0] _GEN_7776 = opcode_3 == 4'hf ? _GEN_5726 : _GEN_7262; // @[executor.scala 466:52]
  wire [7:0] _GEN_7777 = opcode_3 == 4'hf ? _GEN_5727 : _GEN_7263; // @[executor.scala 466:52]
  wire [7:0] _GEN_7778 = opcode_3 == 4'hf ? _GEN_5728 : _GEN_7264; // @[executor.scala 466:52]
  wire [7:0] _GEN_7779 = opcode_3 == 4'hf ? _GEN_5729 : _GEN_7265; // @[executor.scala 466:52]
  wire [7:0] _GEN_7780 = opcode_3 == 4'hf ? _GEN_5730 : _GEN_7266; // @[executor.scala 466:52]
  wire [7:0] _GEN_7781 = opcode_3 == 4'hf ? _GEN_5731 : _GEN_7267; // @[executor.scala 466:52]
  wire [7:0] _GEN_7782 = opcode_3 == 4'hf ? _GEN_5732 : _GEN_7268; // @[executor.scala 466:52]
  wire [7:0] _GEN_7783 = opcode_3 == 4'hf ? _GEN_5733 : _GEN_7269; // @[executor.scala 466:52]
  wire [7:0] _GEN_7784 = opcode_3 == 4'hf ? _GEN_5734 : _GEN_7270; // @[executor.scala 466:52]
  wire [7:0] _GEN_7785 = opcode_3 == 4'hf ? _GEN_5735 : _GEN_7271; // @[executor.scala 466:52]
  wire [7:0] _GEN_7786 = opcode_3 == 4'hf ? _GEN_5736 : _GEN_7272; // @[executor.scala 466:52]
  wire [7:0] _GEN_7787 = opcode_3 == 4'hf ? _GEN_5737 : _GEN_7273; // @[executor.scala 466:52]
  wire [7:0] _GEN_7788 = opcode_3 == 4'hf ? _GEN_5738 : _GEN_7274; // @[executor.scala 466:52]
  wire [7:0] _GEN_7789 = opcode_3 == 4'hf ? _GEN_5739 : _GEN_7275; // @[executor.scala 466:52]
  wire [7:0] _GEN_7790 = opcode_3 == 4'hf ? _GEN_5740 : _GEN_7276; // @[executor.scala 466:52]
  wire [7:0] _GEN_7791 = opcode_3 == 4'hf ? _GEN_5741 : _GEN_7277; // @[executor.scala 466:52]
  wire [7:0] _GEN_7792 = opcode_3 == 4'hf ? _GEN_5742 : _GEN_7278; // @[executor.scala 466:52]
  wire [7:0] _GEN_7793 = opcode_3 == 4'hf ? _GEN_5743 : _GEN_7279; // @[executor.scala 466:52]
  wire [7:0] _GEN_7794 = opcode_3 == 4'hf ? _GEN_5744 : _GEN_7280; // @[executor.scala 466:52]
  wire [7:0] _GEN_7795 = opcode_3 == 4'hf ? _GEN_5745 : _GEN_7281; // @[executor.scala 466:52]
  wire [7:0] _GEN_7796 = opcode_3 == 4'hf ? _GEN_5746 : _GEN_7282; // @[executor.scala 466:52]
  wire [7:0] _GEN_7797 = opcode_3 == 4'hf ? _GEN_5747 : _GEN_7283; // @[executor.scala 466:52]
  wire [7:0] _GEN_7798 = opcode_3 == 4'hf ? _GEN_5748 : _GEN_7284; // @[executor.scala 466:52]
  wire [7:0] _GEN_7799 = opcode_3 == 4'hf ? _GEN_5749 : _GEN_7285; // @[executor.scala 466:52]
  wire [7:0] _GEN_7800 = opcode_3 == 4'hf ? _GEN_5750 : _GEN_7286; // @[executor.scala 466:52]
  wire [7:0] _GEN_7801 = opcode_3 == 4'hf ? _GEN_5751 : _GEN_7287; // @[executor.scala 466:52]
  wire [7:0] _GEN_7802 = opcode_3 == 4'hf ? _GEN_5752 : _GEN_7288; // @[executor.scala 466:52]
  wire [7:0] _GEN_7803 = opcode_3 == 4'hf ? _GEN_5753 : _GEN_7289; // @[executor.scala 466:52]
  wire [7:0] _GEN_7804 = opcode_3 == 4'hf ? _GEN_5754 : _GEN_7290; // @[executor.scala 466:52]
  wire [7:0] _GEN_7805 = opcode_3 == 4'hf ? _GEN_5755 : _GEN_7291; // @[executor.scala 466:52]
  wire [7:0] _GEN_7806 = opcode_3 == 4'hf ? _GEN_5756 : _GEN_7292; // @[executor.scala 466:52]
  wire [7:0] _GEN_7807 = opcode_3 == 4'hf ? _GEN_5757 : _GEN_7293; // @[executor.scala 466:52]
  wire [7:0] _GEN_7808 = opcode_3 == 4'hf ? _GEN_5758 : _GEN_7294; // @[executor.scala 466:52]
  wire [7:0] _GEN_7809 = opcode_3 == 4'hf ? _GEN_5759 : _GEN_7295; // @[executor.scala 466:52]
  wire [7:0] _GEN_7810 = opcode_3 == 4'hf ? _GEN_5760 : _GEN_7296; // @[executor.scala 466:52]
  wire [7:0] _GEN_7811 = opcode_3 == 4'hf ? _GEN_5761 : _GEN_7297; // @[executor.scala 466:52]
  wire [7:0] _GEN_7812 = opcode_3 == 4'hf ? _GEN_5762 : _GEN_7298; // @[executor.scala 466:52]
  wire [7:0] _GEN_7813 = opcode_3 == 4'hf ? _GEN_5763 : _GEN_7299; // @[executor.scala 466:52]
  wire [7:0] _GEN_7814 = opcode_3 == 4'hf ? _GEN_5764 : _GEN_7300; // @[executor.scala 466:52]
  wire [7:0] _GEN_7815 = opcode_3 == 4'hf ? _GEN_5765 : _GEN_7301; // @[executor.scala 466:52]
  wire [7:0] _GEN_7816 = opcode_3 == 4'hf ? _GEN_5766 : _GEN_7302; // @[executor.scala 466:52]
  wire [7:0] _GEN_7817 = opcode_3 == 4'hf ? _GEN_5767 : _GEN_7303; // @[executor.scala 466:52]
  wire [7:0] _GEN_7818 = opcode_3 == 4'hf ? _GEN_5768 : _GEN_7304; // @[executor.scala 466:52]
  wire [7:0] _GEN_7819 = opcode_3 == 4'hf ? _GEN_5769 : _GEN_7305; // @[executor.scala 466:52]
  wire [7:0] _GEN_7820 = opcode_3 == 4'hf ? _GEN_5770 : _GEN_7306; // @[executor.scala 466:52]
  wire [7:0] _GEN_7821 = opcode_3 == 4'hf ? _GEN_5771 : _GEN_7307; // @[executor.scala 466:52]
  wire [7:0] _GEN_7822 = opcode_3 == 4'hf ? _GEN_5772 : _GEN_7308; // @[executor.scala 466:52]
  wire [7:0] _GEN_7823 = opcode_3 == 4'hf ? _GEN_5773 : _GEN_7309; // @[executor.scala 466:52]
  wire [7:0] _GEN_7824 = opcode_3 == 4'hf ? _GEN_5774 : _GEN_7310; // @[executor.scala 466:52]
  wire [7:0] _GEN_7825 = opcode_3 == 4'hf ? _GEN_5775 : _GEN_7311; // @[executor.scala 466:52]
  wire [7:0] _GEN_7826 = opcode_3 == 4'hf ? _GEN_5776 : _GEN_7312; // @[executor.scala 466:52]
  wire [7:0] _GEN_7827 = opcode_3 == 4'hf ? _GEN_5777 : _GEN_7313; // @[executor.scala 466:52]
  wire [7:0] _GEN_7828 = opcode_3 == 4'hf ? _GEN_5778 : _GEN_7314; // @[executor.scala 466:52]
  wire [7:0] _GEN_7829 = opcode_3 == 4'hf ? _GEN_5779 : _GEN_7315; // @[executor.scala 466:52]
  wire [7:0] _GEN_7830 = opcode_3 == 4'hf ? _GEN_5780 : _GEN_7316; // @[executor.scala 466:52]
  wire [7:0] _GEN_7831 = opcode_3 == 4'hf ? _GEN_5781 : _GEN_7317; // @[executor.scala 466:52]
  wire [7:0] _GEN_7832 = opcode_3 == 4'hf ? _GEN_5782 : _GEN_7318; // @[executor.scala 466:52]
  wire [7:0] _GEN_7833 = opcode_3 == 4'hf ? _GEN_5783 : _GEN_7319; // @[executor.scala 466:52]
  wire [7:0] _GEN_7834 = opcode_3 == 4'hf ? _GEN_5784 : _GEN_7320; // @[executor.scala 466:52]
  wire [7:0] _GEN_7835 = opcode_3 == 4'hf ? _GEN_5785 : _GEN_7321; // @[executor.scala 466:52]
  wire [7:0] _GEN_7836 = opcode_3 == 4'hf ? _GEN_5786 : _GEN_7322; // @[executor.scala 466:52]
  wire [7:0] _GEN_7837 = opcode_3 == 4'hf ? _GEN_5787 : _GEN_7323; // @[executor.scala 466:52]
  wire [7:0] _GEN_7838 = opcode_3 == 4'hf ? _GEN_5788 : _GEN_7324; // @[executor.scala 466:52]
  wire [7:0] _GEN_7839 = opcode_3 == 4'hf ? _GEN_5789 : _GEN_7325; // @[executor.scala 466:52]
  wire [7:0] _GEN_7840 = opcode_3 == 4'hf ? _GEN_5790 : _GEN_7326; // @[executor.scala 466:52]
  wire [7:0] _GEN_7841 = opcode_3 == 4'hf ? _GEN_5791 : _GEN_7327; // @[executor.scala 466:52]
  wire [7:0] _GEN_7842 = opcode_3 == 4'hf ? _GEN_5792 : _GEN_7328; // @[executor.scala 466:52]
  wire [7:0] _GEN_7843 = opcode_3 == 4'hf ? _GEN_5793 : _GEN_7329; // @[executor.scala 466:52]
  wire [7:0] _GEN_7844 = opcode_3 == 4'hf ? _GEN_5794 : _GEN_7330; // @[executor.scala 466:52]
  wire [7:0] _GEN_7845 = opcode_3 == 4'hf ? _GEN_5795 : _GEN_7331; // @[executor.scala 466:52]
  wire [7:0] _GEN_7846 = opcode_3 == 4'hf ? _GEN_5796 : _GEN_7332; // @[executor.scala 466:52]
  wire [7:0] _GEN_7847 = opcode_3 == 4'hf ? _GEN_5797 : _GEN_7333; // @[executor.scala 466:52]
  wire [7:0] _GEN_7848 = opcode_3 == 4'hf ? _GEN_5798 : _GEN_7334; // @[executor.scala 466:52]
  wire [7:0] _GEN_7849 = opcode_3 == 4'hf ? _GEN_5799 : _GEN_7335; // @[executor.scala 466:52]
  wire [7:0] _GEN_7850 = opcode_3 == 4'hf ? _GEN_5800 : _GEN_7336; // @[executor.scala 466:52]
  wire [7:0] _GEN_7851 = opcode_3 == 4'hf ? _GEN_5801 : _GEN_7337; // @[executor.scala 466:52]
  wire [7:0] _GEN_7852 = opcode_3 == 4'hf ? _GEN_5802 : _GEN_7338; // @[executor.scala 466:52]
  wire [7:0] _GEN_7853 = opcode_3 == 4'hf ? _GEN_5803 : _GEN_7339; // @[executor.scala 466:52]
  wire [7:0] _GEN_7854 = opcode_3 == 4'hf ? _GEN_5804 : _GEN_7340; // @[executor.scala 466:52]
  wire [7:0] _GEN_7855 = opcode_3 == 4'hf ? _GEN_5805 : _GEN_7341; // @[executor.scala 466:52]
  wire [7:0] _GEN_7856 = opcode_3 == 4'hf ? _GEN_5806 : _GEN_7342; // @[executor.scala 466:52]
  wire [7:0] _GEN_7857 = opcode_3 == 4'hf ? _GEN_5807 : _GEN_7343; // @[executor.scala 466:52]
  wire [7:0] _GEN_7858 = opcode_3 == 4'hf ? _GEN_5808 : _GEN_7344; // @[executor.scala 466:52]
  wire [7:0] _GEN_7859 = opcode_3 == 4'hf ? _GEN_5809 : _GEN_7345; // @[executor.scala 466:52]
  wire [7:0] _GEN_7860 = opcode_3 == 4'hf ? _GEN_5810 : _GEN_7346; // @[executor.scala 466:52]
  wire [7:0] _GEN_7861 = opcode_3 == 4'hf ? _GEN_5811 : _GEN_7347; // @[executor.scala 466:52]
  wire [7:0] _GEN_7862 = opcode_3 == 4'hf ? _GEN_5812 : _GEN_7348; // @[executor.scala 466:52]
  wire [7:0] _GEN_7863 = opcode_3 == 4'hf ? _GEN_5813 : _GEN_7349; // @[executor.scala 466:52]
  wire [7:0] _GEN_7864 = opcode_3 == 4'hf ? _GEN_5814 : _GEN_7350; // @[executor.scala 466:52]
  wire [7:0] _GEN_7865 = opcode_3 == 4'hf ? _GEN_5815 : _GEN_7351; // @[executor.scala 466:52]
  wire [7:0] _GEN_7866 = opcode_3 == 4'hf ? _GEN_5816 : _GEN_7352; // @[executor.scala 466:52]
  wire [7:0] _GEN_7867 = opcode_3 == 4'hf ? _GEN_5817 : _GEN_7353; // @[executor.scala 466:52]
  wire [7:0] _GEN_7868 = opcode_3 == 4'hf ? _GEN_5818 : _GEN_7354; // @[executor.scala 466:52]
  wire [7:0] _GEN_7869 = opcode_3 == 4'hf ? _GEN_5819 : _GEN_7355; // @[executor.scala 466:52]
  wire [7:0] _GEN_7870 = opcode_3 == 4'hf ? _GEN_5820 : _GEN_7356; // @[executor.scala 466:52]
  wire [7:0] _GEN_7871 = opcode_3 == 4'hf ? _GEN_5821 : _GEN_7357; // @[executor.scala 466:52]
  wire [7:0] _GEN_7872 = opcode_3 == 4'hf ? _GEN_5822 : _GEN_7358; // @[executor.scala 466:52]
  wire [7:0] _GEN_7873 = opcode_3 == 4'hf ? _GEN_5823 : _GEN_7359; // @[executor.scala 466:52]
  wire [7:0] _GEN_7874 = opcode_3 == 4'hf ? _GEN_5824 : _GEN_7360; // @[executor.scala 466:52]
  wire [7:0] _GEN_7875 = opcode_3 == 4'hf ? _GEN_5825 : _GEN_7361; // @[executor.scala 466:52]
  wire [7:0] _GEN_7876 = opcode_3 == 4'hf ? _GEN_5826 : _GEN_7362; // @[executor.scala 466:52]
  wire [7:0] _GEN_7877 = opcode_3 == 4'hf ? _GEN_5827 : _GEN_7363; // @[executor.scala 466:52]
  wire [7:0] _GEN_7878 = opcode_3 == 4'hf ? _GEN_5828 : _GEN_7364; // @[executor.scala 466:52]
  wire [7:0] _GEN_7879 = opcode_3 == 4'hf ? _GEN_5829 : _GEN_7365; // @[executor.scala 466:52]
  wire [7:0] _GEN_7880 = opcode_3 == 4'hf ? _GEN_5830 : _GEN_7366; // @[executor.scala 466:52]
  wire [7:0] _GEN_7881 = opcode_3 == 4'hf ? _GEN_5831 : _GEN_7367; // @[executor.scala 466:52]
  wire [7:0] _GEN_7882 = opcode_3 == 4'hf ? _GEN_5832 : _GEN_7368; // @[executor.scala 466:52]
  wire [7:0] _GEN_7883 = opcode_3 == 4'hf ? _GEN_5833 : _GEN_7369; // @[executor.scala 466:52]
  wire [7:0] _GEN_7884 = opcode_3 == 4'hf ? _GEN_5834 : _GEN_7370; // @[executor.scala 466:52]
  wire [7:0] _GEN_7885 = opcode_3 == 4'hf ? _GEN_5835 : _GEN_7371; // @[executor.scala 466:52]
  wire [7:0] _GEN_7886 = opcode_3 == 4'hf ? _GEN_5836 : _GEN_7372; // @[executor.scala 466:52]
  wire [7:0] _GEN_7887 = opcode_3 == 4'hf ? _GEN_5837 : _GEN_7373; // @[executor.scala 466:52]
  wire [7:0] _GEN_7888 = opcode_3 == 4'hf ? _GEN_5838 : _GEN_7374; // @[executor.scala 466:52]
  wire [7:0] _GEN_7889 = opcode_3 == 4'hf ? _GEN_5839 : _GEN_7375; // @[executor.scala 466:52]
  wire [7:0] _GEN_7890 = opcode_3 == 4'hf ? _GEN_5840 : _GEN_7376; // @[executor.scala 466:52]
  wire [7:0] _GEN_7891 = opcode_3 == 4'hf ? _GEN_5841 : _GEN_7377; // @[executor.scala 466:52]
  wire [7:0] _GEN_7892 = opcode_3 == 4'hf ? _GEN_5842 : _GEN_7378; // @[executor.scala 466:52]
  wire [7:0] _GEN_7893 = opcode_3 == 4'hf ? _GEN_5843 : _GEN_7379; // @[executor.scala 466:52]
  wire [7:0] _GEN_7894 = opcode_3 == 4'hf ? _GEN_5844 : _GEN_7380; // @[executor.scala 466:52]
  wire [7:0] _GEN_7895 = opcode_3 == 4'hf ? _GEN_5845 : _GEN_7381; // @[executor.scala 466:52]
  wire [7:0] _GEN_7896 = opcode_3 == 4'hf ? _GEN_5846 : _GEN_7382; // @[executor.scala 466:52]
  wire [7:0] _GEN_7897 = opcode_3 == 4'hf ? _GEN_5847 : _GEN_7383; // @[executor.scala 466:52]
  wire [7:0] _GEN_7898 = opcode_3 == 4'hf ? _GEN_5848 : _GEN_7384; // @[executor.scala 466:52]
  wire [7:0] _GEN_7899 = opcode_3 == 4'hf ? _GEN_5849 : _GEN_7385; // @[executor.scala 466:52]
  wire [7:0] _GEN_7900 = opcode_3 == 4'hf ? _GEN_5850 : _GEN_7386; // @[executor.scala 466:52]
  wire [7:0] _GEN_7901 = opcode_3 == 4'hf ? _GEN_5851 : _GEN_7387; // @[executor.scala 466:52]
  wire [7:0] _GEN_7902 = opcode_3 == 4'hf ? _GEN_5852 : _GEN_7388; // @[executor.scala 466:52]
  wire [7:0] _GEN_7903 = opcode_3 == 4'hf ? _GEN_5853 : _GEN_7389; // @[executor.scala 466:52]
  wire [7:0] _GEN_7904 = opcode_3 == 4'hf ? _GEN_5854 : _GEN_7390; // @[executor.scala 466:52]
  wire [7:0] _GEN_7905 = opcode_3 == 4'hf ? _GEN_5855 : _GEN_7391; // @[executor.scala 466:52]
  wire [7:0] _GEN_7906 = opcode_3 == 4'hf ? _GEN_5856 : _GEN_7392; // @[executor.scala 466:52]
  wire [7:0] _GEN_7907 = opcode_3 == 4'hf ? _GEN_5857 : _GEN_7393; // @[executor.scala 466:52]
  wire [7:0] _GEN_7908 = opcode_3 == 4'hf ? _GEN_5858 : _GEN_7394; // @[executor.scala 466:52]
  wire [7:0] _GEN_7909 = opcode_3 == 4'hf ? _GEN_5859 : _GEN_7395; // @[executor.scala 466:52]
  wire [7:0] _GEN_7910 = opcode_3 == 4'hf ? _GEN_5860 : _GEN_7396; // @[executor.scala 466:52]
  wire [7:0] _GEN_7911 = opcode_3 == 4'hf ? _GEN_5861 : _GEN_7397; // @[executor.scala 466:52]
  wire [7:0] _GEN_7912 = opcode_3 == 4'hf ? _GEN_5862 : _GEN_7398; // @[executor.scala 466:52]
  wire [7:0] _GEN_7913 = opcode_3 == 4'hf ? _GEN_5863 : _GEN_7399; // @[executor.scala 466:52]
  wire [7:0] _GEN_7914 = opcode_3 == 4'hf ? _GEN_5864 : _GEN_7400; // @[executor.scala 466:52]
  wire [7:0] _GEN_7915 = opcode_3 == 4'hf ? _GEN_5865 : _GEN_7401; // @[executor.scala 466:52]
  wire [7:0] _GEN_7916 = opcode_3 == 4'hf ? _GEN_5866 : _GEN_7402; // @[executor.scala 466:52]
  wire [7:0] _GEN_7917 = opcode_3 == 4'hf ? _GEN_5867 : _GEN_7403; // @[executor.scala 466:52]
  wire [7:0] _GEN_7918 = opcode_3 == 4'hf ? _GEN_5868 : _GEN_7404; // @[executor.scala 466:52]
  wire [7:0] _GEN_7919 = opcode_3 == 4'hf ? _GEN_5869 : _GEN_7405; // @[executor.scala 466:52]
  wire [7:0] _GEN_7920 = opcode_3 == 4'hf ? _GEN_5870 : _GEN_7406; // @[executor.scala 466:52]
  wire [7:0] _GEN_7921 = opcode_3 == 4'hf ? _GEN_5871 : _GEN_7407; // @[executor.scala 466:52]
  wire [7:0] _GEN_7922 = opcode_3 == 4'hf ? _GEN_5872 : _GEN_7408; // @[executor.scala 466:52]
  wire [7:0] _GEN_7923 = opcode_3 == 4'hf ? _GEN_5873 : _GEN_7409; // @[executor.scala 466:52]
  wire [7:0] _GEN_7924 = opcode_3 == 4'hf ? _GEN_5874 : _GEN_7410; // @[executor.scala 466:52]
  wire [7:0] _GEN_7925 = opcode_3 == 4'hf ? _GEN_5875 : _GEN_7411; // @[executor.scala 466:52]
  wire [7:0] _GEN_7926 = opcode_3 == 4'hf ? _GEN_5876 : _GEN_7412; // @[executor.scala 466:52]
  wire [7:0] _GEN_7927 = opcode_3 == 4'hf ? _GEN_5877 : _GEN_7413; // @[executor.scala 466:52]
  wire [7:0] _GEN_7928 = opcode_3 == 4'hf ? _GEN_5878 : _GEN_7414; // @[executor.scala 466:52]
  wire [7:0] _GEN_7929 = opcode_3 == 4'hf ? _GEN_5879 : _GEN_7415; // @[executor.scala 466:52]
  wire [7:0] _GEN_7930 = opcode_3 == 4'hf ? _GEN_5880 : _GEN_7416; // @[executor.scala 466:52]
  wire [7:0] _GEN_7931 = opcode_3 == 4'hf ? _GEN_5881 : _GEN_7417; // @[executor.scala 466:52]
  wire [7:0] _GEN_7932 = opcode_3 == 4'hf ? _GEN_5882 : _GEN_7418; // @[executor.scala 466:52]
  wire [7:0] _GEN_7933 = opcode_3 == 4'hf ? _GEN_5883 : _GEN_7419; // @[executor.scala 466:52]
  wire [7:0] _GEN_7934 = opcode_3 == 4'hf ? _GEN_5884 : _GEN_7420; // @[executor.scala 466:52]
  wire [7:0] _GEN_7935 = opcode_3 == 4'hf ? _GEN_5885 : _GEN_7421; // @[executor.scala 466:52]
  wire [7:0] _GEN_7936 = opcode_3 == 4'hf ? _GEN_5886 : _GEN_7422; // @[executor.scala 466:52]
  wire [7:0] _GEN_7937 = opcode_3 == 4'hf ? _GEN_5887 : _GEN_7423; // @[executor.scala 466:52]
  wire [7:0] _GEN_7938 = opcode_3 == 4'hf ? _GEN_5888 : _GEN_7424; // @[executor.scala 466:52]
  wire [7:0] _GEN_7939 = opcode_3 == 4'hf ? _GEN_5889 : _GEN_7425; // @[executor.scala 466:52]
  wire [7:0] _GEN_7940 = opcode_3 == 4'hf ? _GEN_5890 : _GEN_7426; // @[executor.scala 466:52]
  wire [7:0] _GEN_7941 = opcode_3 == 4'hf ? _GEN_5891 : _GEN_7427; // @[executor.scala 466:52]
  wire [7:0] _GEN_7942 = opcode_3 == 4'hf ? _GEN_5892 : _GEN_7428; // @[executor.scala 466:52]
  wire [7:0] _GEN_7943 = opcode_3 == 4'hf ? _GEN_5893 : _GEN_7429; // @[executor.scala 466:52]
  wire [7:0] _GEN_7944 = opcode_3 == 4'hf ? _GEN_5894 : _GEN_7430; // @[executor.scala 466:52]
  wire [7:0] _GEN_7945 = opcode_3 == 4'hf ? _GEN_5895 : _GEN_7431; // @[executor.scala 466:52]
  wire [7:0] _GEN_7946 = opcode_3 == 4'hf ? _GEN_5896 : _GEN_7432; // @[executor.scala 466:52]
  wire [7:0] _GEN_7947 = opcode_3 == 4'hf ? _GEN_5897 : _GEN_7433; // @[executor.scala 466:52]
  wire [7:0] _GEN_7948 = opcode_3 == 4'hf ? _GEN_5898 : _GEN_7434; // @[executor.scala 466:52]
  wire [7:0] _GEN_7949 = opcode_3 == 4'hf ? _GEN_5899 : _GEN_7435; // @[executor.scala 466:52]
  wire [7:0] _GEN_7950 = opcode_3 == 4'hf ? _GEN_5900 : _GEN_7436; // @[executor.scala 466:52]
  wire [7:0] _GEN_7951 = opcode_3 == 4'hf ? _GEN_5901 : _GEN_7437; // @[executor.scala 466:52]
  wire [7:0] _GEN_7952 = opcode_3 == 4'hf ? _GEN_5902 : _GEN_7438; // @[executor.scala 466:52]
  wire [7:0] _GEN_7953 = opcode_3 == 4'hf ? _GEN_5903 : _GEN_7439; // @[executor.scala 466:52]
  wire [7:0] _GEN_7954 = opcode_3 == 4'hf ? _GEN_5904 : _GEN_7440; // @[executor.scala 466:52]
  wire [7:0] _GEN_7955 = opcode_3 == 4'hf ? _GEN_5905 : _GEN_7441; // @[executor.scala 466:52]
  wire [7:0] _GEN_7956 = opcode_3 == 4'hf ? _GEN_5906 : _GEN_7442; // @[executor.scala 466:52]
  wire [7:0] _GEN_7957 = opcode_3 == 4'hf ? _GEN_5907 : _GEN_7443; // @[executor.scala 466:52]
  wire [7:0] _GEN_7958 = opcode_3 == 4'hf ? _GEN_5908 : _GEN_7444; // @[executor.scala 466:52]
  wire [7:0] _GEN_7959 = opcode_3 == 4'hf ? _GEN_5909 : _GEN_7445; // @[executor.scala 466:52]
  wire [7:0] _GEN_7960 = opcode_3 == 4'hf ? _GEN_5910 : _GEN_7446; // @[executor.scala 466:52]
  wire [7:0] _GEN_7961 = opcode_3 == 4'hf ? _GEN_5911 : _GEN_7447; // @[executor.scala 466:52]
  wire [7:0] _GEN_7962 = opcode_3 == 4'hf ? _GEN_5912 : _GEN_7448; // @[executor.scala 466:52]
  wire [7:0] _GEN_7963 = opcode_3 == 4'hf ? _GEN_5913 : _GEN_7449; // @[executor.scala 466:52]
  wire [7:0] _GEN_7964 = opcode_3 == 4'hf ? _GEN_5914 : _GEN_7450; // @[executor.scala 466:52]
  wire [7:0] _GEN_7965 = opcode_3 == 4'hf ? _GEN_5915 : _GEN_7451; // @[executor.scala 466:52]
  wire [7:0] _GEN_7966 = opcode_3 == 4'hf ? _GEN_5916 : _GEN_7452; // @[executor.scala 466:52]
  wire [7:0] _GEN_7967 = opcode_3 == 4'hf ? _GEN_5917 : _GEN_7453; // @[executor.scala 466:52]
  wire [7:0] _GEN_7968 = opcode_3 == 4'hf ? _GEN_5918 : _GEN_7454; // @[executor.scala 466:52]
  wire [7:0] _GEN_7969 = opcode_3 == 4'hf ? _GEN_5919 : _GEN_7455; // @[executor.scala 466:52]
  wire [7:0] _GEN_7970 = opcode_3 == 4'hf ? _GEN_5920 : _GEN_7456; // @[executor.scala 466:52]
  wire [7:0] _GEN_7971 = opcode_3 == 4'hf ? _GEN_5921 : _GEN_7457; // @[executor.scala 466:52]
  wire [7:0] _GEN_7972 = opcode_3 == 4'hf ? _GEN_5922 : _GEN_7458; // @[executor.scala 466:52]
  wire [7:0] _GEN_7973 = opcode_3 == 4'hf ? _GEN_5923 : _GEN_7459; // @[executor.scala 466:52]
  wire [7:0] _GEN_7974 = opcode_3 == 4'hf ? _GEN_5924 : _GEN_7460; // @[executor.scala 466:52]
  wire [7:0] _GEN_7975 = opcode_3 == 4'hf ? _GEN_5925 : _GEN_7461; // @[executor.scala 466:52]
  wire [7:0] _GEN_7976 = opcode_3 == 4'hf ? _GEN_5926 : _GEN_7462; // @[executor.scala 466:52]
  wire [7:0] _GEN_7977 = opcode_3 == 4'hf ? _GEN_5927 : _GEN_7463; // @[executor.scala 466:52]
  wire [7:0] _GEN_7978 = opcode_3 == 4'hf ? _GEN_5928 : _GEN_7464; // @[executor.scala 466:52]
  wire [7:0] _GEN_7979 = opcode_3 == 4'hf ? _GEN_5929 : _GEN_7465; // @[executor.scala 466:52]
  wire [7:0] _GEN_7980 = opcode_3 == 4'hf ? _GEN_5930 : _GEN_7466; // @[executor.scala 466:52]
  wire [7:0] _GEN_7981 = opcode_3 == 4'hf ? _GEN_5931 : _GEN_7467; // @[executor.scala 466:52]
  wire [7:0] _GEN_7982 = opcode_3 == 4'hf ? _GEN_5932 : _GEN_7468; // @[executor.scala 466:52]
  wire [7:0] _GEN_7983 = opcode_3 == 4'hf ? _GEN_5933 : _GEN_7469; // @[executor.scala 466:52]
  wire [7:0] _GEN_7984 = opcode_3 == 4'hf ? _GEN_5934 : _GEN_7470; // @[executor.scala 466:52]
  wire [7:0] _GEN_7985 = opcode_3 == 4'hf ? _GEN_5935 : _GEN_7471; // @[executor.scala 466:52]
  wire [7:0] _GEN_7986 = opcode_3 == 4'hf ? _GEN_5936 : _GEN_7472; // @[executor.scala 466:52]
  wire [7:0] _GEN_7987 = opcode_3 == 4'hf ? _GEN_5937 : _GEN_7473; // @[executor.scala 466:52]
  wire [7:0] _GEN_7988 = opcode_3 == 4'hf ? _GEN_5938 : _GEN_7474; // @[executor.scala 466:52]
  wire [7:0] _GEN_7989 = opcode_3 == 4'hf ? _GEN_5939 : _GEN_7475; // @[executor.scala 466:52]
  wire [7:0] _GEN_7990 = opcode_3 == 4'hf ? _GEN_5940 : _GEN_7476; // @[executor.scala 466:52]
  wire [7:0] _GEN_7991 = opcode_3 == 4'hf ? _GEN_5941 : _GEN_7477; // @[executor.scala 466:52]
  wire [7:0] _GEN_7992 = opcode_3 == 4'hf ? _GEN_5942 : _GEN_7478; // @[executor.scala 466:52]
  wire [7:0] _GEN_7993 = opcode_3 == 4'hf ? _GEN_5943 : _GEN_7479; // @[executor.scala 466:52]
  wire [7:0] _GEN_7994 = opcode_3 == 4'hf ? _GEN_5944 : _GEN_7480; // @[executor.scala 466:52]
  wire [7:0] _GEN_7995 = opcode_3 == 4'hf ? _GEN_5945 : _GEN_7481; // @[executor.scala 466:52]
  wire [7:0] _GEN_7996 = opcode_3 == 4'hf ? _GEN_5946 : _GEN_7482; // @[executor.scala 466:52]
  wire [7:0] _GEN_7997 = opcode_3 == 4'hf ? _GEN_5947 : _GEN_7483; // @[executor.scala 466:52]
  wire [7:0] _GEN_7998 = opcode_3 == 4'hf ? _GEN_5948 : _GEN_7484; // @[executor.scala 466:52]
  wire [7:0] _GEN_7999 = opcode_3 == 4'hf ? _GEN_5949 : _GEN_7485; // @[executor.scala 466:52]
  wire [7:0] _GEN_8000 = opcode_3 == 4'hf ? _GEN_5950 : _GEN_7486; // @[executor.scala 466:52]
  wire [7:0] _GEN_8001 = opcode_3 == 4'hf ? _GEN_5951 : _GEN_7487; // @[executor.scala 466:52]
  wire [7:0] _GEN_8002 = opcode_3 == 4'hf ? _GEN_5952 : _GEN_7488; // @[executor.scala 466:52]
  wire [7:0] _GEN_8003 = opcode_3 == 4'hf ? _GEN_5953 : _GEN_7489; // @[executor.scala 466:52]
  wire [7:0] _GEN_8004 = opcode_3 == 4'hf ? _GEN_5954 : _GEN_7490; // @[executor.scala 466:52]
  wire [7:0] _GEN_8005 = opcode_3 == 4'hf ? _GEN_5955 : _GEN_7491; // @[executor.scala 466:52]
  wire [7:0] _GEN_8006 = opcode_3 == 4'hf ? _GEN_5956 : _GEN_7492; // @[executor.scala 466:52]
  wire [7:0] _GEN_8007 = opcode_3 == 4'hf ? _GEN_5957 : _GEN_7493; // @[executor.scala 466:52]
  wire [7:0] _GEN_8008 = opcode_3 == 4'hf ? _GEN_5958 : _GEN_7494; // @[executor.scala 466:52]
  wire [7:0] _GEN_8009 = opcode_3 == 4'hf ? _GEN_5959 : _GEN_7495; // @[executor.scala 466:52]
  wire [7:0] _GEN_8010 = opcode_3 == 4'hf ? _GEN_5960 : _GEN_7496; // @[executor.scala 466:52]
  wire [7:0] _GEN_8011 = opcode_3 == 4'hf ? _GEN_5961 : _GEN_7497; // @[executor.scala 466:52]
  wire [7:0] _GEN_8012 = opcode_3 == 4'hf ? _GEN_5962 : _GEN_7498; // @[executor.scala 466:52]
  wire [7:0] _GEN_8013 = opcode_3 == 4'hf ? _GEN_5963 : _GEN_7499; // @[executor.scala 466:52]
  wire [7:0] _GEN_8014 = opcode_3 == 4'hf ? _GEN_5964 : _GEN_7500; // @[executor.scala 466:52]
  wire [7:0] _GEN_8015 = opcode_3 == 4'hf ? _GEN_5965 : _GEN_7501; // @[executor.scala 466:52]
  wire [7:0] _GEN_8016 = opcode_3 == 4'hf ? _GEN_5966 : _GEN_7502; // @[executor.scala 466:52]
  wire [7:0] _GEN_8017 = opcode_3 == 4'hf ? _GEN_5967 : _GEN_7503; // @[executor.scala 466:52]
  wire [7:0] _GEN_8018 = opcode_3 == 4'hf ? _GEN_5968 : _GEN_7504; // @[executor.scala 466:52]
  wire [7:0] _GEN_8019 = opcode_3 == 4'hf ? _GEN_5969 : _GEN_7505; // @[executor.scala 466:52]
  wire [7:0] _GEN_8020 = opcode_3 == 4'hf ? _GEN_5970 : _GEN_7506; // @[executor.scala 466:52]
  wire [7:0] _GEN_8021 = opcode_3 == 4'hf ? _GEN_5971 : _GEN_7507; // @[executor.scala 466:52]
  wire [7:0] _GEN_8022 = opcode_3 == 4'hf ? _GEN_5972 : _GEN_7508; // @[executor.scala 466:52]
  wire [7:0] _GEN_8023 = opcode_3 == 4'hf ? _GEN_5973 : _GEN_7509; // @[executor.scala 466:52]
  wire [7:0] _GEN_8024 = opcode_3 == 4'hf ? _GEN_5974 : _GEN_7510; // @[executor.scala 466:52]
  wire [7:0] _GEN_8025 = opcode_3 == 4'hf ? _GEN_5975 : _GEN_7511; // @[executor.scala 466:52]
  wire [7:0] _GEN_8026 = opcode_3 == 4'hf ? _GEN_5976 : _GEN_7512; // @[executor.scala 466:52]
  wire [7:0] _GEN_8027 = opcode_3 == 4'hf ? _GEN_5977 : _GEN_7513; // @[executor.scala 466:52]
  wire [7:0] _GEN_8028 = opcode_3 == 4'hf ? _GEN_5978 : _GEN_7514; // @[executor.scala 466:52]
  wire [7:0] _GEN_8029 = opcode_3 == 4'hf ? _GEN_5979 : _GEN_7515; // @[executor.scala 466:52]
  wire [7:0] _GEN_8030 = opcode_3 == 4'hf ? _GEN_5980 : _GEN_7516; // @[executor.scala 466:52]
  wire [7:0] _GEN_8031 = opcode_3 == 4'hf ? _GEN_5981 : _GEN_7517; // @[executor.scala 466:52]
  wire [7:0] _GEN_8032 = opcode_3 == 4'hf ? _GEN_5982 : _GEN_7518; // @[executor.scala 466:52]
  wire [7:0] _GEN_8033 = opcode_3 == 4'hf ? _GEN_5983 : _GEN_7519; // @[executor.scala 466:52]
  wire [7:0] _GEN_8034 = opcode_3 == 4'hf ? _GEN_5984 : _GEN_7520; // @[executor.scala 466:52]
  wire [7:0] _GEN_8035 = opcode_3 == 4'hf ? _GEN_5985 : _GEN_7521; // @[executor.scala 466:52]
  wire [7:0] _GEN_8036 = opcode_3 == 4'hf ? _GEN_5986 : _GEN_7522; // @[executor.scala 466:52]
  wire [7:0] _GEN_8037 = opcode_3 == 4'hf ? _GEN_5987 : _GEN_7523; // @[executor.scala 466:52]
  wire [7:0] _GEN_8038 = opcode_3 == 4'hf ? _GEN_5988 : _GEN_7524; // @[executor.scala 466:52]
  wire [7:0] _GEN_8039 = opcode_3 == 4'hf ? _GEN_5989 : _GEN_7525; // @[executor.scala 466:52]
  wire [7:0] _GEN_8040 = opcode_3 == 4'hf ? _GEN_5990 : _GEN_7526; // @[executor.scala 466:52]
  wire [7:0] _GEN_8041 = opcode_3 == 4'hf ? _GEN_5991 : _GEN_7527; // @[executor.scala 466:52]
  wire [7:0] _GEN_8042 = opcode_3 == 4'hf ? _GEN_5992 : _GEN_7528; // @[executor.scala 466:52]
  wire [7:0] _GEN_8043 = opcode_3 == 4'hf ? _GEN_5993 : _GEN_7529; // @[executor.scala 466:52]
  wire [7:0] _GEN_8044 = opcode_3 == 4'hf ? _GEN_5994 : _GEN_7530; // @[executor.scala 466:52]
  wire [7:0] _GEN_8045 = opcode_3 == 4'hf ? _GEN_5995 : _GEN_7531; // @[executor.scala 466:52]
  wire [7:0] _GEN_8046 = opcode_3 == 4'hf ? _GEN_5996 : _GEN_7532; // @[executor.scala 466:52]
  wire [7:0] _GEN_8047 = opcode_3 == 4'hf ? _GEN_5997 : _GEN_7533; // @[executor.scala 466:52]
  wire [7:0] _GEN_8048 = opcode_3 == 4'hf ? _GEN_5998 : _GEN_7534; // @[executor.scala 466:52]
  wire [7:0] _GEN_8049 = opcode_3 == 4'hf ? _GEN_5999 : _GEN_7535; // @[executor.scala 466:52]
  wire [7:0] _GEN_8050 = opcode_3 == 4'hf ? _GEN_6000 : _GEN_7536; // @[executor.scala 466:52]
  wire [7:0] _GEN_8051 = opcode_3 == 4'hf ? _GEN_6001 : _GEN_7537; // @[executor.scala 466:52]
  wire [7:0] _GEN_8052 = opcode_3 == 4'hf ? _GEN_6002 : _GEN_7538; // @[executor.scala 466:52]
  wire [7:0] _GEN_8053 = opcode_3 == 4'hf ? _GEN_6003 : _GEN_7539; // @[executor.scala 466:52]
  wire [7:0] _GEN_8054 = opcode_3 == 4'hf ? _GEN_6004 : _GEN_7540; // @[executor.scala 466:52]
  wire [7:0] _GEN_8055 = opcode_3 == 4'hf ? _GEN_6005 : _GEN_7541; // @[executor.scala 466:52]
  wire [7:0] _GEN_8056 = opcode_3 == 4'hf ? _GEN_6006 : _GEN_7542; // @[executor.scala 466:52]
  wire [7:0] _GEN_8057 = opcode_3 == 4'hf ? _GEN_6007 : _GEN_7543; // @[executor.scala 466:52]
  wire [7:0] _GEN_8058 = opcode_3 == 4'hf ? _GEN_6008 : _GEN_7544; // @[executor.scala 466:52]
  wire [7:0] _GEN_8059 = opcode_3 == 4'hf ? _GEN_6009 : _GEN_7545; // @[executor.scala 466:52]
  wire [7:0] _GEN_8060 = opcode_3 == 4'hf ? _GEN_6010 : _GEN_7546; // @[executor.scala 466:52]
  wire [7:0] _GEN_8061 = opcode_3 == 4'hf ? _GEN_6011 : _GEN_7547; // @[executor.scala 466:52]
  wire [7:0] _GEN_8062 = opcode_3 == 4'hf ? _GEN_6012 : _GEN_7548; // @[executor.scala 466:52]
  wire [7:0] _GEN_8063 = opcode_3 == 4'hf ? _GEN_6013 : _GEN_7549; // @[executor.scala 466:52]
  wire [7:0] _GEN_8064 = opcode_3 == 4'hf ? _GEN_6014 : _GEN_7550; // @[executor.scala 466:52]
  wire [7:0] _GEN_8065 = opcode_3 == 4'hf ? _GEN_6015 : _GEN_7551; // @[executor.scala 466:52]
  wire [7:0] _GEN_8066 = opcode_3 == 4'hf ? _GEN_6016 : _GEN_7552; // @[executor.scala 466:52]
  wire [7:0] _GEN_8067 = opcode_3 == 4'hf ? _GEN_6017 : _GEN_7553; // @[executor.scala 466:52]
  wire [7:0] _GEN_8068 = opcode_3 == 4'hf ? _GEN_6018 : _GEN_7554; // @[executor.scala 466:52]
  wire [7:0] _GEN_8069 = opcode_3 == 4'hf ? _GEN_6019 : _GEN_7555; // @[executor.scala 466:52]
  wire [7:0] _GEN_8070 = opcode_3 == 4'hf ? _GEN_6020 : _GEN_7556; // @[executor.scala 466:52]
  wire [7:0] _GEN_8071 = opcode_3 == 4'hf ? _GEN_6021 : _GEN_7557; // @[executor.scala 466:52]
  wire [7:0] _GEN_8072 = opcode_3 == 4'hf ? _GEN_6022 : _GEN_7558; // @[executor.scala 466:52]
  wire [7:0] _GEN_8073 = opcode_3 == 4'hf ? _GEN_6023 : _GEN_7559; // @[executor.scala 466:52]
  wire [7:0] _GEN_8074 = opcode_3 == 4'hf ? _GEN_6024 : _GEN_7560; // @[executor.scala 466:52]
  wire [7:0] _GEN_8075 = opcode_3 == 4'hf ? _GEN_6025 : _GEN_7561; // @[executor.scala 466:52]
  wire [7:0] _GEN_8076 = opcode_3 == 4'hf ? _GEN_6026 : _GEN_7562; // @[executor.scala 466:52]
  wire [7:0] _GEN_8077 = opcode_3 == 4'hf ? _GEN_6027 : _GEN_7563; // @[executor.scala 466:52]
  wire [7:0] _GEN_8078 = opcode_3 == 4'hf ? _GEN_6028 : _GEN_7564; // @[executor.scala 466:52]
  wire [7:0] _GEN_8079 = opcode_3 == 4'hf ? _GEN_6029 : _GEN_7565; // @[executor.scala 466:52]
  wire [7:0] _GEN_8080 = opcode_3 == 4'hf ? _GEN_6030 : _GEN_7566; // @[executor.scala 466:52]
  wire [7:0] _GEN_8081 = opcode_3 == 4'hf ? _GEN_6031 : _GEN_7567; // @[executor.scala 466:52]
  wire [7:0] _GEN_8082 = opcode_3 == 4'hf ? _GEN_6032 : _GEN_7568; // @[executor.scala 466:52]
  wire [7:0] _GEN_8083 = opcode_3 == 4'hf ? _GEN_6033 : _GEN_7569; // @[executor.scala 466:52]
  wire [7:0] _GEN_8084 = opcode_3 == 4'hf ? _GEN_6034 : _GEN_7570; // @[executor.scala 466:52]
  wire [7:0] _GEN_8085 = opcode_3 == 4'hf ? _GEN_6035 : _GEN_7571; // @[executor.scala 466:52]
  wire [7:0] _GEN_8086 = opcode_3 == 4'hf ? _GEN_6036 : _GEN_7572; // @[executor.scala 466:52]
  wire [7:0] _GEN_8087 = opcode_3 == 4'hf ? _GEN_6037 : _GEN_7573; // @[executor.scala 466:52]
  wire [7:0] _GEN_8088 = opcode_3 == 4'hf ? _GEN_6038 : _GEN_7574; // @[executor.scala 466:52]
  wire [7:0] _GEN_8089 = opcode_3 == 4'hf ? _GEN_6039 : _GEN_7575; // @[executor.scala 466:52]
  wire [7:0] _GEN_8090 = opcode_3 == 4'hf ? _GEN_6040 : _GEN_7576; // @[executor.scala 466:52]
  wire [7:0] _GEN_8091 = opcode_3 == 4'hf ? _GEN_6041 : _GEN_7577; // @[executor.scala 466:52]
  wire [7:0] _GEN_8092 = opcode_3 == 4'hf ? _GEN_6042 : _GEN_7578; // @[executor.scala 466:52]
  wire [7:0] _GEN_8093 = opcode_3 == 4'hf ? _GEN_6043 : _GEN_7579; // @[executor.scala 466:52]
  wire [7:0] _GEN_8094 = opcode_3 == 4'hf ? _GEN_6044 : _GEN_7580; // @[executor.scala 466:52]
  wire [7:0] _GEN_8095 = opcode_3 == 4'hf ? _GEN_6045 : _GEN_7581; // @[executor.scala 466:52]
  wire [7:0] _GEN_8096 = opcode_3 == 4'hf ? _GEN_6046 : _GEN_7582; // @[executor.scala 466:52]
  wire [7:0] _GEN_8097 = opcode_3 == 4'hf ? _GEN_6047 : _GEN_7583; // @[executor.scala 466:52]
  wire [7:0] _GEN_8098 = opcode_3 == 4'hf ? _GEN_6048 : _GEN_7584; // @[executor.scala 466:52]
  wire [7:0] _GEN_8099 = opcode_3 == 4'hf ? _GEN_6049 : _GEN_7585; // @[executor.scala 466:52]
  wire [7:0] _GEN_8100 = opcode_3 == 4'hf ? _GEN_6050 : _GEN_7586; // @[executor.scala 466:52]
  wire [7:0] _GEN_8101 = opcode_3 == 4'hf ? _GEN_6051 : _GEN_7587; // @[executor.scala 466:52]
  wire [7:0] _GEN_8102 = opcode_3 == 4'hf ? _GEN_6052 : _GEN_7588; // @[executor.scala 466:52]
  wire [7:0] _GEN_8103 = opcode_3 == 4'hf ? _GEN_6053 : _GEN_7589; // @[executor.scala 466:52]
  wire [7:0] _GEN_8104 = opcode_3 == 4'hf ? _GEN_6054 : _GEN_7590; // @[executor.scala 466:52]
  wire [7:0] _GEN_8105 = opcode_3 == 4'hf ? _GEN_6055 : _GEN_7591; // @[executor.scala 466:52]
  wire [7:0] _GEN_8106 = opcode_3 == 4'hf ? _GEN_6056 : _GEN_7592; // @[executor.scala 466:52]
  wire [7:0] _GEN_8107 = opcode_3 == 4'hf ? _GEN_6057 : _GEN_7593; // @[executor.scala 466:52]
  wire [7:0] _GEN_8108 = opcode_3 == 4'hf ? _GEN_6058 : _GEN_7594; // @[executor.scala 466:52]
  wire [7:0] _GEN_8109 = opcode_3 == 4'hf ? _GEN_6059 : _GEN_7595; // @[executor.scala 466:52]
  wire [7:0] _GEN_8110 = opcode_3 == 4'hf ? _GEN_6060 : _GEN_7596; // @[executor.scala 466:52]
  wire [7:0] _GEN_8111 = opcode_3 == 4'hf ? _GEN_6061 : _GEN_7597; // @[executor.scala 466:52]
  wire [7:0] _GEN_8112 = opcode_3 == 4'hf ? _GEN_6062 : _GEN_7598; // @[executor.scala 466:52]
  wire [7:0] _GEN_8113 = opcode_3 == 4'hf ? _GEN_6063 : _GEN_7599; // @[executor.scala 466:52]
  wire [7:0] _GEN_8114 = opcode_3 == 4'hf ? _GEN_6064 : _GEN_7600; // @[executor.scala 466:52]
  wire [7:0] _GEN_8115 = opcode_3 == 4'hf ? _GEN_6065 : _GEN_7601; // @[executor.scala 466:52]
  wire [7:0] _GEN_8116 = opcode_3 == 4'hf ? _GEN_6066 : _GEN_7602; // @[executor.scala 466:52]
  wire [7:0] _GEN_8117 = opcode_3 == 4'hf ? _GEN_6067 : _GEN_7603; // @[executor.scala 466:52]
  wire [7:0] _GEN_8118 = opcode_3 == 4'hf ? _GEN_6068 : _GEN_7604; // @[executor.scala 466:52]
  wire [7:0] _GEN_8119 = opcode_3 == 4'hf ? _GEN_6069 : _GEN_7605; // @[executor.scala 466:52]
  wire [7:0] _GEN_8120 = opcode_3 == 4'hf ? _GEN_6070 : _GEN_7606; // @[executor.scala 466:52]
  wire [7:0] _GEN_8121 = opcode_3 == 4'hf ? _GEN_6071 : _GEN_7607; // @[executor.scala 466:52]
  wire [7:0] _GEN_8122 = opcode_3 == 4'hf ? _GEN_6072 : _GEN_7608; // @[executor.scala 466:52]
  wire [7:0] _GEN_8123 = opcode_3 == 4'hf ? _GEN_6073 : _GEN_7609; // @[executor.scala 466:52]
  wire [7:0] _GEN_8124 = opcode_3 == 4'hf ? _GEN_6074 : _GEN_7610; // @[executor.scala 466:52]
  wire [7:0] _GEN_8125 = opcode_3 == 4'hf ? _GEN_6075 : _GEN_7611; // @[executor.scala 466:52]
  wire [7:0] _GEN_8126 = opcode_3 == 4'hf ? _GEN_6076 : _GEN_7612; // @[executor.scala 466:52]
  wire [7:0] _GEN_8127 = opcode_3 == 4'hf ? _GEN_6077 : _GEN_7613; // @[executor.scala 466:52]
  wire [7:0] _GEN_8128 = opcode_3 == 4'hf ? _GEN_6078 : _GEN_7614; // @[executor.scala 466:52]
  wire [7:0] _GEN_8129 = opcode_3 == 4'hf ? _GEN_6079 : _GEN_7615; // @[executor.scala 466:52]
  wire [7:0] _GEN_8130 = opcode_3 == 4'hf ? _GEN_6080 : _GEN_7616; // @[executor.scala 466:52]
  wire [7:0] _GEN_8131 = opcode_3 == 4'hf ? _GEN_6081 : _GEN_7617; // @[executor.scala 466:52]
  wire [7:0] _GEN_8132 = opcode_3 == 4'hf ? _GEN_6082 : _GEN_7618; // @[executor.scala 466:52]
  wire [7:0] _GEN_8133 = opcode_3 == 4'hf ? _GEN_6083 : _GEN_7619; // @[executor.scala 466:52]
  wire [7:0] _GEN_8134 = opcode_3 == 4'hf ? _GEN_6084 : _GEN_7620; // @[executor.scala 466:52]
  wire [7:0] _GEN_8135 = opcode_3 == 4'hf ? _GEN_6085 : _GEN_7621; // @[executor.scala 466:52]
  wire [7:0] _GEN_8136 = opcode_3 == 4'hf ? _GEN_6086 : _GEN_7622; // @[executor.scala 466:52]
  wire [7:0] _GEN_8137 = opcode_3 == 4'hf ? _GEN_6087 : _GEN_7623; // @[executor.scala 466:52]
  wire [7:0] _GEN_8138 = opcode_3 == 4'hf ? _GEN_6088 : _GEN_7624; // @[executor.scala 466:52]
  wire [7:0] _GEN_8139 = opcode_3 == 4'hf ? _GEN_6089 : _GEN_7625; // @[executor.scala 466:52]
  wire [7:0] _GEN_8140 = opcode_3 == 4'hf ? _GEN_6090 : _GEN_7626; // @[executor.scala 466:52]
  wire [7:0] _GEN_8141 = opcode_3 == 4'hf ? _GEN_6091 : _GEN_7627; // @[executor.scala 466:52]
  wire [7:0] _GEN_8142 = opcode_3 == 4'hf ? _GEN_6092 : _GEN_7628; // @[executor.scala 466:52]
  wire [7:0] _GEN_8143 = opcode_3 == 4'hf ? _GEN_6093 : _GEN_7629; // @[executor.scala 466:52]
  wire [7:0] _GEN_8144 = opcode_3 == 4'hf ? _GEN_6094 : _GEN_7630; // @[executor.scala 466:52]
  wire [7:0] _GEN_8145 = opcode_3 == 4'hf ? _GEN_6095 : _GEN_7631; // @[executor.scala 466:52]
  wire [7:0] _GEN_8146 = opcode_3 == 4'hf ? _GEN_6096 : _GEN_7632; // @[executor.scala 466:52]
  wire [7:0] _GEN_8147 = opcode_3 == 4'hf ? _GEN_6097 : _GEN_7633; // @[executor.scala 466:52]
  wire [7:0] _GEN_8148 = opcode_3 == 4'hf ? _GEN_6098 : _GEN_7634; // @[executor.scala 466:52]
  wire [7:0] _GEN_8149 = opcode_3 == 4'hf ? _GEN_6099 : _GEN_7635; // @[executor.scala 466:52]
  wire [7:0] _GEN_8150 = opcode_3 == 4'hf ? _GEN_6100 : _GEN_7636; // @[executor.scala 466:52]
  wire [7:0] _GEN_8151 = opcode_3 == 4'hf ? _GEN_6101 : _GEN_7637; // @[executor.scala 466:52]
  wire [7:0] _GEN_8152 = opcode_3 == 4'hf ? _GEN_6102 : _GEN_7638; // @[executor.scala 466:52]
  wire [7:0] _GEN_8153 = opcode_3 == 4'hf ? _GEN_6103 : _GEN_7639; // @[executor.scala 466:52]
  wire [7:0] _GEN_8154 = opcode_3 == 4'hf ? _GEN_6104 : _GEN_7640; // @[executor.scala 466:52]
  wire [7:0] _GEN_8155 = opcode_3 == 4'hf ? _GEN_6105 : _GEN_7641; // @[executor.scala 466:52]
  wire [7:0] _GEN_8156 = opcode_3 == 4'hf ? _GEN_6106 : _GEN_7642; // @[executor.scala 466:52]
  wire [7:0] _GEN_8157 = opcode_3 == 4'hf ? _GEN_6107 : _GEN_7643; // @[executor.scala 466:52]
  wire [7:0] _GEN_8158 = opcode_3 == 4'hf ? _GEN_6108 : _GEN_7644; // @[executor.scala 466:52]
  wire [7:0] _GEN_8159 = opcode_3 == 4'hf ? _GEN_6109 : _GEN_7645; // @[executor.scala 466:52]
  wire [7:0] _GEN_8160 = opcode_3 == 4'hf ? _GEN_6110 : _GEN_7646; // @[executor.scala 466:52]
  wire [7:0] _GEN_8161 = opcode_3 == 4'hf ? _GEN_6111 : _GEN_7647; // @[executor.scala 466:52]
  wire [7:0] _GEN_8162 = opcode_3 == 4'hf ? _GEN_6112 : _GEN_7648; // @[executor.scala 466:52]
  wire [7:0] _GEN_8163 = opcode_3 == 4'hf ? _GEN_6113 : _GEN_7649; // @[executor.scala 466:52]
  wire [7:0] _GEN_8164 = opcode_3 == 4'hf ? _GEN_6114 : _GEN_7650; // @[executor.scala 466:52]
  wire [7:0] _GEN_8165 = opcode_3 == 4'hf ? _GEN_6115 : _GEN_7651; // @[executor.scala 466:52]
  wire [7:0] _GEN_8166 = opcode_3 == 4'hf ? _GEN_6116 : _GEN_7652; // @[executor.scala 466:52]
  wire [7:0] _GEN_8167 = opcode_3 == 4'hf ? _GEN_6117 : _GEN_7653; // @[executor.scala 466:52]
  wire [7:0] _GEN_8168 = opcode_3 == 4'hf ? _GEN_6118 : _GEN_7654; // @[executor.scala 466:52]
  wire [7:0] _GEN_8169 = opcode_3 == 4'hf ? _GEN_6119 : _GEN_7655; // @[executor.scala 466:52]
  wire [7:0] _GEN_8170 = opcode_3 == 4'hf ? _GEN_6120 : _GEN_7656; // @[executor.scala 466:52]
  wire [7:0] _GEN_8171 = opcode_3 == 4'hf ? _GEN_6121 : _GEN_7657; // @[executor.scala 466:52]
  wire [7:0] _GEN_8172 = opcode_3 == 4'hf ? _GEN_6122 : _GEN_7658; // @[executor.scala 466:52]
  wire [7:0] _GEN_8173 = opcode_3 == 4'hf ? _GEN_6123 : _GEN_7659; // @[executor.scala 466:52]
  wire [7:0] _GEN_8174 = opcode_3 == 4'hf ? _GEN_6124 : _GEN_7660; // @[executor.scala 466:52]
  wire [7:0] _GEN_8175 = opcode_3 == 4'hf ? _GEN_6125 : _GEN_7661; // @[executor.scala 466:52]
  wire [7:0] _GEN_8176 = opcode_3 == 4'hf ? _GEN_6126 : _GEN_7662; // @[executor.scala 466:52]
  wire [7:0] _GEN_8177 = opcode_3 == 4'hf ? _GEN_6127 : _GEN_7663; // @[executor.scala 466:52]
  wire [7:0] _GEN_8178 = opcode_3 == 4'hf ? _GEN_6128 : _GEN_7664; // @[executor.scala 466:52]
  wire [7:0] _GEN_8179 = opcode_3 == 4'hf ? _GEN_6129 : _GEN_7665; // @[executor.scala 466:52]
  wire [7:0] _GEN_8180 = opcode_3 == 4'hf ? _GEN_6130 : _GEN_7666; // @[executor.scala 466:52]
  wire [7:0] _GEN_8181 = opcode_3 == 4'hf ? _GEN_6131 : _GEN_7667; // @[executor.scala 466:52]
  wire [7:0] _GEN_8182 = opcode_3 == 4'hf ? _GEN_6132 : _GEN_7668; // @[executor.scala 466:52]
  wire [7:0] _GEN_8183 = opcode_3 == 4'hf ? _GEN_6133 : _GEN_7669; // @[executor.scala 466:52]
  wire [7:0] _GEN_8184 = opcode_3 == 4'hf ? _GEN_6134 : _GEN_7670; // @[executor.scala 466:52]
  wire [7:0] _GEN_8185 = opcode_3 == 4'hf ? _GEN_6135 : _GEN_7671; // @[executor.scala 466:52]
  wire [7:0] _GEN_8186 = opcode_3 == 4'hf ? _GEN_6136 : _GEN_7672; // @[executor.scala 466:52]
  wire [7:0] _GEN_8187 = opcode_3 == 4'hf ? _GEN_6137 : _GEN_7673; // @[executor.scala 466:52]
  wire [7:0] _GEN_8188 = opcode_3 == 4'hf ? _GEN_6138 : _GEN_7674; // @[executor.scala 466:52]
  wire [7:0] _GEN_8189 = opcode_3 == 4'hf ? _GEN_6139 : _GEN_7675; // @[executor.scala 466:52]
  wire [7:0] _GEN_8190 = opcode_3 == 4'hf ? _GEN_6140 : _GEN_7676; // @[executor.scala 466:52]
  wire [7:0] _GEN_8191 = opcode_3 == 4'hf ? _GEN_6141 : _GEN_7677; // @[executor.scala 466:52]
  wire [7:0] _GEN_8192 = opcode_3 == 4'hf ? _GEN_6142 : _GEN_7678; // @[executor.scala 466:52]
  wire [7:0] _GEN_8193 = opcode_3 == 4'hf ? _GEN_6143 : _GEN_7679; // @[executor.scala 466:52]
  wire [7:0] _GEN_8194 = opcode_3 == 4'hf ? _GEN_6144 : _GEN_7680; // @[executor.scala 466:52]
  wire [7:0] _GEN_8195 = opcode_3 == 4'hf ? _GEN_6145 : _GEN_7681; // @[executor.scala 466:52]
  wire [7:0] _GEN_8196 = opcode_3 == 4'hf ? _GEN_6146 : _GEN_7682; // @[executor.scala 466:52]
  wire [7:0] _GEN_8197 = opcode_3 == 4'hf ? _GEN_6147 : _GEN_7683; // @[executor.scala 466:52]
  wire [7:0] _GEN_8198 = opcode_3 == 4'hf ? _GEN_6148 : _GEN_7684; // @[executor.scala 466:52]
  wire [7:0] _GEN_8199 = opcode_3 == 4'hf ? _GEN_6149 : _GEN_7685; // @[executor.scala 466:52]
  assign io_pipe_phv_out_data_0 = phv_is_valid_processor ? _GEN_7691 : phv_data_0; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_1 = phv_is_valid_processor ? _GEN_7690 : phv_data_1; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_2 = phv_is_valid_processor ? _GEN_7689 : phv_data_2; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_3 = phv_is_valid_processor ? _GEN_7688 : phv_data_3; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_4 = phv_is_valid_processor ? _GEN_7695 : phv_data_4; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_5 = phv_is_valid_processor ? _GEN_7694 : phv_data_5; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_6 = phv_is_valid_processor ? _GEN_7693 : phv_data_6; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_7 = phv_is_valid_processor ? _GEN_7692 : phv_data_7; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_8 = phv_is_valid_processor ? _GEN_7699 : phv_data_8; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_9 = phv_is_valid_processor ? _GEN_7698 : phv_data_9; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_10 = phv_is_valid_processor ? _GEN_7697 : phv_data_10; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_11 = phv_is_valid_processor ? _GEN_7696 : phv_data_11; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_12 = phv_is_valid_processor ? _GEN_7703 : phv_data_12; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_13 = phv_is_valid_processor ? _GEN_7702 : phv_data_13; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_14 = phv_is_valid_processor ? _GEN_7701 : phv_data_14; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_15 = phv_is_valid_processor ? _GEN_7700 : phv_data_15; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_16 = phv_is_valid_processor ? _GEN_7707 : phv_data_16; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_17 = phv_is_valid_processor ? _GEN_7706 : phv_data_17; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_18 = phv_is_valid_processor ? _GEN_7705 : phv_data_18; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_19 = phv_is_valid_processor ? _GEN_7704 : phv_data_19; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_20 = phv_is_valid_processor ? _GEN_7711 : phv_data_20; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_21 = phv_is_valid_processor ? _GEN_7710 : phv_data_21; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_22 = phv_is_valid_processor ? _GEN_7709 : phv_data_22; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_23 = phv_is_valid_processor ? _GEN_7708 : phv_data_23; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_24 = phv_is_valid_processor ? _GEN_7715 : phv_data_24; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_25 = phv_is_valid_processor ? _GEN_7714 : phv_data_25; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_26 = phv_is_valid_processor ? _GEN_7713 : phv_data_26; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_27 = phv_is_valid_processor ? _GEN_7712 : phv_data_27; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_28 = phv_is_valid_processor ? _GEN_7719 : phv_data_28; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_29 = phv_is_valid_processor ? _GEN_7718 : phv_data_29; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_30 = phv_is_valid_processor ? _GEN_7717 : phv_data_30; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_31 = phv_is_valid_processor ? _GEN_7716 : phv_data_31; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_32 = phv_is_valid_processor ? _GEN_7723 : phv_data_32; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_33 = phv_is_valid_processor ? _GEN_7722 : phv_data_33; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_34 = phv_is_valid_processor ? _GEN_7721 : phv_data_34; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_35 = phv_is_valid_processor ? _GEN_7720 : phv_data_35; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_36 = phv_is_valid_processor ? _GEN_7727 : phv_data_36; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_37 = phv_is_valid_processor ? _GEN_7726 : phv_data_37; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_38 = phv_is_valid_processor ? _GEN_7725 : phv_data_38; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_39 = phv_is_valid_processor ? _GEN_7724 : phv_data_39; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_40 = phv_is_valid_processor ? _GEN_7731 : phv_data_40; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_41 = phv_is_valid_processor ? _GEN_7730 : phv_data_41; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_42 = phv_is_valid_processor ? _GEN_7729 : phv_data_42; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_43 = phv_is_valid_processor ? _GEN_7728 : phv_data_43; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_44 = phv_is_valid_processor ? _GEN_7735 : phv_data_44; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_45 = phv_is_valid_processor ? _GEN_7734 : phv_data_45; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_46 = phv_is_valid_processor ? _GEN_7733 : phv_data_46; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_47 = phv_is_valid_processor ? _GEN_7732 : phv_data_47; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_48 = phv_is_valid_processor ? _GEN_7739 : phv_data_48; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_49 = phv_is_valid_processor ? _GEN_7738 : phv_data_49; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_50 = phv_is_valid_processor ? _GEN_7737 : phv_data_50; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_51 = phv_is_valid_processor ? _GEN_7736 : phv_data_51; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_52 = phv_is_valid_processor ? _GEN_7743 : phv_data_52; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_53 = phv_is_valid_processor ? _GEN_7742 : phv_data_53; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_54 = phv_is_valid_processor ? _GEN_7741 : phv_data_54; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_55 = phv_is_valid_processor ? _GEN_7740 : phv_data_55; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_56 = phv_is_valid_processor ? _GEN_7747 : phv_data_56; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_57 = phv_is_valid_processor ? _GEN_7746 : phv_data_57; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_58 = phv_is_valid_processor ? _GEN_7745 : phv_data_58; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_59 = phv_is_valid_processor ? _GEN_7744 : phv_data_59; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_60 = phv_is_valid_processor ? _GEN_7751 : phv_data_60; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_61 = phv_is_valid_processor ? _GEN_7750 : phv_data_61; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_62 = phv_is_valid_processor ? _GEN_7749 : phv_data_62; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_63 = phv_is_valid_processor ? _GEN_7748 : phv_data_63; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_64 = phv_is_valid_processor ? _GEN_7755 : phv_data_64; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_65 = phv_is_valid_processor ? _GEN_7754 : phv_data_65; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_66 = phv_is_valid_processor ? _GEN_7753 : phv_data_66; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_67 = phv_is_valid_processor ? _GEN_7752 : phv_data_67; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_68 = phv_is_valid_processor ? _GEN_7759 : phv_data_68; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_69 = phv_is_valid_processor ? _GEN_7758 : phv_data_69; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_70 = phv_is_valid_processor ? _GEN_7757 : phv_data_70; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_71 = phv_is_valid_processor ? _GEN_7756 : phv_data_71; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_72 = phv_is_valid_processor ? _GEN_7763 : phv_data_72; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_73 = phv_is_valid_processor ? _GEN_7762 : phv_data_73; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_74 = phv_is_valid_processor ? _GEN_7761 : phv_data_74; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_75 = phv_is_valid_processor ? _GEN_7760 : phv_data_75; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_76 = phv_is_valid_processor ? _GEN_7767 : phv_data_76; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_77 = phv_is_valid_processor ? _GEN_7766 : phv_data_77; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_78 = phv_is_valid_processor ? _GEN_7765 : phv_data_78; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_79 = phv_is_valid_processor ? _GEN_7764 : phv_data_79; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_80 = phv_is_valid_processor ? _GEN_7771 : phv_data_80; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_81 = phv_is_valid_processor ? _GEN_7770 : phv_data_81; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_82 = phv_is_valid_processor ? _GEN_7769 : phv_data_82; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_83 = phv_is_valid_processor ? _GEN_7768 : phv_data_83; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_84 = phv_is_valid_processor ? _GEN_7775 : phv_data_84; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_85 = phv_is_valid_processor ? _GEN_7774 : phv_data_85; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_86 = phv_is_valid_processor ? _GEN_7773 : phv_data_86; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_87 = phv_is_valid_processor ? _GEN_7772 : phv_data_87; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_88 = phv_is_valid_processor ? _GEN_7779 : phv_data_88; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_89 = phv_is_valid_processor ? _GEN_7778 : phv_data_89; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_90 = phv_is_valid_processor ? _GEN_7777 : phv_data_90; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_91 = phv_is_valid_processor ? _GEN_7776 : phv_data_91; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_92 = phv_is_valid_processor ? _GEN_7783 : phv_data_92; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_93 = phv_is_valid_processor ? _GEN_7782 : phv_data_93; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_94 = phv_is_valid_processor ? _GEN_7781 : phv_data_94; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_95 = phv_is_valid_processor ? _GEN_7780 : phv_data_95; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_96 = phv_is_valid_processor ? _GEN_7787 : phv_data_96; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_97 = phv_is_valid_processor ? _GEN_7786 : phv_data_97; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_98 = phv_is_valid_processor ? _GEN_7785 : phv_data_98; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_99 = phv_is_valid_processor ? _GEN_7784 : phv_data_99; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_100 = phv_is_valid_processor ? _GEN_7791 : phv_data_100; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_101 = phv_is_valid_processor ? _GEN_7790 : phv_data_101; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_102 = phv_is_valid_processor ? _GEN_7789 : phv_data_102; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_103 = phv_is_valid_processor ? _GEN_7788 : phv_data_103; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_104 = phv_is_valid_processor ? _GEN_7795 : phv_data_104; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_105 = phv_is_valid_processor ? _GEN_7794 : phv_data_105; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_106 = phv_is_valid_processor ? _GEN_7793 : phv_data_106; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_107 = phv_is_valid_processor ? _GEN_7792 : phv_data_107; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_108 = phv_is_valid_processor ? _GEN_7799 : phv_data_108; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_109 = phv_is_valid_processor ? _GEN_7798 : phv_data_109; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_110 = phv_is_valid_processor ? _GEN_7797 : phv_data_110; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_111 = phv_is_valid_processor ? _GEN_7796 : phv_data_111; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_112 = phv_is_valid_processor ? _GEN_7803 : phv_data_112; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_113 = phv_is_valid_processor ? _GEN_7802 : phv_data_113; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_114 = phv_is_valid_processor ? _GEN_7801 : phv_data_114; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_115 = phv_is_valid_processor ? _GEN_7800 : phv_data_115; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_116 = phv_is_valid_processor ? _GEN_7807 : phv_data_116; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_117 = phv_is_valid_processor ? _GEN_7806 : phv_data_117; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_118 = phv_is_valid_processor ? _GEN_7805 : phv_data_118; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_119 = phv_is_valid_processor ? _GEN_7804 : phv_data_119; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_120 = phv_is_valid_processor ? _GEN_7811 : phv_data_120; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_121 = phv_is_valid_processor ? _GEN_7810 : phv_data_121; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_122 = phv_is_valid_processor ? _GEN_7809 : phv_data_122; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_123 = phv_is_valid_processor ? _GEN_7808 : phv_data_123; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_124 = phv_is_valid_processor ? _GEN_7815 : phv_data_124; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_125 = phv_is_valid_processor ? _GEN_7814 : phv_data_125; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_126 = phv_is_valid_processor ? _GEN_7813 : phv_data_126; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_127 = phv_is_valid_processor ? _GEN_7812 : phv_data_127; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_128 = phv_is_valid_processor ? _GEN_7819 : phv_data_128; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_129 = phv_is_valid_processor ? _GEN_7818 : phv_data_129; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_130 = phv_is_valid_processor ? _GEN_7817 : phv_data_130; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_131 = phv_is_valid_processor ? _GEN_7816 : phv_data_131; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_132 = phv_is_valid_processor ? _GEN_7823 : phv_data_132; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_133 = phv_is_valid_processor ? _GEN_7822 : phv_data_133; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_134 = phv_is_valid_processor ? _GEN_7821 : phv_data_134; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_135 = phv_is_valid_processor ? _GEN_7820 : phv_data_135; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_136 = phv_is_valid_processor ? _GEN_7827 : phv_data_136; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_137 = phv_is_valid_processor ? _GEN_7826 : phv_data_137; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_138 = phv_is_valid_processor ? _GEN_7825 : phv_data_138; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_139 = phv_is_valid_processor ? _GEN_7824 : phv_data_139; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_140 = phv_is_valid_processor ? _GEN_7831 : phv_data_140; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_141 = phv_is_valid_processor ? _GEN_7830 : phv_data_141; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_142 = phv_is_valid_processor ? _GEN_7829 : phv_data_142; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_143 = phv_is_valid_processor ? _GEN_7828 : phv_data_143; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_144 = phv_is_valid_processor ? _GEN_7835 : phv_data_144; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_145 = phv_is_valid_processor ? _GEN_7834 : phv_data_145; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_146 = phv_is_valid_processor ? _GEN_7833 : phv_data_146; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_147 = phv_is_valid_processor ? _GEN_7832 : phv_data_147; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_148 = phv_is_valid_processor ? _GEN_7839 : phv_data_148; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_149 = phv_is_valid_processor ? _GEN_7838 : phv_data_149; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_150 = phv_is_valid_processor ? _GEN_7837 : phv_data_150; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_151 = phv_is_valid_processor ? _GEN_7836 : phv_data_151; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_152 = phv_is_valid_processor ? _GEN_7843 : phv_data_152; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_153 = phv_is_valid_processor ? _GEN_7842 : phv_data_153; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_154 = phv_is_valid_processor ? _GEN_7841 : phv_data_154; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_155 = phv_is_valid_processor ? _GEN_7840 : phv_data_155; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_156 = phv_is_valid_processor ? _GEN_7847 : phv_data_156; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_157 = phv_is_valid_processor ? _GEN_7846 : phv_data_157; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_158 = phv_is_valid_processor ? _GEN_7845 : phv_data_158; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_159 = phv_is_valid_processor ? _GEN_7844 : phv_data_159; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_160 = phv_is_valid_processor ? _GEN_7851 : phv_data_160; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_161 = phv_is_valid_processor ? _GEN_7850 : phv_data_161; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_162 = phv_is_valid_processor ? _GEN_7849 : phv_data_162; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_163 = phv_is_valid_processor ? _GEN_7848 : phv_data_163; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_164 = phv_is_valid_processor ? _GEN_7855 : phv_data_164; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_165 = phv_is_valid_processor ? _GEN_7854 : phv_data_165; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_166 = phv_is_valid_processor ? _GEN_7853 : phv_data_166; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_167 = phv_is_valid_processor ? _GEN_7852 : phv_data_167; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_168 = phv_is_valid_processor ? _GEN_7859 : phv_data_168; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_169 = phv_is_valid_processor ? _GEN_7858 : phv_data_169; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_170 = phv_is_valid_processor ? _GEN_7857 : phv_data_170; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_171 = phv_is_valid_processor ? _GEN_7856 : phv_data_171; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_172 = phv_is_valid_processor ? _GEN_7863 : phv_data_172; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_173 = phv_is_valid_processor ? _GEN_7862 : phv_data_173; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_174 = phv_is_valid_processor ? _GEN_7861 : phv_data_174; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_175 = phv_is_valid_processor ? _GEN_7860 : phv_data_175; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_176 = phv_is_valid_processor ? _GEN_7867 : phv_data_176; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_177 = phv_is_valid_processor ? _GEN_7866 : phv_data_177; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_178 = phv_is_valid_processor ? _GEN_7865 : phv_data_178; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_179 = phv_is_valid_processor ? _GEN_7864 : phv_data_179; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_180 = phv_is_valid_processor ? _GEN_7871 : phv_data_180; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_181 = phv_is_valid_processor ? _GEN_7870 : phv_data_181; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_182 = phv_is_valid_processor ? _GEN_7869 : phv_data_182; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_183 = phv_is_valid_processor ? _GEN_7868 : phv_data_183; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_184 = phv_is_valid_processor ? _GEN_7875 : phv_data_184; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_185 = phv_is_valid_processor ? _GEN_7874 : phv_data_185; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_186 = phv_is_valid_processor ? _GEN_7873 : phv_data_186; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_187 = phv_is_valid_processor ? _GEN_7872 : phv_data_187; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_188 = phv_is_valid_processor ? _GEN_7879 : phv_data_188; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_189 = phv_is_valid_processor ? _GEN_7878 : phv_data_189; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_190 = phv_is_valid_processor ? _GEN_7877 : phv_data_190; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_191 = phv_is_valid_processor ? _GEN_7876 : phv_data_191; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_192 = phv_is_valid_processor ? _GEN_7883 : phv_data_192; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_193 = phv_is_valid_processor ? _GEN_7882 : phv_data_193; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_194 = phv_is_valid_processor ? _GEN_7881 : phv_data_194; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_195 = phv_is_valid_processor ? _GEN_7880 : phv_data_195; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_196 = phv_is_valid_processor ? _GEN_7887 : phv_data_196; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_197 = phv_is_valid_processor ? _GEN_7886 : phv_data_197; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_198 = phv_is_valid_processor ? _GEN_7885 : phv_data_198; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_199 = phv_is_valid_processor ? _GEN_7884 : phv_data_199; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_200 = phv_is_valid_processor ? _GEN_7891 : phv_data_200; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_201 = phv_is_valid_processor ? _GEN_7890 : phv_data_201; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_202 = phv_is_valid_processor ? _GEN_7889 : phv_data_202; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_203 = phv_is_valid_processor ? _GEN_7888 : phv_data_203; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_204 = phv_is_valid_processor ? _GEN_7895 : phv_data_204; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_205 = phv_is_valid_processor ? _GEN_7894 : phv_data_205; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_206 = phv_is_valid_processor ? _GEN_7893 : phv_data_206; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_207 = phv_is_valid_processor ? _GEN_7892 : phv_data_207; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_208 = phv_is_valid_processor ? _GEN_7899 : phv_data_208; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_209 = phv_is_valid_processor ? _GEN_7898 : phv_data_209; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_210 = phv_is_valid_processor ? _GEN_7897 : phv_data_210; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_211 = phv_is_valid_processor ? _GEN_7896 : phv_data_211; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_212 = phv_is_valid_processor ? _GEN_7903 : phv_data_212; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_213 = phv_is_valid_processor ? _GEN_7902 : phv_data_213; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_214 = phv_is_valid_processor ? _GEN_7901 : phv_data_214; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_215 = phv_is_valid_processor ? _GEN_7900 : phv_data_215; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_216 = phv_is_valid_processor ? _GEN_7907 : phv_data_216; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_217 = phv_is_valid_processor ? _GEN_7906 : phv_data_217; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_218 = phv_is_valid_processor ? _GEN_7905 : phv_data_218; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_219 = phv_is_valid_processor ? _GEN_7904 : phv_data_219; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_220 = phv_is_valid_processor ? _GEN_7911 : phv_data_220; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_221 = phv_is_valid_processor ? _GEN_7910 : phv_data_221; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_222 = phv_is_valid_processor ? _GEN_7909 : phv_data_222; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_223 = phv_is_valid_processor ? _GEN_7908 : phv_data_223; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_224 = phv_is_valid_processor ? _GEN_7915 : phv_data_224; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_225 = phv_is_valid_processor ? _GEN_7914 : phv_data_225; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_226 = phv_is_valid_processor ? _GEN_7913 : phv_data_226; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_227 = phv_is_valid_processor ? _GEN_7912 : phv_data_227; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_228 = phv_is_valid_processor ? _GEN_7919 : phv_data_228; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_229 = phv_is_valid_processor ? _GEN_7918 : phv_data_229; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_230 = phv_is_valid_processor ? _GEN_7917 : phv_data_230; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_231 = phv_is_valid_processor ? _GEN_7916 : phv_data_231; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_232 = phv_is_valid_processor ? _GEN_7923 : phv_data_232; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_233 = phv_is_valid_processor ? _GEN_7922 : phv_data_233; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_234 = phv_is_valid_processor ? _GEN_7921 : phv_data_234; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_235 = phv_is_valid_processor ? _GEN_7920 : phv_data_235; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_236 = phv_is_valid_processor ? _GEN_7927 : phv_data_236; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_237 = phv_is_valid_processor ? _GEN_7926 : phv_data_237; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_238 = phv_is_valid_processor ? _GEN_7925 : phv_data_238; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_239 = phv_is_valid_processor ? _GEN_7924 : phv_data_239; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_240 = phv_is_valid_processor ? _GEN_7931 : phv_data_240; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_241 = phv_is_valid_processor ? _GEN_7930 : phv_data_241; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_242 = phv_is_valid_processor ? _GEN_7929 : phv_data_242; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_243 = phv_is_valid_processor ? _GEN_7928 : phv_data_243; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_244 = phv_is_valid_processor ? _GEN_7935 : phv_data_244; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_245 = phv_is_valid_processor ? _GEN_7934 : phv_data_245; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_246 = phv_is_valid_processor ? _GEN_7933 : phv_data_246; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_247 = phv_is_valid_processor ? _GEN_7932 : phv_data_247; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_248 = phv_is_valid_processor ? _GEN_7939 : phv_data_248; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_249 = phv_is_valid_processor ? _GEN_7938 : phv_data_249; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_250 = phv_is_valid_processor ? _GEN_7937 : phv_data_250; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_251 = phv_is_valid_processor ? _GEN_7936 : phv_data_251; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_252 = phv_is_valid_processor ? _GEN_7943 : phv_data_252; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_253 = phv_is_valid_processor ? _GEN_7942 : phv_data_253; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_254 = phv_is_valid_processor ? _GEN_7941 : phv_data_254; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_255 = phv_is_valid_processor ? _GEN_7940 : phv_data_255; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_256 = phv_is_valid_processor ? _GEN_7947 : phv_data_256; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_257 = phv_is_valid_processor ? _GEN_7946 : phv_data_257; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_258 = phv_is_valid_processor ? _GEN_7945 : phv_data_258; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_259 = phv_is_valid_processor ? _GEN_7944 : phv_data_259; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_260 = phv_is_valid_processor ? _GEN_7951 : phv_data_260; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_261 = phv_is_valid_processor ? _GEN_7950 : phv_data_261; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_262 = phv_is_valid_processor ? _GEN_7949 : phv_data_262; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_263 = phv_is_valid_processor ? _GEN_7948 : phv_data_263; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_264 = phv_is_valid_processor ? _GEN_7955 : phv_data_264; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_265 = phv_is_valid_processor ? _GEN_7954 : phv_data_265; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_266 = phv_is_valid_processor ? _GEN_7953 : phv_data_266; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_267 = phv_is_valid_processor ? _GEN_7952 : phv_data_267; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_268 = phv_is_valid_processor ? _GEN_7959 : phv_data_268; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_269 = phv_is_valid_processor ? _GEN_7958 : phv_data_269; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_270 = phv_is_valid_processor ? _GEN_7957 : phv_data_270; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_271 = phv_is_valid_processor ? _GEN_7956 : phv_data_271; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_272 = phv_is_valid_processor ? _GEN_7963 : phv_data_272; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_273 = phv_is_valid_processor ? _GEN_7962 : phv_data_273; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_274 = phv_is_valid_processor ? _GEN_7961 : phv_data_274; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_275 = phv_is_valid_processor ? _GEN_7960 : phv_data_275; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_276 = phv_is_valid_processor ? _GEN_7967 : phv_data_276; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_277 = phv_is_valid_processor ? _GEN_7966 : phv_data_277; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_278 = phv_is_valid_processor ? _GEN_7965 : phv_data_278; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_279 = phv_is_valid_processor ? _GEN_7964 : phv_data_279; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_280 = phv_is_valid_processor ? _GEN_7971 : phv_data_280; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_281 = phv_is_valid_processor ? _GEN_7970 : phv_data_281; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_282 = phv_is_valid_processor ? _GEN_7969 : phv_data_282; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_283 = phv_is_valid_processor ? _GEN_7968 : phv_data_283; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_284 = phv_is_valid_processor ? _GEN_7975 : phv_data_284; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_285 = phv_is_valid_processor ? _GEN_7974 : phv_data_285; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_286 = phv_is_valid_processor ? _GEN_7973 : phv_data_286; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_287 = phv_is_valid_processor ? _GEN_7972 : phv_data_287; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_288 = phv_is_valid_processor ? _GEN_7979 : phv_data_288; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_289 = phv_is_valid_processor ? _GEN_7978 : phv_data_289; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_290 = phv_is_valid_processor ? _GEN_7977 : phv_data_290; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_291 = phv_is_valid_processor ? _GEN_7976 : phv_data_291; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_292 = phv_is_valid_processor ? _GEN_7983 : phv_data_292; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_293 = phv_is_valid_processor ? _GEN_7982 : phv_data_293; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_294 = phv_is_valid_processor ? _GEN_7981 : phv_data_294; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_295 = phv_is_valid_processor ? _GEN_7980 : phv_data_295; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_296 = phv_is_valid_processor ? _GEN_7987 : phv_data_296; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_297 = phv_is_valid_processor ? _GEN_7986 : phv_data_297; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_298 = phv_is_valid_processor ? _GEN_7985 : phv_data_298; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_299 = phv_is_valid_processor ? _GEN_7984 : phv_data_299; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_300 = phv_is_valid_processor ? _GEN_7991 : phv_data_300; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_301 = phv_is_valid_processor ? _GEN_7990 : phv_data_301; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_302 = phv_is_valid_processor ? _GEN_7989 : phv_data_302; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_303 = phv_is_valid_processor ? _GEN_7988 : phv_data_303; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_304 = phv_is_valid_processor ? _GEN_7995 : phv_data_304; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_305 = phv_is_valid_processor ? _GEN_7994 : phv_data_305; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_306 = phv_is_valid_processor ? _GEN_7993 : phv_data_306; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_307 = phv_is_valid_processor ? _GEN_7992 : phv_data_307; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_308 = phv_is_valid_processor ? _GEN_7999 : phv_data_308; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_309 = phv_is_valid_processor ? _GEN_7998 : phv_data_309; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_310 = phv_is_valid_processor ? _GEN_7997 : phv_data_310; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_311 = phv_is_valid_processor ? _GEN_7996 : phv_data_311; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_312 = phv_is_valid_processor ? _GEN_8003 : phv_data_312; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_313 = phv_is_valid_processor ? _GEN_8002 : phv_data_313; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_314 = phv_is_valid_processor ? _GEN_8001 : phv_data_314; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_315 = phv_is_valid_processor ? _GEN_8000 : phv_data_315; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_316 = phv_is_valid_processor ? _GEN_8007 : phv_data_316; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_317 = phv_is_valid_processor ? _GEN_8006 : phv_data_317; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_318 = phv_is_valid_processor ? _GEN_8005 : phv_data_318; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_319 = phv_is_valid_processor ? _GEN_8004 : phv_data_319; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_320 = phv_is_valid_processor ? _GEN_8011 : phv_data_320; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_321 = phv_is_valid_processor ? _GEN_8010 : phv_data_321; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_322 = phv_is_valid_processor ? _GEN_8009 : phv_data_322; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_323 = phv_is_valid_processor ? _GEN_8008 : phv_data_323; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_324 = phv_is_valid_processor ? _GEN_8015 : phv_data_324; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_325 = phv_is_valid_processor ? _GEN_8014 : phv_data_325; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_326 = phv_is_valid_processor ? _GEN_8013 : phv_data_326; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_327 = phv_is_valid_processor ? _GEN_8012 : phv_data_327; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_328 = phv_is_valid_processor ? _GEN_8019 : phv_data_328; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_329 = phv_is_valid_processor ? _GEN_8018 : phv_data_329; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_330 = phv_is_valid_processor ? _GEN_8017 : phv_data_330; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_331 = phv_is_valid_processor ? _GEN_8016 : phv_data_331; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_332 = phv_is_valid_processor ? _GEN_8023 : phv_data_332; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_333 = phv_is_valid_processor ? _GEN_8022 : phv_data_333; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_334 = phv_is_valid_processor ? _GEN_8021 : phv_data_334; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_335 = phv_is_valid_processor ? _GEN_8020 : phv_data_335; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_336 = phv_is_valid_processor ? _GEN_8027 : phv_data_336; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_337 = phv_is_valid_processor ? _GEN_8026 : phv_data_337; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_338 = phv_is_valid_processor ? _GEN_8025 : phv_data_338; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_339 = phv_is_valid_processor ? _GEN_8024 : phv_data_339; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_340 = phv_is_valid_processor ? _GEN_8031 : phv_data_340; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_341 = phv_is_valid_processor ? _GEN_8030 : phv_data_341; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_342 = phv_is_valid_processor ? _GEN_8029 : phv_data_342; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_343 = phv_is_valid_processor ? _GEN_8028 : phv_data_343; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_344 = phv_is_valid_processor ? _GEN_8035 : phv_data_344; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_345 = phv_is_valid_processor ? _GEN_8034 : phv_data_345; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_346 = phv_is_valid_processor ? _GEN_8033 : phv_data_346; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_347 = phv_is_valid_processor ? _GEN_8032 : phv_data_347; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_348 = phv_is_valid_processor ? _GEN_8039 : phv_data_348; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_349 = phv_is_valid_processor ? _GEN_8038 : phv_data_349; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_350 = phv_is_valid_processor ? _GEN_8037 : phv_data_350; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_351 = phv_is_valid_processor ? _GEN_8036 : phv_data_351; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_352 = phv_is_valid_processor ? _GEN_8043 : phv_data_352; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_353 = phv_is_valid_processor ? _GEN_8042 : phv_data_353; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_354 = phv_is_valid_processor ? _GEN_8041 : phv_data_354; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_355 = phv_is_valid_processor ? _GEN_8040 : phv_data_355; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_356 = phv_is_valid_processor ? _GEN_8047 : phv_data_356; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_357 = phv_is_valid_processor ? _GEN_8046 : phv_data_357; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_358 = phv_is_valid_processor ? _GEN_8045 : phv_data_358; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_359 = phv_is_valid_processor ? _GEN_8044 : phv_data_359; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_360 = phv_is_valid_processor ? _GEN_8051 : phv_data_360; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_361 = phv_is_valid_processor ? _GEN_8050 : phv_data_361; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_362 = phv_is_valid_processor ? _GEN_8049 : phv_data_362; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_363 = phv_is_valid_processor ? _GEN_8048 : phv_data_363; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_364 = phv_is_valid_processor ? _GEN_8055 : phv_data_364; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_365 = phv_is_valid_processor ? _GEN_8054 : phv_data_365; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_366 = phv_is_valid_processor ? _GEN_8053 : phv_data_366; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_367 = phv_is_valid_processor ? _GEN_8052 : phv_data_367; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_368 = phv_is_valid_processor ? _GEN_8059 : phv_data_368; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_369 = phv_is_valid_processor ? _GEN_8058 : phv_data_369; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_370 = phv_is_valid_processor ? _GEN_8057 : phv_data_370; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_371 = phv_is_valid_processor ? _GEN_8056 : phv_data_371; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_372 = phv_is_valid_processor ? _GEN_8063 : phv_data_372; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_373 = phv_is_valid_processor ? _GEN_8062 : phv_data_373; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_374 = phv_is_valid_processor ? _GEN_8061 : phv_data_374; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_375 = phv_is_valid_processor ? _GEN_8060 : phv_data_375; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_376 = phv_is_valid_processor ? _GEN_8067 : phv_data_376; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_377 = phv_is_valid_processor ? _GEN_8066 : phv_data_377; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_378 = phv_is_valid_processor ? _GEN_8065 : phv_data_378; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_379 = phv_is_valid_processor ? _GEN_8064 : phv_data_379; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_380 = phv_is_valid_processor ? _GEN_8071 : phv_data_380; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_381 = phv_is_valid_processor ? _GEN_8070 : phv_data_381; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_382 = phv_is_valid_processor ? _GEN_8069 : phv_data_382; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_383 = phv_is_valid_processor ? _GEN_8068 : phv_data_383; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_384 = phv_is_valid_processor ? _GEN_8075 : phv_data_384; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_385 = phv_is_valid_processor ? _GEN_8074 : phv_data_385; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_386 = phv_is_valid_processor ? _GEN_8073 : phv_data_386; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_387 = phv_is_valid_processor ? _GEN_8072 : phv_data_387; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_388 = phv_is_valid_processor ? _GEN_8079 : phv_data_388; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_389 = phv_is_valid_processor ? _GEN_8078 : phv_data_389; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_390 = phv_is_valid_processor ? _GEN_8077 : phv_data_390; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_391 = phv_is_valid_processor ? _GEN_8076 : phv_data_391; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_392 = phv_is_valid_processor ? _GEN_8083 : phv_data_392; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_393 = phv_is_valid_processor ? _GEN_8082 : phv_data_393; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_394 = phv_is_valid_processor ? _GEN_8081 : phv_data_394; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_395 = phv_is_valid_processor ? _GEN_8080 : phv_data_395; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_396 = phv_is_valid_processor ? _GEN_8087 : phv_data_396; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_397 = phv_is_valid_processor ? _GEN_8086 : phv_data_397; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_398 = phv_is_valid_processor ? _GEN_8085 : phv_data_398; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_399 = phv_is_valid_processor ? _GEN_8084 : phv_data_399; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_400 = phv_is_valid_processor ? _GEN_8091 : phv_data_400; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_401 = phv_is_valid_processor ? _GEN_8090 : phv_data_401; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_402 = phv_is_valid_processor ? _GEN_8089 : phv_data_402; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_403 = phv_is_valid_processor ? _GEN_8088 : phv_data_403; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_404 = phv_is_valid_processor ? _GEN_8095 : phv_data_404; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_405 = phv_is_valid_processor ? _GEN_8094 : phv_data_405; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_406 = phv_is_valid_processor ? _GEN_8093 : phv_data_406; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_407 = phv_is_valid_processor ? _GEN_8092 : phv_data_407; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_408 = phv_is_valid_processor ? _GEN_8099 : phv_data_408; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_409 = phv_is_valid_processor ? _GEN_8098 : phv_data_409; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_410 = phv_is_valid_processor ? _GEN_8097 : phv_data_410; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_411 = phv_is_valid_processor ? _GEN_8096 : phv_data_411; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_412 = phv_is_valid_processor ? _GEN_8103 : phv_data_412; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_413 = phv_is_valid_processor ? _GEN_8102 : phv_data_413; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_414 = phv_is_valid_processor ? _GEN_8101 : phv_data_414; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_415 = phv_is_valid_processor ? _GEN_8100 : phv_data_415; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_416 = phv_is_valid_processor ? _GEN_8107 : phv_data_416; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_417 = phv_is_valid_processor ? _GEN_8106 : phv_data_417; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_418 = phv_is_valid_processor ? _GEN_8105 : phv_data_418; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_419 = phv_is_valid_processor ? _GEN_8104 : phv_data_419; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_420 = phv_is_valid_processor ? _GEN_8111 : phv_data_420; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_421 = phv_is_valid_processor ? _GEN_8110 : phv_data_421; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_422 = phv_is_valid_processor ? _GEN_8109 : phv_data_422; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_423 = phv_is_valid_processor ? _GEN_8108 : phv_data_423; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_424 = phv_is_valid_processor ? _GEN_8115 : phv_data_424; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_425 = phv_is_valid_processor ? _GEN_8114 : phv_data_425; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_426 = phv_is_valid_processor ? _GEN_8113 : phv_data_426; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_427 = phv_is_valid_processor ? _GEN_8112 : phv_data_427; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_428 = phv_is_valid_processor ? _GEN_8119 : phv_data_428; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_429 = phv_is_valid_processor ? _GEN_8118 : phv_data_429; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_430 = phv_is_valid_processor ? _GEN_8117 : phv_data_430; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_431 = phv_is_valid_processor ? _GEN_8116 : phv_data_431; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_432 = phv_is_valid_processor ? _GEN_8123 : phv_data_432; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_433 = phv_is_valid_processor ? _GEN_8122 : phv_data_433; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_434 = phv_is_valid_processor ? _GEN_8121 : phv_data_434; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_435 = phv_is_valid_processor ? _GEN_8120 : phv_data_435; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_436 = phv_is_valid_processor ? _GEN_8127 : phv_data_436; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_437 = phv_is_valid_processor ? _GEN_8126 : phv_data_437; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_438 = phv_is_valid_processor ? _GEN_8125 : phv_data_438; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_439 = phv_is_valid_processor ? _GEN_8124 : phv_data_439; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_440 = phv_is_valid_processor ? _GEN_8131 : phv_data_440; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_441 = phv_is_valid_processor ? _GEN_8130 : phv_data_441; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_442 = phv_is_valid_processor ? _GEN_8129 : phv_data_442; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_443 = phv_is_valid_processor ? _GEN_8128 : phv_data_443; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_444 = phv_is_valid_processor ? _GEN_8135 : phv_data_444; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_445 = phv_is_valid_processor ? _GEN_8134 : phv_data_445; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_446 = phv_is_valid_processor ? _GEN_8133 : phv_data_446; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_447 = phv_is_valid_processor ? _GEN_8132 : phv_data_447; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_448 = phv_is_valid_processor ? _GEN_8139 : phv_data_448; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_449 = phv_is_valid_processor ? _GEN_8138 : phv_data_449; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_450 = phv_is_valid_processor ? _GEN_8137 : phv_data_450; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_451 = phv_is_valid_processor ? _GEN_8136 : phv_data_451; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_452 = phv_is_valid_processor ? _GEN_8143 : phv_data_452; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_453 = phv_is_valid_processor ? _GEN_8142 : phv_data_453; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_454 = phv_is_valid_processor ? _GEN_8141 : phv_data_454; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_455 = phv_is_valid_processor ? _GEN_8140 : phv_data_455; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_456 = phv_is_valid_processor ? _GEN_8147 : phv_data_456; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_457 = phv_is_valid_processor ? _GEN_8146 : phv_data_457; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_458 = phv_is_valid_processor ? _GEN_8145 : phv_data_458; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_459 = phv_is_valid_processor ? _GEN_8144 : phv_data_459; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_460 = phv_is_valid_processor ? _GEN_8151 : phv_data_460; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_461 = phv_is_valid_processor ? _GEN_8150 : phv_data_461; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_462 = phv_is_valid_processor ? _GEN_8149 : phv_data_462; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_463 = phv_is_valid_processor ? _GEN_8148 : phv_data_463; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_464 = phv_is_valid_processor ? _GEN_8155 : phv_data_464; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_465 = phv_is_valid_processor ? _GEN_8154 : phv_data_465; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_466 = phv_is_valid_processor ? _GEN_8153 : phv_data_466; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_467 = phv_is_valid_processor ? _GEN_8152 : phv_data_467; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_468 = phv_is_valid_processor ? _GEN_8159 : phv_data_468; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_469 = phv_is_valid_processor ? _GEN_8158 : phv_data_469; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_470 = phv_is_valid_processor ? _GEN_8157 : phv_data_470; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_471 = phv_is_valid_processor ? _GEN_8156 : phv_data_471; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_472 = phv_is_valid_processor ? _GEN_8163 : phv_data_472; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_473 = phv_is_valid_processor ? _GEN_8162 : phv_data_473; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_474 = phv_is_valid_processor ? _GEN_8161 : phv_data_474; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_475 = phv_is_valid_processor ? _GEN_8160 : phv_data_475; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_476 = phv_is_valid_processor ? _GEN_8167 : phv_data_476; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_477 = phv_is_valid_processor ? _GEN_8166 : phv_data_477; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_478 = phv_is_valid_processor ? _GEN_8165 : phv_data_478; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_479 = phv_is_valid_processor ? _GEN_8164 : phv_data_479; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_480 = phv_is_valid_processor ? _GEN_8171 : phv_data_480; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_481 = phv_is_valid_processor ? _GEN_8170 : phv_data_481; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_482 = phv_is_valid_processor ? _GEN_8169 : phv_data_482; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_483 = phv_is_valid_processor ? _GEN_8168 : phv_data_483; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_484 = phv_is_valid_processor ? _GEN_8175 : phv_data_484; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_485 = phv_is_valid_processor ? _GEN_8174 : phv_data_485; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_486 = phv_is_valid_processor ? _GEN_8173 : phv_data_486; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_487 = phv_is_valid_processor ? _GEN_8172 : phv_data_487; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_488 = phv_is_valid_processor ? _GEN_8179 : phv_data_488; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_489 = phv_is_valid_processor ? _GEN_8178 : phv_data_489; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_490 = phv_is_valid_processor ? _GEN_8177 : phv_data_490; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_491 = phv_is_valid_processor ? _GEN_8176 : phv_data_491; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_492 = phv_is_valid_processor ? _GEN_8183 : phv_data_492; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_493 = phv_is_valid_processor ? _GEN_8182 : phv_data_493; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_494 = phv_is_valid_processor ? _GEN_8181 : phv_data_494; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_495 = phv_is_valid_processor ? _GEN_8180 : phv_data_495; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_496 = phv_is_valid_processor ? _GEN_8187 : phv_data_496; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_497 = phv_is_valid_processor ? _GEN_8186 : phv_data_497; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_498 = phv_is_valid_processor ? _GEN_8185 : phv_data_498; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_499 = phv_is_valid_processor ? _GEN_8184 : phv_data_499; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_500 = phv_is_valid_processor ? _GEN_8191 : phv_data_500; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_501 = phv_is_valid_processor ? _GEN_8190 : phv_data_501; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_502 = phv_is_valid_processor ? _GEN_8189 : phv_data_502; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_503 = phv_is_valid_processor ? _GEN_8188 : phv_data_503; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_504 = phv_is_valid_processor ? _GEN_8195 : phv_data_504; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_505 = phv_is_valid_processor ? _GEN_8194 : phv_data_505; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_506 = phv_is_valid_processor ? _GEN_8193 : phv_data_506; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_507 = phv_is_valid_processor ? _GEN_8192 : phv_data_507; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_508 = phv_is_valid_processor ? _GEN_8199 : phv_data_508; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_509 = phv_is_valid_processor ? _GEN_8198 : phv_data_509; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_510 = phv_is_valid_processor ? _GEN_8197 : phv_data_510; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_data_511 = phv_is_valid_processor ? _GEN_8196 : phv_data_511; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 450:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 450:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 450:25]
  assign io_pipe_phv_out_next_processor_id = phv_is_valid_processor ? _GEN_7686 : phv_next_processor_id; // @[executor.scala 461:39 executor.scala 450:25]
  assign io_pipe_phv_out_next_config_id = phv_is_valid_processor ? _GEN_7687 : phv_next_config_id; // @[executor.scala 461:39 executor.scala 450:25]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 449:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 449:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 449:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 449:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 449:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 449:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 449:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 449:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 449:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 449:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 449:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 449:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 449:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 449:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 449:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 449:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 449:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 449:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 449:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 449:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 449:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 449:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 449:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 449:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 449:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 449:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 449:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 449:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 449:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 449:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 449:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 449:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 449:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 449:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 449:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 449:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 449:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 449:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 449:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 449:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 449:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 449:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 449:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 449:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 449:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 449:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 449:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 449:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 449:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 449:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 449:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 449:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 449:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 449:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 449:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 449:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 449:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 449:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 449:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 449:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 449:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 449:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 449:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 449:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 449:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 449:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 449:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 449:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 449:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 449:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 449:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 449:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 449:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 449:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 449:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 449:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 449:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 449:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 449:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 449:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 449:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 449:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 449:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 449:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 449:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 449:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 449:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 449:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 449:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 449:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 449:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 449:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 449:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 449:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 449:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 449:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor.scala 449:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor.scala 449:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor.scala 449:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor.scala 449:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor.scala 449:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor.scala 449:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor.scala 449:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor.scala 449:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor.scala 449:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor.scala 449:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor.scala 449:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor.scala 449:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor.scala 449:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor.scala 449:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor.scala 449:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor.scala 449:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor.scala 449:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor.scala 449:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor.scala 449:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor.scala 449:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor.scala 449:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor.scala 449:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor.scala 449:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor.scala 449:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor.scala 449:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor.scala 449:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor.scala 449:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor.scala 449:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor.scala 449:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor.scala 449:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor.scala 449:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor.scala 449:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor.scala 449:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor.scala 449:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor.scala 449:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor.scala 449:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor.scala 449:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor.scala 449:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor.scala 449:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor.scala 449:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor.scala 449:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor.scala 449:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor.scala 449:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor.scala 449:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor.scala 449:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor.scala 449:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor.scala 449:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor.scala 449:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor.scala 449:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor.scala 449:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor.scala 449:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor.scala 449:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor.scala 449:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor.scala 449:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor.scala 449:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor.scala 449:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor.scala 449:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor.scala 449:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor.scala 449:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor.scala 449:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor.scala 449:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor.scala 449:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor.scala 449:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor.scala 449:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor.scala 449:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor.scala 449:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor.scala 449:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor.scala 449:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor.scala 449:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor.scala 449:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor.scala 449:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor.scala 449:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor.scala 449:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor.scala 449:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor.scala 449:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor.scala 449:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor.scala 449:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor.scala 449:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor.scala 449:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor.scala 449:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor.scala 449:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor.scala 449:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor.scala 449:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor.scala 449:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor.scala 449:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor.scala 449:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor.scala 449:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor.scala 449:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor.scala 449:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor.scala 449:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor.scala 449:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor.scala 449:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor.scala 449:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor.scala 449:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor.scala 449:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor.scala 449:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor.scala 449:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor.scala 449:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor.scala 449:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor.scala 449:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor.scala 449:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor.scala 449:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor.scala 449:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor.scala 449:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor.scala 449:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor.scala 449:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor.scala 449:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor.scala 449:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor.scala 449:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor.scala 449:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor.scala 449:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor.scala 449:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor.scala 449:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor.scala 449:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor.scala 449:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor.scala 449:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor.scala 449:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor.scala 449:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor.scala 449:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor.scala 449:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor.scala 449:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor.scala 449:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor.scala 449:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor.scala 449:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor.scala 449:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor.scala 449:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor.scala 449:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor.scala 449:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor.scala 449:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor.scala 449:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor.scala 449:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor.scala 449:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor.scala 449:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor.scala 449:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor.scala 449:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor.scala 449:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor.scala 449:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor.scala 449:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor.scala 449:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor.scala 449:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor.scala 449:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor.scala 449:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor.scala 449:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor.scala 449:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor.scala 449:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor.scala 449:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor.scala 449:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor.scala 449:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor.scala 449:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor.scala 449:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor.scala 449:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor.scala 449:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor.scala 449:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor.scala 449:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor.scala 449:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor.scala 449:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor.scala 449:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor.scala 449:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor.scala 449:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor.scala 449:13]
    phv_data_256 <= io_pipe_phv_in_data_256; // @[executor.scala 449:13]
    phv_data_257 <= io_pipe_phv_in_data_257; // @[executor.scala 449:13]
    phv_data_258 <= io_pipe_phv_in_data_258; // @[executor.scala 449:13]
    phv_data_259 <= io_pipe_phv_in_data_259; // @[executor.scala 449:13]
    phv_data_260 <= io_pipe_phv_in_data_260; // @[executor.scala 449:13]
    phv_data_261 <= io_pipe_phv_in_data_261; // @[executor.scala 449:13]
    phv_data_262 <= io_pipe_phv_in_data_262; // @[executor.scala 449:13]
    phv_data_263 <= io_pipe_phv_in_data_263; // @[executor.scala 449:13]
    phv_data_264 <= io_pipe_phv_in_data_264; // @[executor.scala 449:13]
    phv_data_265 <= io_pipe_phv_in_data_265; // @[executor.scala 449:13]
    phv_data_266 <= io_pipe_phv_in_data_266; // @[executor.scala 449:13]
    phv_data_267 <= io_pipe_phv_in_data_267; // @[executor.scala 449:13]
    phv_data_268 <= io_pipe_phv_in_data_268; // @[executor.scala 449:13]
    phv_data_269 <= io_pipe_phv_in_data_269; // @[executor.scala 449:13]
    phv_data_270 <= io_pipe_phv_in_data_270; // @[executor.scala 449:13]
    phv_data_271 <= io_pipe_phv_in_data_271; // @[executor.scala 449:13]
    phv_data_272 <= io_pipe_phv_in_data_272; // @[executor.scala 449:13]
    phv_data_273 <= io_pipe_phv_in_data_273; // @[executor.scala 449:13]
    phv_data_274 <= io_pipe_phv_in_data_274; // @[executor.scala 449:13]
    phv_data_275 <= io_pipe_phv_in_data_275; // @[executor.scala 449:13]
    phv_data_276 <= io_pipe_phv_in_data_276; // @[executor.scala 449:13]
    phv_data_277 <= io_pipe_phv_in_data_277; // @[executor.scala 449:13]
    phv_data_278 <= io_pipe_phv_in_data_278; // @[executor.scala 449:13]
    phv_data_279 <= io_pipe_phv_in_data_279; // @[executor.scala 449:13]
    phv_data_280 <= io_pipe_phv_in_data_280; // @[executor.scala 449:13]
    phv_data_281 <= io_pipe_phv_in_data_281; // @[executor.scala 449:13]
    phv_data_282 <= io_pipe_phv_in_data_282; // @[executor.scala 449:13]
    phv_data_283 <= io_pipe_phv_in_data_283; // @[executor.scala 449:13]
    phv_data_284 <= io_pipe_phv_in_data_284; // @[executor.scala 449:13]
    phv_data_285 <= io_pipe_phv_in_data_285; // @[executor.scala 449:13]
    phv_data_286 <= io_pipe_phv_in_data_286; // @[executor.scala 449:13]
    phv_data_287 <= io_pipe_phv_in_data_287; // @[executor.scala 449:13]
    phv_data_288 <= io_pipe_phv_in_data_288; // @[executor.scala 449:13]
    phv_data_289 <= io_pipe_phv_in_data_289; // @[executor.scala 449:13]
    phv_data_290 <= io_pipe_phv_in_data_290; // @[executor.scala 449:13]
    phv_data_291 <= io_pipe_phv_in_data_291; // @[executor.scala 449:13]
    phv_data_292 <= io_pipe_phv_in_data_292; // @[executor.scala 449:13]
    phv_data_293 <= io_pipe_phv_in_data_293; // @[executor.scala 449:13]
    phv_data_294 <= io_pipe_phv_in_data_294; // @[executor.scala 449:13]
    phv_data_295 <= io_pipe_phv_in_data_295; // @[executor.scala 449:13]
    phv_data_296 <= io_pipe_phv_in_data_296; // @[executor.scala 449:13]
    phv_data_297 <= io_pipe_phv_in_data_297; // @[executor.scala 449:13]
    phv_data_298 <= io_pipe_phv_in_data_298; // @[executor.scala 449:13]
    phv_data_299 <= io_pipe_phv_in_data_299; // @[executor.scala 449:13]
    phv_data_300 <= io_pipe_phv_in_data_300; // @[executor.scala 449:13]
    phv_data_301 <= io_pipe_phv_in_data_301; // @[executor.scala 449:13]
    phv_data_302 <= io_pipe_phv_in_data_302; // @[executor.scala 449:13]
    phv_data_303 <= io_pipe_phv_in_data_303; // @[executor.scala 449:13]
    phv_data_304 <= io_pipe_phv_in_data_304; // @[executor.scala 449:13]
    phv_data_305 <= io_pipe_phv_in_data_305; // @[executor.scala 449:13]
    phv_data_306 <= io_pipe_phv_in_data_306; // @[executor.scala 449:13]
    phv_data_307 <= io_pipe_phv_in_data_307; // @[executor.scala 449:13]
    phv_data_308 <= io_pipe_phv_in_data_308; // @[executor.scala 449:13]
    phv_data_309 <= io_pipe_phv_in_data_309; // @[executor.scala 449:13]
    phv_data_310 <= io_pipe_phv_in_data_310; // @[executor.scala 449:13]
    phv_data_311 <= io_pipe_phv_in_data_311; // @[executor.scala 449:13]
    phv_data_312 <= io_pipe_phv_in_data_312; // @[executor.scala 449:13]
    phv_data_313 <= io_pipe_phv_in_data_313; // @[executor.scala 449:13]
    phv_data_314 <= io_pipe_phv_in_data_314; // @[executor.scala 449:13]
    phv_data_315 <= io_pipe_phv_in_data_315; // @[executor.scala 449:13]
    phv_data_316 <= io_pipe_phv_in_data_316; // @[executor.scala 449:13]
    phv_data_317 <= io_pipe_phv_in_data_317; // @[executor.scala 449:13]
    phv_data_318 <= io_pipe_phv_in_data_318; // @[executor.scala 449:13]
    phv_data_319 <= io_pipe_phv_in_data_319; // @[executor.scala 449:13]
    phv_data_320 <= io_pipe_phv_in_data_320; // @[executor.scala 449:13]
    phv_data_321 <= io_pipe_phv_in_data_321; // @[executor.scala 449:13]
    phv_data_322 <= io_pipe_phv_in_data_322; // @[executor.scala 449:13]
    phv_data_323 <= io_pipe_phv_in_data_323; // @[executor.scala 449:13]
    phv_data_324 <= io_pipe_phv_in_data_324; // @[executor.scala 449:13]
    phv_data_325 <= io_pipe_phv_in_data_325; // @[executor.scala 449:13]
    phv_data_326 <= io_pipe_phv_in_data_326; // @[executor.scala 449:13]
    phv_data_327 <= io_pipe_phv_in_data_327; // @[executor.scala 449:13]
    phv_data_328 <= io_pipe_phv_in_data_328; // @[executor.scala 449:13]
    phv_data_329 <= io_pipe_phv_in_data_329; // @[executor.scala 449:13]
    phv_data_330 <= io_pipe_phv_in_data_330; // @[executor.scala 449:13]
    phv_data_331 <= io_pipe_phv_in_data_331; // @[executor.scala 449:13]
    phv_data_332 <= io_pipe_phv_in_data_332; // @[executor.scala 449:13]
    phv_data_333 <= io_pipe_phv_in_data_333; // @[executor.scala 449:13]
    phv_data_334 <= io_pipe_phv_in_data_334; // @[executor.scala 449:13]
    phv_data_335 <= io_pipe_phv_in_data_335; // @[executor.scala 449:13]
    phv_data_336 <= io_pipe_phv_in_data_336; // @[executor.scala 449:13]
    phv_data_337 <= io_pipe_phv_in_data_337; // @[executor.scala 449:13]
    phv_data_338 <= io_pipe_phv_in_data_338; // @[executor.scala 449:13]
    phv_data_339 <= io_pipe_phv_in_data_339; // @[executor.scala 449:13]
    phv_data_340 <= io_pipe_phv_in_data_340; // @[executor.scala 449:13]
    phv_data_341 <= io_pipe_phv_in_data_341; // @[executor.scala 449:13]
    phv_data_342 <= io_pipe_phv_in_data_342; // @[executor.scala 449:13]
    phv_data_343 <= io_pipe_phv_in_data_343; // @[executor.scala 449:13]
    phv_data_344 <= io_pipe_phv_in_data_344; // @[executor.scala 449:13]
    phv_data_345 <= io_pipe_phv_in_data_345; // @[executor.scala 449:13]
    phv_data_346 <= io_pipe_phv_in_data_346; // @[executor.scala 449:13]
    phv_data_347 <= io_pipe_phv_in_data_347; // @[executor.scala 449:13]
    phv_data_348 <= io_pipe_phv_in_data_348; // @[executor.scala 449:13]
    phv_data_349 <= io_pipe_phv_in_data_349; // @[executor.scala 449:13]
    phv_data_350 <= io_pipe_phv_in_data_350; // @[executor.scala 449:13]
    phv_data_351 <= io_pipe_phv_in_data_351; // @[executor.scala 449:13]
    phv_data_352 <= io_pipe_phv_in_data_352; // @[executor.scala 449:13]
    phv_data_353 <= io_pipe_phv_in_data_353; // @[executor.scala 449:13]
    phv_data_354 <= io_pipe_phv_in_data_354; // @[executor.scala 449:13]
    phv_data_355 <= io_pipe_phv_in_data_355; // @[executor.scala 449:13]
    phv_data_356 <= io_pipe_phv_in_data_356; // @[executor.scala 449:13]
    phv_data_357 <= io_pipe_phv_in_data_357; // @[executor.scala 449:13]
    phv_data_358 <= io_pipe_phv_in_data_358; // @[executor.scala 449:13]
    phv_data_359 <= io_pipe_phv_in_data_359; // @[executor.scala 449:13]
    phv_data_360 <= io_pipe_phv_in_data_360; // @[executor.scala 449:13]
    phv_data_361 <= io_pipe_phv_in_data_361; // @[executor.scala 449:13]
    phv_data_362 <= io_pipe_phv_in_data_362; // @[executor.scala 449:13]
    phv_data_363 <= io_pipe_phv_in_data_363; // @[executor.scala 449:13]
    phv_data_364 <= io_pipe_phv_in_data_364; // @[executor.scala 449:13]
    phv_data_365 <= io_pipe_phv_in_data_365; // @[executor.scala 449:13]
    phv_data_366 <= io_pipe_phv_in_data_366; // @[executor.scala 449:13]
    phv_data_367 <= io_pipe_phv_in_data_367; // @[executor.scala 449:13]
    phv_data_368 <= io_pipe_phv_in_data_368; // @[executor.scala 449:13]
    phv_data_369 <= io_pipe_phv_in_data_369; // @[executor.scala 449:13]
    phv_data_370 <= io_pipe_phv_in_data_370; // @[executor.scala 449:13]
    phv_data_371 <= io_pipe_phv_in_data_371; // @[executor.scala 449:13]
    phv_data_372 <= io_pipe_phv_in_data_372; // @[executor.scala 449:13]
    phv_data_373 <= io_pipe_phv_in_data_373; // @[executor.scala 449:13]
    phv_data_374 <= io_pipe_phv_in_data_374; // @[executor.scala 449:13]
    phv_data_375 <= io_pipe_phv_in_data_375; // @[executor.scala 449:13]
    phv_data_376 <= io_pipe_phv_in_data_376; // @[executor.scala 449:13]
    phv_data_377 <= io_pipe_phv_in_data_377; // @[executor.scala 449:13]
    phv_data_378 <= io_pipe_phv_in_data_378; // @[executor.scala 449:13]
    phv_data_379 <= io_pipe_phv_in_data_379; // @[executor.scala 449:13]
    phv_data_380 <= io_pipe_phv_in_data_380; // @[executor.scala 449:13]
    phv_data_381 <= io_pipe_phv_in_data_381; // @[executor.scala 449:13]
    phv_data_382 <= io_pipe_phv_in_data_382; // @[executor.scala 449:13]
    phv_data_383 <= io_pipe_phv_in_data_383; // @[executor.scala 449:13]
    phv_data_384 <= io_pipe_phv_in_data_384; // @[executor.scala 449:13]
    phv_data_385 <= io_pipe_phv_in_data_385; // @[executor.scala 449:13]
    phv_data_386 <= io_pipe_phv_in_data_386; // @[executor.scala 449:13]
    phv_data_387 <= io_pipe_phv_in_data_387; // @[executor.scala 449:13]
    phv_data_388 <= io_pipe_phv_in_data_388; // @[executor.scala 449:13]
    phv_data_389 <= io_pipe_phv_in_data_389; // @[executor.scala 449:13]
    phv_data_390 <= io_pipe_phv_in_data_390; // @[executor.scala 449:13]
    phv_data_391 <= io_pipe_phv_in_data_391; // @[executor.scala 449:13]
    phv_data_392 <= io_pipe_phv_in_data_392; // @[executor.scala 449:13]
    phv_data_393 <= io_pipe_phv_in_data_393; // @[executor.scala 449:13]
    phv_data_394 <= io_pipe_phv_in_data_394; // @[executor.scala 449:13]
    phv_data_395 <= io_pipe_phv_in_data_395; // @[executor.scala 449:13]
    phv_data_396 <= io_pipe_phv_in_data_396; // @[executor.scala 449:13]
    phv_data_397 <= io_pipe_phv_in_data_397; // @[executor.scala 449:13]
    phv_data_398 <= io_pipe_phv_in_data_398; // @[executor.scala 449:13]
    phv_data_399 <= io_pipe_phv_in_data_399; // @[executor.scala 449:13]
    phv_data_400 <= io_pipe_phv_in_data_400; // @[executor.scala 449:13]
    phv_data_401 <= io_pipe_phv_in_data_401; // @[executor.scala 449:13]
    phv_data_402 <= io_pipe_phv_in_data_402; // @[executor.scala 449:13]
    phv_data_403 <= io_pipe_phv_in_data_403; // @[executor.scala 449:13]
    phv_data_404 <= io_pipe_phv_in_data_404; // @[executor.scala 449:13]
    phv_data_405 <= io_pipe_phv_in_data_405; // @[executor.scala 449:13]
    phv_data_406 <= io_pipe_phv_in_data_406; // @[executor.scala 449:13]
    phv_data_407 <= io_pipe_phv_in_data_407; // @[executor.scala 449:13]
    phv_data_408 <= io_pipe_phv_in_data_408; // @[executor.scala 449:13]
    phv_data_409 <= io_pipe_phv_in_data_409; // @[executor.scala 449:13]
    phv_data_410 <= io_pipe_phv_in_data_410; // @[executor.scala 449:13]
    phv_data_411 <= io_pipe_phv_in_data_411; // @[executor.scala 449:13]
    phv_data_412 <= io_pipe_phv_in_data_412; // @[executor.scala 449:13]
    phv_data_413 <= io_pipe_phv_in_data_413; // @[executor.scala 449:13]
    phv_data_414 <= io_pipe_phv_in_data_414; // @[executor.scala 449:13]
    phv_data_415 <= io_pipe_phv_in_data_415; // @[executor.scala 449:13]
    phv_data_416 <= io_pipe_phv_in_data_416; // @[executor.scala 449:13]
    phv_data_417 <= io_pipe_phv_in_data_417; // @[executor.scala 449:13]
    phv_data_418 <= io_pipe_phv_in_data_418; // @[executor.scala 449:13]
    phv_data_419 <= io_pipe_phv_in_data_419; // @[executor.scala 449:13]
    phv_data_420 <= io_pipe_phv_in_data_420; // @[executor.scala 449:13]
    phv_data_421 <= io_pipe_phv_in_data_421; // @[executor.scala 449:13]
    phv_data_422 <= io_pipe_phv_in_data_422; // @[executor.scala 449:13]
    phv_data_423 <= io_pipe_phv_in_data_423; // @[executor.scala 449:13]
    phv_data_424 <= io_pipe_phv_in_data_424; // @[executor.scala 449:13]
    phv_data_425 <= io_pipe_phv_in_data_425; // @[executor.scala 449:13]
    phv_data_426 <= io_pipe_phv_in_data_426; // @[executor.scala 449:13]
    phv_data_427 <= io_pipe_phv_in_data_427; // @[executor.scala 449:13]
    phv_data_428 <= io_pipe_phv_in_data_428; // @[executor.scala 449:13]
    phv_data_429 <= io_pipe_phv_in_data_429; // @[executor.scala 449:13]
    phv_data_430 <= io_pipe_phv_in_data_430; // @[executor.scala 449:13]
    phv_data_431 <= io_pipe_phv_in_data_431; // @[executor.scala 449:13]
    phv_data_432 <= io_pipe_phv_in_data_432; // @[executor.scala 449:13]
    phv_data_433 <= io_pipe_phv_in_data_433; // @[executor.scala 449:13]
    phv_data_434 <= io_pipe_phv_in_data_434; // @[executor.scala 449:13]
    phv_data_435 <= io_pipe_phv_in_data_435; // @[executor.scala 449:13]
    phv_data_436 <= io_pipe_phv_in_data_436; // @[executor.scala 449:13]
    phv_data_437 <= io_pipe_phv_in_data_437; // @[executor.scala 449:13]
    phv_data_438 <= io_pipe_phv_in_data_438; // @[executor.scala 449:13]
    phv_data_439 <= io_pipe_phv_in_data_439; // @[executor.scala 449:13]
    phv_data_440 <= io_pipe_phv_in_data_440; // @[executor.scala 449:13]
    phv_data_441 <= io_pipe_phv_in_data_441; // @[executor.scala 449:13]
    phv_data_442 <= io_pipe_phv_in_data_442; // @[executor.scala 449:13]
    phv_data_443 <= io_pipe_phv_in_data_443; // @[executor.scala 449:13]
    phv_data_444 <= io_pipe_phv_in_data_444; // @[executor.scala 449:13]
    phv_data_445 <= io_pipe_phv_in_data_445; // @[executor.scala 449:13]
    phv_data_446 <= io_pipe_phv_in_data_446; // @[executor.scala 449:13]
    phv_data_447 <= io_pipe_phv_in_data_447; // @[executor.scala 449:13]
    phv_data_448 <= io_pipe_phv_in_data_448; // @[executor.scala 449:13]
    phv_data_449 <= io_pipe_phv_in_data_449; // @[executor.scala 449:13]
    phv_data_450 <= io_pipe_phv_in_data_450; // @[executor.scala 449:13]
    phv_data_451 <= io_pipe_phv_in_data_451; // @[executor.scala 449:13]
    phv_data_452 <= io_pipe_phv_in_data_452; // @[executor.scala 449:13]
    phv_data_453 <= io_pipe_phv_in_data_453; // @[executor.scala 449:13]
    phv_data_454 <= io_pipe_phv_in_data_454; // @[executor.scala 449:13]
    phv_data_455 <= io_pipe_phv_in_data_455; // @[executor.scala 449:13]
    phv_data_456 <= io_pipe_phv_in_data_456; // @[executor.scala 449:13]
    phv_data_457 <= io_pipe_phv_in_data_457; // @[executor.scala 449:13]
    phv_data_458 <= io_pipe_phv_in_data_458; // @[executor.scala 449:13]
    phv_data_459 <= io_pipe_phv_in_data_459; // @[executor.scala 449:13]
    phv_data_460 <= io_pipe_phv_in_data_460; // @[executor.scala 449:13]
    phv_data_461 <= io_pipe_phv_in_data_461; // @[executor.scala 449:13]
    phv_data_462 <= io_pipe_phv_in_data_462; // @[executor.scala 449:13]
    phv_data_463 <= io_pipe_phv_in_data_463; // @[executor.scala 449:13]
    phv_data_464 <= io_pipe_phv_in_data_464; // @[executor.scala 449:13]
    phv_data_465 <= io_pipe_phv_in_data_465; // @[executor.scala 449:13]
    phv_data_466 <= io_pipe_phv_in_data_466; // @[executor.scala 449:13]
    phv_data_467 <= io_pipe_phv_in_data_467; // @[executor.scala 449:13]
    phv_data_468 <= io_pipe_phv_in_data_468; // @[executor.scala 449:13]
    phv_data_469 <= io_pipe_phv_in_data_469; // @[executor.scala 449:13]
    phv_data_470 <= io_pipe_phv_in_data_470; // @[executor.scala 449:13]
    phv_data_471 <= io_pipe_phv_in_data_471; // @[executor.scala 449:13]
    phv_data_472 <= io_pipe_phv_in_data_472; // @[executor.scala 449:13]
    phv_data_473 <= io_pipe_phv_in_data_473; // @[executor.scala 449:13]
    phv_data_474 <= io_pipe_phv_in_data_474; // @[executor.scala 449:13]
    phv_data_475 <= io_pipe_phv_in_data_475; // @[executor.scala 449:13]
    phv_data_476 <= io_pipe_phv_in_data_476; // @[executor.scala 449:13]
    phv_data_477 <= io_pipe_phv_in_data_477; // @[executor.scala 449:13]
    phv_data_478 <= io_pipe_phv_in_data_478; // @[executor.scala 449:13]
    phv_data_479 <= io_pipe_phv_in_data_479; // @[executor.scala 449:13]
    phv_data_480 <= io_pipe_phv_in_data_480; // @[executor.scala 449:13]
    phv_data_481 <= io_pipe_phv_in_data_481; // @[executor.scala 449:13]
    phv_data_482 <= io_pipe_phv_in_data_482; // @[executor.scala 449:13]
    phv_data_483 <= io_pipe_phv_in_data_483; // @[executor.scala 449:13]
    phv_data_484 <= io_pipe_phv_in_data_484; // @[executor.scala 449:13]
    phv_data_485 <= io_pipe_phv_in_data_485; // @[executor.scala 449:13]
    phv_data_486 <= io_pipe_phv_in_data_486; // @[executor.scala 449:13]
    phv_data_487 <= io_pipe_phv_in_data_487; // @[executor.scala 449:13]
    phv_data_488 <= io_pipe_phv_in_data_488; // @[executor.scala 449:13]
    phv_data_489 <= io_pipe_phv_in_data_489; // @[executor.scala 449:13]
    phv_data_490 <= io_pipe_phv_in_data_490; // @[executor.scala 449:13]
    phv_data_491 <= io_pipe_phv_in_data_491; // @[executor.scala 449:13]
    phv_data_492 <= io_pipe_phv_in_data_492; // @[executor.scala 449:13]
    phv_data_493 <= io_pipe_phv_in_data_493; // @[executor.scala 449:13]
    phv_data_494 <= io_pipe_phv_in_data_494; // @[executor.scala 449:13]
    phv_data_495 <= io_pipe_phv_in_data_495; // @[executor.scala 449:13]
    phv_data_496 <= io_pipe_phv_in_data_496; // @[executor.scala 449:13]
    phv_data_497 <= io_pipe_phv_in_data_497; // @[executor.scala 449:13]
    phv_data_498 <= io_pipe_phv_in_data_498; // @[executor.scala 449:13]
    phv_data_499 <= io_pipe_phv_in_data_499; // @[executor.scala 449:13]
    phv_data_500 <= io_pipe_phv_in_data_500; // @[executor.scala 449:13]
    phv_data_501 <= io_pipe_phv_in_data_501; // @[executor.scala 449:13]
    phv_data_502 <= io_pipe_phv_in_data_502; // @[executor.scala 449:13]
    phv_data_503 <= io_pipe_phv_in_data_503; // @[executor.scala 449:13]
    phv_data_504 <= io_pipe_phv_in_data_504; // @[executor.scala 449:13]
    phv_data_505 <= io_pipe_phv_in_data_505; // @[executor.scala 449:13]
    phv_data_506 <= io_pipe_phv_in_data_506; // @[executor.scala 449:13]
    phv_data_507 <= io_pipe_phv_in_data_507; // @[executor.scala 449:13]
    phv_data_508 <= io_pipe_phv_in_data_508; // @[executor.scala 449:13]
    phv_data_509 <= io_pipe_phv_in_data_509; // @[executor.scala 449:13]
    phv_data_510 <= io_pipe_phv_in_data_510; // @[executor.scala 449:13]
    phv_data_511 <= io_pipe_phv_in_data_511; // @[executor.scala 449:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 449:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 449:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 449:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 449:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 449:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 449:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 449:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 449:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 449:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 449:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 449:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 449:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 449:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 449:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 449:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 449:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 449:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 449:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 449:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 449:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor.scala 449:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 449:13]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 453:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 453:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 453:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 453:14]
    field_0 <= io_field_in_0; // @[executor.scala 455:15]
    field_1 <= io_field_in_1; // @[executor.scala 455:15]
    field_2 <= io_field_in_2; // @[executor.scala 455:15]
    field_3 <= io_field_in_3; // @[executor.scala 455:15]
    mask_0 <= io_mask_in_0; // @[executor.scala 457:14]
    mask_1 <= io_mask_in_1; // @[executor.scala 457:14]
    mask_2 <= io_mask_in_2; // @[executor.scala 457:14]
    mask_3 <= io_mask_in_3; // @[executor.scala 457:14]
    dst_offset_0 <= io_dst_offset_in_0; // @[executor.scala 459:20]
    dst_offset_1 <= io_dst_offset_in_1; // @[executor.scala 459:20]
    dst_offset_2 <= io_dst_offset_in_2; // @[executor.scala 459:20]
    dst_offset_3 <= io_dst_offset_in_3; // @[executor.scala 459:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_data_256 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  phv_data_257 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  phv_data_258 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  phv_data_259 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  phv_data_260 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  phv_data_261 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  phv_data_262 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  phv_data_263 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  phv_data_264 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  phv_data_265 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  phv_data_266 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  phv_data_267 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  phv_data_268 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  phv_data_269 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  phv_data_270 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  phv_data_271 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  phv_data_272 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_data_273 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_data_274 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  phv_data_275 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  phv_data_276 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  phv_data_277 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  phv_data_278 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  phv_data_279 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  phv_data_280 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  phv_data_281 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  phv_data_282 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  phv_data_283 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  phv_data_284 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  phv_data_285 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  phv_data_286 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  phv_data_287 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  phv_data_288 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  phv_data_289 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  phv_data_290 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  phv_data_291 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  phv_data_292 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  phv_data_293 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  phv_data_294 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  phv_data_295 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  phv_data_296 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  phv_data_297 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  phv_data_298 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  phv_data_299 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  phv_data_300 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  phv_data_301 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  phv_data_302 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  phv_data_303 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  phv_data_304 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  phv_data_305 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  phv_data_306 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  phv_data_307 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  phv_data_308 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  phv_data_309 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  phv_data_310 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  phv_data_311 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  phv_data_312 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  phv_data_313 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  phv_data_314 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  phv_data_315 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  phv_data_316 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  phv_data_317 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  phv_data_318 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  phv_data_319 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  phv_data_320 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  phv_data_321 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  phv_data_322 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  phv_data_323 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  phv_data_324 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  phv_data_325 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  phv_data_326 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  phv_data_327 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  phv_data_328 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  phv_data_329 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  phv_data_330 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  phv_data_331 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  phv_data_332 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  phv_data_333 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  phv_data_334 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  phv_data_335 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  phv_data_336 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  phv_data_337 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  phv_data_338 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  phv_data_339 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  phv_data_340 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  phv_data_341 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  phv_data_342 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  phv_data_343 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  phv_data_344 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  phv_data_345 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  phv_data_346 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  phv_data_347 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  phv_data_348 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  phv_data_349 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  phv_data_350 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  phv_data_351 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  phv_data_352 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  phv_data_353 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  phv_data_354 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  phv_data_355 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  phv_data_356 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  phv_data_357 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  phv_data_358 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  phv_data_359 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  phv_data_360 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  phv_data_361 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  phv_data_362 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  phv_data_363 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  phv_data_364 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  phv_data_365 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  phv_data_366 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  phv_data_367 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  phv_data_368 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  phv_data_369 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  phv_data_370 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  phv_data_371 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  phv_data_372 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  phv_data_373 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  phv_data_374 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  phv_data_375 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  phv_data_376 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  phv_data_377 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  phv_data_378 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  phv_data_379 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  phv_data_380 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  phv_data_381 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  phv_data_382 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  phv_data_383 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  phv_data_384 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  phv_data_385 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  phv_data_386 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  phv_data_387 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  phv_data_388 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  phv_data_389 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  phv_data_390 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  phv_data_391 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  phv_data_392 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  phv_data_393 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  phv_data_394 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  phv_data_395 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  phv_data_396 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  phv_data_397 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  phv_data_398 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  phv_data_399 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  phv_data_400 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  phv_data_401 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  phv_data_402 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  phv_data_403 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  phv_data_404 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  phv_data_405 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  phv_data_406 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  phv_data_407 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  phv_data_408 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  phv_data_409 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  phv_data_410 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  phv_data_411 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  phv_data_412 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  phv_data_413 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  phv_data_414 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  phv_data_415 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  phv_data_416 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  phv_data_417 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  phv_data_418 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  phv_data_419 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  phv_data_420 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  phv_data_421 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  phv_data_422 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  phv_data_423 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  phv_data_424 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  phv_data_425 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  phv_data_426 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  phv_data_427 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  phv_data_428 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  phv_data_429 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  phv_data_430 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  phv_data_431 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  phv_data_432 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  phv_data_433 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  phv_data_434 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  phv_data_435 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  phv_data_436 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  phv_data_437 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  phv_data_438 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  phv_data_439 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  phv_data_440 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  phv_data_441 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  phv_data_442 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  phv_data_443 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  phv_data_444 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  phv_data_445 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  phv_data_446 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  phv_data_447 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  phv_data_448 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  phv_data_449 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  phv_data_450 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  phv_data_451 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  phv_data_452 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  phv_data_453 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  phv_data_454 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  phv_data_455 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  phv_data_456 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  phv_data_457 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  phv_data_458 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  phv_data_459 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  phv_data_460 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  phv_data_461 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  phv_data_462 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  phv_data_463 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  phv_data_464 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  phv_data_465 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  phv_data_466 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  phv_data_467 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  phv_data_468 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  phv_data_469 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  phv_data_470 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  phv_data_471 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  phv_data_472 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  phv_data_473 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  phv_data_474 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  phv_data_475 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  phv_data_476 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  phv_data_477 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  phv_data_478 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  phv_data_479 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  phv_data_480 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  phv_data_481 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  phv_data_482 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  phv_data_483 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  phv_data_484 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  phv_data_485 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  phv_data_486 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  phv_data_487 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  phv_data_488 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  phv_data_489 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  phv_data_490 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  phv_data_491 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  phv_data_492 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  phv_data_493 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  phv_data_494 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  phv_data_495 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  phv_data_496 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  phv_data_497 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  phv_data_498 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  phv_data_499 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  phv_data_500 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  phv_data_501 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  phv_data_502 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  phv_data_503 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  phv_data_504 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  phv_data_505 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  phv_data_506 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  phv_data_507 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  phv_data_508 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  phv_data_509 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  phv_data_510 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  phv_data_511 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  phv_header_0 = _RAND_512[15:0];
  _RAND_513 = {1{`RANDOM}};
  phv_header_1 = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  phv_header_2 = _RAND_514[15:0];
  _RAND_515 = {1{`RANDOM}};
  phv_header_3 = _RAND_515[15:0];
  _RAND_516 = {1{`RANDOM}};
  phv_header_4 = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  phv_header_5 = _RAND_517[15:0];
  _RAND_518 = {1{`RANDOM}};
  phv_header_6 = _RAND_518[15:0];
  _RAND_519 = {1{`RANDOM}};
  phv_header_7 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  phv_header_8 = _RAND_520[15:0];
  _RAND_521 = {1{`RANDOM}};
  phv_header_9 = _RAND_521[15:0];
  _RAND_522 = {1{`RANDOM}};
  phv_header_10 = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  phv_header_11 = _RAND_523[15:0];
  _RAND_524 = {1{`RANDOM}};
  phv_header_12 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  phv_header_13 = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  phv_header_14 = _RAND_526[15:0];
  _RAND_527 = {1{`RANDOM}};
  phv_header_15 = _RAND_527[15:0];
  _RAND_528 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_530[15:0];
  _RAND_531 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  phv_next_config_id = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  vliw_0 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  vliw_1 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  vliw_2 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  vliw_3 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  field_0 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  field_1 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  field_2 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  field_3 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  mask_0 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  mask_1 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  mask_2 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  mask_3 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  dst_offset_0 = _RAND_546[5:0];
  _RAND_547 = {1{`RANDOM}};
  dst_offset_1 = _RAND_547[5:0];
  _RAND_548 = {1{`RANDOM}};
  dst_offset_2 = _RAND_548[5:0];
  _RAND_549 = {1{`RANDOM}};
  dst_offset_3 = _RAND_549[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
