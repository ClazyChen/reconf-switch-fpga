module InPort(
  input        clock,
  input        reset,
  output [7:0] io_phv_out_data_0,
  output [7:0] io_phv_out_data_1,
  output [7:0] io_phv_out_data_2,
  output [7:0] io_phv_out_data_3,
  output [7:0] io_phv_out_data_4,
  output [7:0] io_phv_out_data_5,
  output [7:0] io_phv_out_data_6,
  output [7:0] io_phv_out_data_7,
  output [7:0] io_phv_out_data_8,
  output [7:0] io_phv_out_data_9,
  output [7:0] io_phv_out_data_10,
  output [7:0] io_phv_out_data_11,
  output [7:0] io_phv_out_data_12,
  output [7:0] io_phv_out_data_13,
  output [7:0] io_phv_out_data_14,
  output [7:0] io_phv_out_data_15,
  output [7:0] io_phv_out_data_16,
  output [7:0] io_phv_out_data_17,
  output [7:0] io_phv_out_data_18,
  output [7:0] io_phv_out_data_19,
  output [7:0] io_phv_out_data_20,
  output [7:0] io_phv_out_data_21,
  output [7:0] io_phv_out_data_22,
  output [7:0] io_phv_out_data_23,
  output [7:0] io_phv_out_data_24,
  output [7:0] io_phv_out_data_25,
  output [7:0] io_phv_out_data_26,
  output [7:0] io_phv_out_data_27,
  output [7:0] io_phv_out_data_28,
  output [7:0] io_phv_out_data_29,
  output [7:0] io_phv_out_data_30,
  output [7:0] io_phv_out_data_31,
  output [7:0] io_phv_out_data_32,
  output [7:0] io_phv_out_data_33,
  output [7:0] io_phv_out_data_34,
  output [7:0] io_phv_out_data_35,
  output [7:0] io_phv_out_data_36,
  output [7:0] io_phv_out_data_37,
  output [7:0] io_phv_out_data_38,
  output [7:0] io_phv_out_data_39,
  output [7:0] io_phv_out_data_40,
  output [7:0] io_phv_out_data_41,
  output [7:0] io_phv_out_data_42,
  output [7:0] io_phv_out_data_43,
  output [7:0] io_phv_out_data_44,
  output [7:0] io_phv_out_data_45,
  output [7:0] io_phv_out_data_46,
  output [7:0] io_phv_out_data_47,
  output [7:0] io_phv_out_data_48,
  output [7:0] io_phv_out_data_49,
  output [7:0] io_phv_out_data_50,
  output [7:0] io_phv_out_data_51,
  output [7:0] io_phv_out_data_52,
  output [7:0] io_phv_out_data_53,
  output [7:0] io_phv_out_data_54,
  output [7:0] io_phv_out_data_55,
  output [7:0] io_phv_out_data_56,
  output [7:0] io_phv_out_data_57,
  output [7:0] io_phv_out_data_58,
  output [7:0] io_phv_out_data_59,
  output [7:0] io_phv_out_data_60,
  output [7:0] io_phv_out_data_61,
  output [7:0] io_phv_out_data_62,
  output [7:0] io_phv_out_data_63,
  output [7:0] io_phv_out_data_64,
  output [7:0] io_phv_out_data_65,
  output [7:0] io_phv_out_data_66,
  output [7:0] io_phv_out_data_67,
  output [7:0] io_phv_out_data_68,
  output [7:0] io_phv_out_data_69,
  output [7:0] io_phv_out_data_70,
  output [7:0] io_phv_out_data_71,
  output [7:0] io_phv_out_data_72,
  output [7:0] io_phv_out_data_73,
  output [7:0] io_phv_out_data_74,
  output [7:0] io_phv_out_data_75,
  output [7:0] io_phv_out_data_76,
  output [7:0] io_phv_out_data_77,
  output [7:0] io_phv_out_data_78,
  output [7:0] io_phv_out_data_79,
  output [7:0] io_phv_out_data_80,
  output [7:0] io_phv_out_data_81,
  output [7:0] io_phv_out_data_82,
  output [7:0] io_phv_out_data_83,
  output [7:0] io_phv_out_data_84,
  output [7:0] io_phv_out_data_85,
  output [7:0] io_phv_out_data_86,
  output [7:0] io_phv_out_data_87,
  output [7:0] io_phv_out_data_88,
  output [7:0] io_phv_out_data_89,
  output [7:0] io_phv_out_data_90,
  output [7:0] io_phv_out_data_91,
  output [7:0] io_phv_out_data_92,
  output [7:0] io_phv_out_data_93,
  output [7:0] io_phv_out_data_94,
  output [7:0] io_phv_out_data_95,
  output [7:0] io_phv_out_data_96,
  output [7:0] io_phv_out_data_97,
  output [7:0] io_phv_out_data_98,
  output [7:0] io_phv_out_data_99,
  output [7:0] io_phv_out_data_100,
  output [7:0] io_phv_out_data_101,
  output [7:0] io_phv_out_data_102,
  output [7:0] io_phv_out_data_103,
  output [7:0] io_phv_out_data_104,
  output [7:0] io_phv_out_data_105,
  output [7:0] io_phv_out_data_106,
  output [7:0] io_phv_out_data_107,
  output [7:0] io_phv_out_data_108,
  output [7:0] io_phv_out_data_109,
  output [7:0] io_phv_out_data_110,
  output [7:0] io_phv_out_data_111,
  output [7:0] io_phv_out_data_112,
  output [7:0] io_phv_out_data_113,
  output [7:0] io_phv_out_data_114,
  output [7:0] io_phv_out_data_115,
  output [7:0] io_phv_out_data_116,
  output [7:0] io_phv_out_data_117,
  output [7:0] io_phv_out_data_118,
  output [7:0] io_phv_out_data_119,
  output [7:0] io_phv_out_data_120,
  output [7:0] io_phv_out_data_121,
  output [7:0] io_phv_out_data_122,
  output [7:0] io_phv_out_data_123,
  output [7:0] io_phv_out_data_124,
  output [7:0] io_phv_out_data_125,
  output [7:0] io_phv_out_data_126,
  output [7:0] io_phv_out_data_127,
  output [7:0] io_phv_out_data_128,
  output [7:0] io_phv_out_data_129,
  output [7:0] io_phv_out_data_130,
  output [7:0] io_phv_out_data_131,
  output [7:0] io_phv_out_data_132,
  output [7:0] io_phv_out_data_133,
  output [7:0] io_phv_out_data_134,
  output [7:0] io_phv_out_data_135,
  output [7:0] io_phv_out_data_136,
  output [7:0] io_phv_out_data_137,
  output [7:0] io_phv_out_data_138,
  output [7:0] io_phv_out_data_139,
  output [7:0] io_phv_out_data_140,
  output [7:0] io_phv_out_data_141,
  output [7:0] io_phv_out_data_142,
  output [7:0] io_phv_out_data_143,
  output [7:0] io_phv_out_data_144,
  output [7:0] io_phv_out_data_145,
  output [7:0] io_phv_out_data_146,
  output [7:0] io_phv_out_data_147,
  output [7:0] io_phv_out_data_148,
  output [7:0] io_phv_out_data_149,
  output [7:0] io_phv_out_data_150,
  output [7:0] io_phv_out_data_151,
  output [7:0] io_phv_out_data_152,
  output [7:0] io_phv_out_data_153,
  output [7:0] io_phv_out_data_154,
  output [7:0] io_phv_out_data_155,
  output [7:0] io_phv_out_data_156,
  output [7:0] io_phv_out_data_157,
  output [7:0] io_phv_out_data_158,
  output [7:0] io_phv_out_data_159,
  output [7:0] io_phv_out_data_160,
  output [7:0] io_phv_out_data_161,
  output [7:0] io_phv_out_data_162,
  output [7:0] io_phv_out_data_163,
  output [7:0] io_phv_out_data_164,
  output [7:0] io_phv_out_data_165,
  output [7:0] io_phv_out_data_166,
  output [7:0] io_phv_out_data_167,
  output [7:0] io_phv_out_data_168,
  output [7:0] io_phv_out_data_169,
  output [7:0] io_phv_out_data_170,
  output [7:0] io_phv_out_data_171,
  output [7:0] io_phv_out_data_172,
  output [7:0] io_phv_out_data_173,
  output [7:0] io_phv_out_data_174,
  output [7:0] io_phv_out_data_175,
  output [7:0] io_phv_out_data_176,
  output [7:0] io_phv_out_data_177,
  output [7:0] io_phv_out_data_178,
  output [7:0] io_phv_out_data_179,
  output [7:0] io_phv_out_data_180,
  output [7:0] io_phv_out_data_181,
  output [7:0] io_phv_out_data_182,
  output [7:0] io_phv_out_data_183,
  output [7:0] io_phv_out_data_184,
  output [7:0] io_phv_out_data_185,
  output [7:0] io_phv_out_data_186,
  output [7:0] io_phv_out_data_187,
  output [7:0] io_phv_out_data_188,
  output [7:0] io_phv_out_data_189,
  output [7:0] io_phv_out_data_190,
  output [7:0] io_phv_out_data_191,
  output [7:0] io_phv_out_data_192,
  output [7:0] io_phv_out_data_193,
  output [7:0] io_phv_out_data_194,
  output [7:0] io_phv_out_data_195,
  output [7:0] io_phv_out_data_196,
  output [7:0] io_phv_out_data_197,
  output [7:0] io_phv_out_data_198,
  output [7:0] io_phv_out_data_199,
  output [7:0] io_phv_out_data_200,
  output [7:0] io_phv_out_data_201,
  output [7:0] io_phv_out_data_202,
  output [7:0] io_phv_out_data_203,
  output [7:0] io_phv_out_data_204,
  output [7:0] io_phv_out_data_205,
  output [7:0] io_phv_out_data_206,
  output [7:0] io_phv_out_data_207,
  output [7:0] io_phv_out_data_208,
  output [7:0] io_phv_out_data_209,
  output [7:0] io_phv_out_data_210,
  output [7:0] io_phv_out_data_211,
  output [7:0] io_phv_out_data_212,
  output [7:0] io_phv_out_data_213,
  output [7:0] io_phv_out_data_214,
  output [7:0] io_phv_out_data_215,
  output [7:0] io_phv_out_data_216,
  output [7:0] io_phv_out_data_217,
  output [7:0] io_phv_out_data_218,
  output [7:0] io_phv_out_data_219,
  output [7:0] io_phv_out_data_220,
  output [7:0] io_phv_out_data_221,
  output [7:0] io_phv_out_data_222,
  output [7:0] io_phv_out_data_223,
  output [7:0] io_phv_out_data_224,
  output [7:0] io_phv_out_data_225,
  output [7:0] io_phv_out_data_226,
  output [7:0] io_phv_out_data_227,
  output [7:0] io_phv_out_data_228,
  output [7:0] io_phv_out_data_229,
  output [7:0] io_phv_out_data_230,
  output [7:0] io_phv_out_data_231,
  output [7:0] io_phv_out_data_232,
  output [7:0] io_phv_out_data_233,
  output [7:0] io_phv_out_data_234,
  output [7:0] io_phv_out_data_235,
  output [7:0] io_phv_out_data_236,
  output [7:0] io_phv_out_data_237,
  output [7:0] io_phv_out_data_238,
  output [7:0] io_phv_out_data_239,
  output [7:0] io_phv_out_data_240,
  output [7:0] io_phv_out_data_241,
  output [7:0] io_phv_out_data_242,
  output [7:0] io_phv_out_data_243,
  output [7:0] io_phv_out_data_244,
  output [7:0] io_phv_out_data_245,
  output [7:0] io_phv_out_data_246,
  output [7:0] io_phv_out_data_247,
  output [7:0] io_phv_out_data_248,
  output [7:0] io_phv_out_data_249,
  output [7:0] io_phv_out_data_250,
  output [7:0] io_phv_out_data_251,
  output [7:0] io_phv_out_data_252,
  output [7:0] io_phv_out_data_253,
  output [7:0] io_phv_out_data_254,
  output [7:0] io_phv_out_data_255,
  output [7:0] io_phv_out_data_256,
  output [7:0] io_phv_out_data_257,
  output [7:0] io_phv_out_data_258,
  output [7:0] io_phv_out_data_259,
  output [7:0] io_phv_out_data_260,
  output [7:0] io_phv_out_data_261,
  output [7:0] io_phv_out_data_262,
  output [7:0] io_phv_out_data_263,
  output [7:0] io_phv_out_data_264,
  output [7:0] io_phv_out_data_265,
  output [7:0] io_phv_out_data_266,
  output [7:0] io_phv_out_data_267,
  output [7:0] io_phv_out_data_268,
  output [7:0] io_phv_out_data_269,
  output [7:0] io_phv_out_data_270,
  output [7:0] io_phv_out_data_271,
  output [7:0] io_phv_out_data_272,
  output [7:0] io_phv_out_data_273,
  output [7:0] io_phv_out_data_274,
  output [7:0] io_phv_out_data_275,
  output [7:0] io_phv_out_data_276,
  output [7:0] io_phv_out_data_277,
  output [7:0] io_phv_out_data_278,
  output [7:0] io_phv_out_data_279,
  output [7:0] io_phv_out_data_280,
  output [7:0] io_phv_out_data_281,
  output [7:0] io_phv_out_data_282,
  output [7:0] io_phv_out_data_283,
  output [7:0] io_phv_out_data_284,
  output [7:0] io_phv_out_data_285,
  output [7:0] io_phv_out_data_286,
  output [7:0] io_phv_out_data_287,
  output [7:0] io_phv_out_data_288,
  output [7:0] io_phv_out_data_289,
  output [7:0] io_phv_out_data_290,
  output [7:0] io_phv_out_data_291,
  output [7:0] io_phv_out_data_292,
  output [7:0] io_phv_out_data_293,
  output [7:0] io_phv_out_data_294,
  output [7:0] io_phv_out_data_295,
  output [7:0] io_phv_out_data_296,
  output [7:0] io_phv_out_data_297,
  output [7:0] io_phv_out_data_298,
  output [7:0] io_phv_out_data_299,
  output [7:0] io_phv_out_data_300,
  output [7:0] io_phv_out_data_301,
  output [7:0] io_phv_out_data_302,
  output [7:0] io_phv_out_data_303,
  output [7:0] io_phv_out_data_304,
  output [7:0] io_phv_out_data_305,
  output [7:0] io_phv_out_data_306,
  output [7:0] io_phv_out_data_307,
  output [7:0] io_phv_out_data_308,
  output [7:0] io_phv_out_data_309,
  output [7:0] io_phv_out_data_310,
  output [7:0] io_phv_out_data_311,
  output [7:0] io_phv_out_data_312,
  output [7:0] io_phv_out_data_313,
  output [7:0] io_phv_out_data_314,
  output [7:0] io_phv_out_data_315,
  output [7:0] io_phv_out_data_316,
  output [7:0] io_phv_out_data_317,
  output [7:0] io_phv_out_data_318,
  output [7:0] io_phv_out_data_319,
  output [7:0] io_phv_out_data_320,
  output [7:0] io_phv_out_data_321,
  output [7:0] io_phv_out_data_322,
  output [7:0] io_phv_out_data_323,
  output [7:0] io_phv_out_data_324,
  output [7:0] io_phv_out_data_325,
  output [7:0] io_phv_out_data_326,
  output [7:0] io_phv_out_data_327,
  output [7:0] io_phv_out_data_328,
  output [7:0] io_phv_out_data_329,
  output [7:0] io_phv_out_data_330,
  output [7:0] io_phv_out_data_331,
  output [7:0] io_phv_out_data_332,
  output [7:0] io_phv_out_data_333,
  output [7:0] io_phv_out_data_334,
  output [7:0] io_phv_out_data_335,
  output [7:0] io_phv_out_data_336,
  output [7:0] io_phv_out_data_337,
  output [7:0] io_phv_out_data_338,
  output [7:0] io_phv_out_data_339,
  output [7:0] io_phv_out_data_340,
  output [7:0] io_phv_out_data_341,
  output [7:0] io_phv_out_data_342,
  output [7:0] io_phv_out_data_343,
  output [7:0] io_phv_out_data_344,
  output [7:0] io_phv_out_data_345,
  output [7:0] io_phv_out_data_346,
  output [7:0] io_phv_out_data_347,
  output [7:0] io_phv_out_data_348,
  output [7:0] io_phv_out_data_349,
  output [7:0] io_phv_out_data_350,
  output [7:0] io_phv_out_data_351,
  output [7:0] io_phv_out_data_352,
  output [7:0] io_phv_out_data_353,
  output [7:0] io_phv_out_data_354,
  output [7:0] io_phv_out_data_355,
  output [7:0] io_phv_out_data_356,
  output [7:0] io_phv_out_data_357,
  output [7:0] io_phv_out_data_358,
  output [7:0] io_phv_out_data_359,
  output [7:0] io_phv_out_data_360,
  output [7:0] io_phv_out_data_361,
  output [7:0] io_phv_out_data_362,
  output [7:0] io_phv_out_data_363,
  output [7:0] io_phv_out_data_364,
  output [7:0] io_phv_out_data_365,
  output [7:0] io_phv_out_data_366,
  output [7:0] io_phv_out_data_367,
  output [7:0] io_phv_out_data_368,
  output [7:0] io_phv_out_data_369,
  output [7:0] io_phv_out_data_370,
  output [7:0] io_phv_out_data_371,
  output [7:0] io_phv_out_data_372,
  output [7:0] io_phv_out_data_373,
  output [7:0] io_phv_out_data_374,
  output [7:0] io_phv_out_data_375,
  output [7:0] io_phv_out_data_376,
  output [7:0] io_phv_out_data_377,
  output [7:0] io_phv_out_data_378,
  output [7:0] io_phv_out_data_379,
  output [7:0] io_phv_out_data_380,
  output [7:0] io_phv_out_data_381,
  output [7:0] io_phv_out_data_382,
  output [7:0] io_phv_out_data_383
);
  wire  rand_exe_prng_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_1_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_2_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_3_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_4_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_5_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_6_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_7_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_8_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_9_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_10_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_11_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_12_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_13_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_14_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_15_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_16_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_17_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_18_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_19_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_20_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_21_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_22_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_23_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_24_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_25_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_26_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_27_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_28_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_29_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_30_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_31_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_32_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_33_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_34_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_35_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_36_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_37_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_38_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_39_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_40_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_41_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_42_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_43_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_44_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_45_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_46_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_47_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_48_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_49_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_50_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_51_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_52_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_53_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_54_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_55_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_56_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_57_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_58_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_59_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_60_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_61_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_62_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_63_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_64_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_65_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_66_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_67_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_68_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_69_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_70_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_71_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_72_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_73_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_74_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_75_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_76_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_77_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_78_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_79_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_80_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_81_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_82_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_83_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_84_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_85_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_86_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_87_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_88_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_89_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_90_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_91_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_92_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_93_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_94_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_95_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_96_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_97_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_98_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_99_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_100_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_101_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_102_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_103_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_104_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_105_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_106_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_107_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_108_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_109_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_110_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_111_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_112_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_113_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_114_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_115_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_116_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_117_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_118_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_119_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_120_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_121_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_122_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_123_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_124_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_125_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_126_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_127_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_128_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_129_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_130_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_131_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_132_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_133_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_134_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_135_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_136_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_137_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_138_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_139_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_140_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_141_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_142_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_143_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_144_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_145_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_146_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_147_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_148_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_149_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_150_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_151_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_152_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_153_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_154_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_155_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_156_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_157_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_158_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_159_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_160_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_161_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_162_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_163_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_164_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_165_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_166_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_167_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_168_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_169_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_170_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_171_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_172_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_173_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_174_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_175_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_176_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_177_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_178_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_179_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_180_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_181_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_182_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_183_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_184_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_185_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_186_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_187_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_188_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_189_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_190_io_out_15; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_clock; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_reset; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_0; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_1; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_2; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_3; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_4; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_5; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_6; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_7; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_8; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_9; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_10; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_11; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_12; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_13; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_14; // @[PRNG.scala 82:22]
  wire  rand_exe_prng_191_io_out_15; // @[PRNG.scala 82:22]
  wire [7:0] rand_exe_lo = {rand_exe_prng_io_out_7,rand_exe_prng_io_out_6,rand_exe_prng_io_out_5,rand_exe_prng_io_out_4,
    rand_exe_prng_io_out_3,rand_exe_prng_io_out_2,rand_exe_prng_io_out_1,rand_exe_prng_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_0 = {rand_exe_prng_io_out_15,rand_exe_prng_io_out_14,rand_exe_prng_io_out_13,rand_exe_prng_io_out_12,
    rand_exe_prng_io_out_11,rand_exe_prng_io_out_10,rand_exe_prng_io_out_9,rand_exe_prng_io_out_8,rand_exe_lo}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_1 = {rand_exe_prng_1_io_out_7,rand_exe_prng_1_io_out_6,rand_exe_prng_1_io_out_5,
    rand_exe_prng_1_io_out_4,rand_exe_prng_1_io_out_3,rand_exe_prng_1_io_out_2,rand_exe_prng_1_io_out_1,
    rand_exe_prng_1_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_1 = {rand_exe_prng_1_io_out_15,rand_exe_prng_1_io_out_14,rand_exe_prng_1_io_out_13,
    rand_exe_prng_1_io_out_12,rand_exe_prng_1_io_out_11,rand_exe_prng_1_io_out_10,rand_exe_prng_1_io_out_9,
    rand_exe_prng_1_io_out_8,rand_exe_lo_1}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_2 = {rand_exe_prng_2_io_out_7,rand_exe_prng_2_io_out_6,rand_exe_prng_2_io_out_5,
    rand_exe_prng_2_io_out_4,rand_exe_prng_2_io_out_3,rand_exe_prng_2_io_out_2,rand_exe_prng_2_io_out_1,
    rand_exe_prng_2_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_2 = {rand_exe_prng_2_io_out_15,rand_exe_prng_2_io_out_14,rand_exe_prng_2_io_out_13,
    rand_exe_prng_2_io_out_12,rand_exe_prng_2_io_out_11,rand_exe_prng_2_io_out_10,rand_exe_prng_2_io_out_9,
    rand_exe_prng_2_io_out_8,rand_exe_lo_2}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_3 = {rand_exe_prng_3_io_out_7,rand_exe_prng_3_io_out_6,rand_exe_prng_3_io_out_5,
    rand_exe_prng_3_io_out_4,rand_exe_prng_3_io_out_3,rand_exe_prng_3_io_out_2,rand_exe_prng_3_io_out_1,
    rand_exe_prng_3_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_3 = {rand_exe_prng_3_io_out_15,rand_exe_prng_3_io_out_14,rand_exe_prng_3_io_out_13,
    rand_exe_prng_3_io_out_12,rand_exe_prng_3_io_out_11,rand_exe_prng_3_io_out_10,rand_exe_prng_3_io_out_9,
    rand_exe_prng_3_io_out_8,rand_exe_lo_3}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_4 = {rand_exe_prng_4_io_out_7,rand_exe_prng_4_io_out_6,rand_exe_prng_4_io_out_5,
    rand_exe_prng_4_io_out_4,rand_exe_prng_4_io_out_3,rand_exe_prng_4_io_out_2,rand_exe_prng_4_io_out_1,
    rand_exe_prng_4_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_4 = {rand_exe_prng_4_io_out_15,rand_exe_prng_4_io_out_14,rand_exe_prng_4_io_out_13,
    rand_exe_prng_4_io_out_12,rand_exe_prng_4_io_out_11,rand_exe_prng_4_io_out_10,rand_exe_prng_4_io_out_9,
    rand_exe_prng_4_io_out_8,rand_exe_lo_4}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_5 = {rand_exe_prng_5_io_out_7,rand_exe_prng_5_io_out_6,rand_exe_prng_5_io_out_5,
    rand_exe_prng_5_io_out_4,rand_exe_prng_5_io_out_3,rand_exe_prng_5_io_out_2,rand_exe_prng_5_io_out_1,
    rand_exe_prng_5_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_5 = {rand_exe_prng_5_io_out_15,rand_exe_prng_5_io_out_14,rand_exe_prng_5_io_out_13,
    rand_exe_prng_5_io_out_12,rand_exe_prng_5_io_out_11,rand_exe_prng_5_io_out_10,rand_exe_prng_5_io_out_9,
    rand_exe_prng_5_io_out_8,rand_exe_lo_5}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_6 = {rand_exe_prng_6_io_out_7,rand_exe_prng_6_io_out_6,rand_exe_prng_6_io_out_5,
    rand_exe_prng_6_io_out_4,rand_exe_prng_6_io_out_3,rand_exe_prng_6_io_out_2,rand_exe_prng_6_io_out_1,
    rand_exe_prng_6_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_6 = {rand_exe_prng_6_io_out_15,rand_exe_prng_6_io_out_14,rand_exe_prng_6_io_out_13,
    rand_exe_prng_6_io_out_12,rand_exe_prng_6_io_out_11,rand_exe_prng_6_io_out_10,rand_exe_prng_6_io_out_9,
    rand_exe_prng_6_io_out_8,rand_exe_lo_6}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_7 = {rand_exe_prng_7_io_out_7,rand_exe_prng_7_io_out_6,rand_exe_prng_7_io_out_5,
    rand_exe_prng_7_io_out_4,rand_exe_prng_7_io_out_3,rand_exe_prng_7_io_out_2,rand_exe_prng_7_io_out_1,
    rand_exe_prng_7_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_7 = {rand_exe_prng_7_io_out_15,rand_exe_prng_7_io_out_14,rand_exe_prng_7_io_out_13,
    rand_exe_prng_7_io_out_12,rand_exe_prng_7_io_out_11,rand_exe_prng_7_io_out_10,rand_exe_prng_7_io_out_9,
    rand_exe_prng_7_io_out_8,rand_exe_lo_7}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_8 = {rand_exe_prng_8_io_out_7,rand_exe_prng_8_io_out_6,rand_exe_prng_8_io_out_5,
    rand_exe_prng_8_io_out_4,rand_exe_prng_8_io_out_3,rand_exe_prng_8_io_out_2,rand_exe_prng_8_io_out_1,
    rand_exe_prng_8_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_8 = {rand_exe_prng_8_io_out_15,rand_exe_prng_8_io_out_14,rand_exe_prng_8_io_out_13,
    rand_exe_prng_8_io_out_12,rand_exe_prng_8_io_out_11,rand_exe_prng_8_io_out_10,rand_exe_prng_8_io_out_9,
    rand_exe_prng_8_io_out_8,rand_exe_lo_8}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_9 = {rand_exe_prng_9_io_out_7,rand_exe_prng_9_io_out_6,rand_exe_prng_9_io_out_5,
    rand_exe_prng_9_io_out_4,rand_exe_prng_9_io_out_3,rand_exe_prng_9_io_out_2,rand_exe_prng_9_io_out_1,
    rand_exe_prng_9_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_9 = {rand_exe_prng_9_io_out_15,rand_exe_prng_9_io_out_14,rand_exe_prng_9_io_out_13,
    rand_exe_prng_9_io_out_12,rand_exe_prng_9_io_out_11,rand_exe_prng_9_io_out_10,rand_exe_prng_9_io_out_9,
    rand_exe_prng_9_io_out_8,rand_exe_lo_9}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_10 = {rand_exe_prng_10_io_out_7,rand_exe_prng_10_io_out_6,rand_exe_prng_10_io_out_5,
    rand_exe_prng_10_io_out_4,rand_exe_prng_10_io_out_3,rand_exe_prng_10_io_out_2,rand_exe_prng_10_io_out_1,
    rand_exe_prng_10_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_10 = {rand_exe_prng_10_io_out_15,rand_exe_prng_10_io_out_14,rand_exe_prng_10_io_out_13,
    rand_exe_prng_10_io_out_12,rand_exe_prng_10_io_out_11,rand_exe_prng_10_io_out_10,rand_exe_prng_10_io_out_9,
    rand_exe_prng_10_io_out_8,rand_exe_lo_10}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_11 = {rand_exe_prng_11_io_out_7,rand_exe_prng_11_io_out_6,rand_exe_prng_11_io_out_5,
    rand_exe_prng_11_io_out_4,rand_exe_prng_11_io_out_3,rand_exe_prng_11_io_out_2,rand_exe_prng_11_io_out_1,
    rand_exe_prng_11_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_11 = {rand_exe_prng_11_io_out_15,rand_exe_prng_11_io_out_14,rand_exe_prng_11_io_out_13,
    rand_exe_prng_11_io_out_12,rand_exe_prng_11_io_out_11,rand_exe_prng_11_io_out_10,rand_exe_prng_11_io_out_9,
    rand_exe_prng_11_io_out_8,rand_exe_lo_11}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_12 = {rand_exe_prng_12_io_out_7,rand_exe_prng_12_io_out_6,rand_exe_prng_12_io_out_5,
    rand_exe_prng_12_io_out_4,rand_exe_prng_12_io_out_3,rand_exe_prng_12_io_out_2,rand_exe_prng_12_io_out_1,
    rand_exe_prng_12_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_12 = {rand_exe_prng_12_io_out_15,rand_exe_prng_12_io_out_14,rand_exe_prng_12_io_out_13,
    rand_exe_prng_12_io_out_12,rand_exe_prng_12_io_out_11,rand_exe_prng_12_io_out_10,rand_exe_prng_12_io_out_9,
    rand_exe_prng_12_io_out_8,rand_exe_lo_12}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_13 = {rand_exe_prng_13_io_out_7,rand_exe_prng_13_io_out_6,rand_exe_prng_13_io_out_5,
    rand_exe_prng_13_io_out_4,rand_exe_prng_13_io_out_3,rand_exe_prng_13_io_out_2,rand_exe_prng_13_io_out_1,
    rand_exe_prng_13_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_13 = {rand_exe_prng_13_io_out_15,rand_exe_prng_13_io_out_14,rand_exe_prng_13_io_out_13,
    rand_exe_prng_13_io_out_12,rand_exe_prng_13_io_out_11,rand_exe_prng_13_io_out_10,rand_exe_prng_13_io_out_9,
    rand_exe_prng_13_io_out_8,rand_exe_lo_13}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_14 = {rand_exe_prng_14_io_out_7,rand_exe_prng_14_io_out_6,rand_exe_prng_14_io_out_5,
    rand_exe_prng_14_io_out_4,rand_exe_prng_14_io_out_3,rand_exe_prng_14_io_out_2,rand_exe_prng_14_io_out_1,
    rand_exe_prng_14_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_14 = {rand_exe_prng_14_io_out_15,rand_exe_prng_14_io_out_14,rand_exe_prng_14_io_out_13,
    rand_exe_prng_14_io_out_12,rand_exe_prng_14_io_out_11,rand_exe_prng_14_io_out_10,rand_exe_prng_14_io_out_9,
    rand_exe_prng_14_io_out_8,rand_exe_lo_14}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_15 = {rand_exe_prng_15_io_out_7,rand_exe_prng_15_io_out_6,rand_exe_prng_15_io_out_5,
    rand_exe_prng_15_io_out_4,rand_exe_prng_15_io_out_3,rand_exe_prng_15_io_out_2,rand_exe_prng_15_io_out_1,
    rand_exe_prng_15_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_15 = {rand_exe_prng_15_io_out_15,rand_exe_prng_15_io_out_14,rand_exe_prng_15_io_out_13,
    rand_exe_prng_15_io_out_12,rand_exe_prng_15_io_out_11,rand_exe_prng_15_io_out_10,rand_exe_prng_15_io_out_9,
    rand_exe_prng_15_io_out_8,rand_exe_lo_15}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_16 = {rand_exe_prng_16_io_out_7,rand_exe_prng_16_io_out_6,rand_exe_prng_16_io_out_5,
    rand_exe_prng_16_io_out_4,rand_exe_prng_16_io_out_3,rand_exe_prng_16_io_out_2,rand_exe_prng_16_io_out_1,
    rand_exe_prng_16_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_16 = {rand_exe_prng_16_io_out_15,rand_exe_prng_16_io_out_14,rand_exe_prng_16_io_out_13,
    rand_exe_prng_16_io_out_12,rand_exe_prng_16_io_out_11,rand_exe_prng_16_io_out_10,rand_exe_prng_16_io_out_9,
    rand_exe_prng_16_io_out_8,rand_exe_lo_16}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_17 = {rand_exe_prng_17_io_out_7,rand_exe_prng_17_io_out_6,rand_exe_prng_17_io_out_5,
    rand_exe_prng_17_io_out_4,rand_exe_prng_17_io_out_3,rand_exe_prng_17_io_out_2,rand_exe_prng_17_io_out_1,
    rand_exe_prng_17_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_17 = {rand_exe_prng_17_io_out_15,rand_exe_prng_17_io_out_14,rand_exe_prng_17_io_out_13,
    rand_exe_prng_17_io_out_12,rand_exe_prng_17_io_out_11,rand_exe_prng_17_io_out_10,rand_exe_prng_17_io_out_9,
    rand_exe_prng_17_io_out_8,rand_exe_lo_17}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_18 = {rand_exe_prng_18_io_out_7,rand_exe_prng_18_io_out_6,rand_exe_prng_18_io_out_5,
    rand_exe_prng_18_io_out_4,rand_exe_prng_18_io_out_3,rand_exe_prng_18_io_out_2,rand_exe_prng_18_io_out_1,
    rand_exe_prng_18_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_18 = {rand_exe_prng_18_io_out_15,rand_exe_prng_18_io_out_14,rand_exe_prng_18_io_out_13,
    rand_exe_prng_18_io_out_12,rand_exe_prng_18_io_out_11,rand_exe_prng_18_io_out_10,rand_exe_prng_18_io_out_9,
    rand_exe_prng_18_io_out_8,rand_exe_lo_18}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_19 = {rand_exe_prng_19_io_out_7,rand_exe_prng_19_io_out_6,rand_exe_prng_19_io_out_5,
    rand_exe_prng_19_io_out_4,rand_exe_prng_19_io_out_3,rand_exe_prng_19_io_out_2,rand_exe_prng_19_io_out_1,
    rand_exe_prng_19_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_19 = {rand_exe_prng_19_io_out_15,rand_exe_prng_19_io_out_14,rand_exe_prng_19_io_out_13,
    rand_exe_prng_19_io_out_12,rand_exe_prng_19_io_out_11,rand_exe_prng_19_io_out_10,rand_exe_prng_19_io_out_9,
    rand_exe_prng_19_io_out_8,rand_exe_lo_19}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_20 = {rand_exe_prng_20_io_out_7,rand_exe_prng_20_io_out_6,rand_exe_prng_20_io_out_5,
    rand_exe_prng_20_io_out_4,rand_exe_prng_20_io_out_3,rand_exe_prng_20_io_out_2,rand_exe_prng_20_io_out_1,
    rand_exe_prng_20_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_20 = {rand_exe_prng_20_io_out_15,rand_exe_prng_20_io_out_14,rand_exe_prng_20_io_out_13,
    rand_exe_prng_20_io_out_12,rand_exe_prng_20_io_out_11,rand_exe_prng_20_io_out_10,rand_exe_prng_20_io_out_9,
    rand_exe_prng_20_io_out_8,rand_exe_lo_20}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_21 = {rand_exe_prng_21_io_out_7,rand_exe_prng_21_io_out_6,rand_exe_prng_21_io_out_5,
    rand_exe_prng_21_io_out_4,rand_exe_prng_21_io_out_3,rand_exe_prng_21_io_out_2,rand_exe_prng_21_io_out_1,
    rand_exe_prng_21_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_21 = {rand_exe_prng_21_io_out_15,rand_exe_prng_21_io_out_14,rand_exe_prng_21_io_out_13,
    rand_exe_prng_21_io_out_12,rand_exe_prng_21_io_out_11,rand_exe_prng_21_io_out_10,rand_exe_prng_21_io_out_9,
    rand_exe_prng_21_io_out_8,rand_exe_lo_21}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_22 = {rand_exe_prng_22_io_out_7,rand_exe_prng_22_io_out_6,rand_exe_prng_22_io_out_5,
    rand_exe_prng_22_io_out_4,rand_exe_prng_22_io_out_3,rand_exe_prng_22_io_out_2,rand_exe_prng_22_io_out_1,
    rand_exe_prng_22_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_22 = {rand_exe_prng_22_io_out_15,rand_exe_prng_22_io_out_14,rand_exe_prng_22_io_out_13,
    rand_exe_prng_22_io_out_12,rand_exe_prng_22_io_out_11,rand_exe_prng_22_io_out_10,rand_exe_prng_22_io_out_9,
    rand_exe_prng_22_io_out_8,rand_exe_lo_22}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_23 = {rand_exe_prng_23_io_out_7,rand_exe_prng_23_io_out_6,rand_exe_prng_23_io_out_5,
    rand_exe_prng_23_io_out_4,rand_exe_prng_23_io_out_3,rand_exe_prng_23_io_out_2,rand_exe_prng_23_io_out_1,
    rand_exe_prng_23_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_23 = {rand_exe_prng_23_io_out_15,rand_exe_prng_23_io_out_14,rand_exe_prng_23_io_out_13,
    rand_exe_prng_23_io_out_12,rand_exe_prng_23_io_out_11,rand_exe_prng_23_io_out_10,rand_exe_prng_23_io_out_9,
    rand_exe_prng_23_io_out_8,rand_exe_lo_23}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_24 = {rand_exe_prng_24_io_out_7,rand_exe_prng_24_io_out_6,rand_exe_prng_24_io_out_5,
    rand_exe_prng_24_io_out_4,rand_exe_prng_24_io_out_3,rand_exe_prng_24_io_out_2,rand_exe_prng_24_io_out_1,
    rand_exe_prng_24_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_24 = {rand_exe_prng_24_io_out_15,rand_exe_prng_24_io_out_14,rand_exe_prng_24_io_out_13,
    rand_exe_prng_24_io_out_12,rand_exe_prng_24_io_out_11,rand_exe_prng_24_io_out_10,rand_exe_prng_24_io_out_9,
    rand_exe_prng_24_io_out_8,rand_exe_lo_24}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_25 = {rand_exe_prng_25_io_out_7,rand_exe_prng_25_io_out_6,rand_exe_prng_25_io_out_5,
    rand_exe_prng_25_io_out_4,rand_exe_prng_25_io_out_3,rand_exe_prng_25_io_out_2,rand_exe_prng_25_io_out_1,
    rand_exe_prng_25_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_25 = {rand_exe_prng_25_io_out_15,rand_exe_prng_25_io_out_14,rand_exe_prng_25_io_out_13,
    rand_exe_prng_25_io_out_12,rand_exe_prng_25_io_out_11,rand_exe_prng_25_io_out_10,rand_exe_prng_25_io_out_9,
    rand_exe_prng_25_io_out_8,rand_exe_lo_25}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_26 = {rand_exe_prng_26_io_out_7,rand_exe_prng_26_io_out_6,rand_exe_prng_26_io_out_5,
    rand_exe_prng_26_io_out_4,rand_exe_prng_26_io_out_3,rand_exe_prng_26_io_out_2,rand_exe_prng_26_io_out_1,
    rand_exe_prng_26_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_26 = {rand_exe_prng_26_io_out_15,rand_exe_prng_26_io_out_14,rand_exe_prng_26_io_out_13,
    rand_exe_prng_26_io_out_12,rand_exe_prng_26_io_out_11,rand_exe_prng_26_io_out_10,rand_exe_prng_26_io_out_9,
    rand_exe_prng_26_io_out_8,rand_exe_lo_26}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_27 = {rand_exe_prng_27_io_out_7,rand_exe_prng_27_io_out_6,rand_exe_prng_27_io_out_5,
    rand_exe_prng_27_io_out_4,rand_exe_prng_27_io_out_3,rand_exe_prng_27_io_out_2,rand_exe_prng_27_io_out_1,
    rand_exe_prng_27_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_27 = {rand_exe_prng_27_io_out_15,rand_exe_prng_27_io_out_14,rand_exe_prng_27_io_out_13,
    rand_exe_prng_27_io_out_12,rand_exe_prng_27_io_out_11,rand_exe_prng_27_io_out_10,rand_exe_prng_27_io_out_9,
    rand_exe_prng_27_io_out_8,rand_exe_lo_27}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_28 = {rand_exe_prng_28_io_out_7,rand_exe_prng_28_io_out_6,rand_exe_prng_28_io_out_5,
    rand_exe_prng_28_io_out_4,rand_exe_prng_28_io_out_3,rand_exe_prng_28_io_out_2,rand_exe_prng_28_io_out_1,
    rand_exe_prng_28_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_28 = {rand_exe_prng_28_io_out_15,rand_exe_prng_28_io_out_14,rand_exe_prng_28_io_out_13,
    rand_exe_prng_28_io_out_12,rand_exe_prng_28_io_out_11,rand_exe_prng_28_io_out_10,rand_exe_prng_28_io_out_9,
    rand_exe_prng_28_io_out_8,rand_exe_lo_28}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_29 = {rand_exe_prng_29_io_out_7,rand_exe_prng_29_io_out_6,rand_exe_prng_29_io_out_5,
    rand_exe_prng_29_io_out_4,rand_exe_prng_29_io_out_3,rand_exe_prng_29_io_out_2,rand_exe_prng_29_io_out_1,
    rand_exe_prng_29_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_29 = {rand_exe_prng_29_io_out_15,rand_exe_prng_29_io_out_14,rand_exe_prng_29_io_out_13,
    rand_exe_prng_29_io_out_12,rand_exe_prng_29_io_out_11,rand_exe_prng_29_io_out_10,rand_exe_prng_29_io_out_9,
    rand_exe_prng_29_io_out_8,rand_exe_lo_29}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_30 = {rand_exe_prng_30_io_out_7,rand_exe_prng_30_io_out_6,rand_exe_prng_30_io_out_5,
    rand_exe_prng_30_io_out_4,rand_exe_prng_30_io_out_3,rand_exe_prng_30_io_out_2,rand_exe_prng_30_io_out_1,
    rand_exe_prng_30_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_30 = {rand_exe_prng_30_io_out_15,rand_exe_prng_30_io_out_14,rand_exe_prng_30_io_out_13,
    rand_exe_prng_30_io_out_12,rand_exe_prng_30_io_out_11,rand_exe_prng_30_io_out_10,rand_exe_prng_30_io_out_9,
    rand_exe_prng_30_io_out_8,rand_exe_lo_30}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_31 = {rand_exe_prng_31_io_out_7,rand_exe_prng_31_io_out_6,rand_exe_prng_31_io_out_5,
    rand_exe_prng_31_io_out_4,rand_exe_prng_31_io_out_3,rand_exe_prng_31_io_out_2,rand_exe_prng_31_io_out_1,
    rand_exe_prng_31_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_31 = {rand_exe_prng_31_io_out_15,rand_exe_prng_31_io_out_14,rand_exe_prng_31_io_out_13,
    rand_exe_prng_31_io_out_12,rand_exe_prng_31_io_out_11,rand_exe_prng_31_io_out_10,rand_exe_prng_31_io_out_9,
    rand_exe_prng_31_io_out_8,rand_exe_lo_31}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_32 = {rand_exe_prng_32_io_out_7,rand_exe_prng_32_io_out_6,rand_exe_prng_32_io_out_5,
    rand_exe_prng_32_io_out_4,rand_exe_prng_32_io_out_3,rand_exe_prng_32_io_out_2,rand_exe_prng_32_io_out_1,
    rand_exe_prng_32_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_32 = {rand_exe_prng_32_io_out_15,rand_exe_prng_32_io_out_14,rand_exe_prng_32_io_out_13,
    rand_exe_prng_32_io_out_12,rand_exe_prng_32_io_out_11,rand_exe_prng_32_io_out_10,rand_exe_prng_32_io_out_9,
    rand_exe_prng_32_io_out_8,rand_exe_lo_32}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_33 = {rand_exe_prng_33_io_out_7,rand_exe_prng_33_io_out_6,rand_exe_prng_33_io_out_5,
    rand_exe_prng_33_io_out_4,rand_exe_prng_33_io_out_3,rand_exe_prng_33_io_out_2,rand_exe_prng_33_io_out_1,
    rand_exe_prng_33_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_33 = {rand_exe_prng_33_io_out_15,rand_exe_prng_33_io_out_14,rand_exe_prng_33_io_out_13,
    rand_exe_prng_33_io_out_12,rand_exe_prng_33_io_out_11,rand_exe_prng_33_io_out_10,rand_exe_prng_33_io_out_9,
    rand_exe_prng_33_io_out_8,rand_exe_lo_33}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_34 = {rand_exe_prng_34_io_out_7,rand_exe_prng_34_io_out_6,rand_exe_prng_34_io_out_5,
    rand_exe_prng_34_io_out_4,rand_exe_prng_34_io_out_3,rand_exe_prng_34_io_out_2,rand_exe_prng_34_io_out_1,
    rand_exe_prng_34_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_34 = {rand_exe_prng_34_io_out_15,rand_exe_prng_34_io_out_14,rand_exe_prng_34_io_out_13,
    rand_exe_prng_34_io_out_12,rand_exe_prng_34_io_out_11,rand_exe_prng_34_io_out_10,rand_exe_prng_34_io_out_9,
    rand_exe_prng_34_io_out_8,rand_exe_lo_34}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_35 = {rand_exe_prng_35_io_out_7,rand_exe_prng_35_io_out_6,rand_exe_prng_35_io_out_5,
    rand_exe_prng_35_io_out_4,rand_exe_prng_35_io_out_3,rand_exe_prng_35_io_out_2,rand_exe_prng_35_io_out_1,
    rand_exe_prng_35_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_35 = {rand_exe_prng_35_io_out_15,rand_exe_prng_35_io_out_14,rand_exe_prng_35_io_out_13,
    rand_exe_prng_35_io_out_12,rand_exe_prng_35_io_out_11,rand_exe_prng_35_io_out_10,rand_exe_prng_35_io_out_9,
    rand_exe_prng_35_io_out_8,rand_exe_lo_35}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_36 = {rand_exe_prng_36_io_out_7,rand_exe_prng_36_io_out_6,rand_exe_prng_36_io_out_5,
    rand_exe_prng_36_io_out_4,rand_exe_prng_36_io_out_3,rand_exe_prng_36_io_out_2,rand_exe_prng_36_io_out_1,
    rand_exe_prng_36_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_36 = {rand_exe_prng_36_io_out_15,rand_exe_prng_36_io_out_14,rand_exe_prng_36_io_out_13,
    rand_exe_prng_36_io_out_12,rand_exe_prng_36_io_out_11,rand_exe_prng_36_io_out_10,rand_exe_prng_36_io_out_9,
    rand_exe_prng_36_io_out_8,rand_exe_lo_36}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_37 = {rand_exe_prng_37_io_out_7,rand_exe_prng_37_io_out_6,rand_exe_prng_37_io_out_5,
    rand_exe_prng_37_io_out_4,rand_exe_prng_37_io_out_3,rand_exe_prng_37_io_out_2,rand_exe_prng_37_io_out_1,
    rand_exe_prng_37_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_37 = {rand_exe_prng_37_io_out_15,rand_exe_prng_37_io_out_14,rand_exe_prng_37_io_out_13,
    rand_exe_prng_37_io_out_12,rand_exe_prng_37_io_out_11,rand_exe_prng_37_io_out_10,rand_exe_prng_37_io_out_9,
    rand_exe_prng_37_io_out_8,rand_exe_lo_37}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_38 = {rand_exe_prng_38_io_out_7,rand_exe_prng_38_io_out_6,rand_exe_prng_38_io_out_5,
    rand_exe_prng_38_io_out_4,rand_exe_prng_38_io_out_3,rand_exe_prng_38_io_out_2,rand_exe_prng_38_io_out_1,
    rand_exe_prng_38_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_38 = {rand_exe_prng_38_io_out_15,rand_exe_prng_38_io_out_14,rand_exe_prng_38_io_out_13,
    rand_exe_prng_38_io_out_12,rand_exe_prng_38_io_out_11,rand_exe_prng_38_io_out_10,rand_exe_prng_38_io_out_9,
    rand_exe_prng_38_io_out_8,rand_exe_lo_38}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_39 = {rand_exe_prng_39_io_out_7,rand_exe_prng_39_io_out_6,rand_exe_prng_39_io_out_5,
    rand_exe_prng_39_io_out_4,rand_exe_prng_39_io_out_3,rand_exe_prng_39_io_out_2,rand_exe_prng_39_io_out_1,
    rand_exe_prng_39_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_39 = {rand_exe_prng_39_io_out_15,rand_exe_prng_39_io_out_14,rand_exe_prng_39_io_out_13,
    rand_exe_prng_39_io_out_12,rand_exe_prng_39_io_out_11,rand_exe_prng_39_io_out_10,rand_exe_prng_39_io_out_9,
    rand_exe_prng_39_io_out_8,rand_exe_lo_39}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_40 = {rand_exe_prng_40_io_out_7,rand_exe_prng_40_io_out_6,rand_exe_prng_40_io_out_5,
    rand_exe_prng_40_io_out_4,rand_exe_prng_40_io_out_3,rand_exe_prng_40_io_out_2,rand_exe_prng_40_io_out_1,
    rand_exe_prng_40_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_40 = {rand_exe_prng_40_io_out_15,rand_exe_prng_40_io_out_14,rand_exe_prng_40_io_out_13,
    rand_exe_prng_40_io_out_12,rand_exe_prng_40_io_out_11,rand_exe_prng_40_io_out_10,rand_exe_prng_40_io_out_9,
    rand_exe_prng_40_io_out_8,rand_exe_lo_40}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_41 = {rand_exe_prng_41_io_out_7,rand_exe_prng_41_io_out_6,rand_exe_prng_41_io_out_5,
    rand_exe_prng_41_io_out_4,rand_exe_prng_41_io_out_3,rand_exe_prng_41_io_out_2,rand_exe_prng_41_io_out_1,
    rand_exe_prng_41_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_41 = {rand_exe_prng_41_io_out_15,rand_exe_prng_41_io_out_14,rand_exe_prng_41_io_out_13,
    rand_exe_prng_41_io_out_12,rand_exe_prng_41_io_out_11,rand_exe_prng_41_io_out_10,rand_exe_prng_41_io_out_9,
    rand_exe_prng_41_io_out_8,rand_exe_lo_41}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_42 = {rand_exe_prng_42_io_out_7,rand_exe_prng_42_io_out_6,rand_exe_prng_42_io_out_5,
    rand_exe_prng_42_io_out_4,rand_exe_prng_42_io_out_3,rand_exe_prng_42_io_out_2,rand_exe_prng_42_io_out_1,
    rand_exe_prng_42_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_42 = {rand_exe_prng_42_io_out_15,rand_exe_prng_42_io_out_14,rand_exe_prng_42_io_out_13,
    rand_exe_prng_42_io_out_12,rand_exe_prng_42_io_out_11,rand_exe_prng_42_io_out_10,rand_exe_prng_42_io_out_9,
    rand_exe_prng_42_io_out_8,rand_exe_lo_42}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_43 = {rand_exe_prng_43_io_out_7,rand_exe_prng_43_io_out_6,rand_exe_prng_43_io_out_5,
    rand_exe_prng_43_io_out_4,rand_exe_prng_43_io_out_3,rand_exe_prng_43_io_out_2,rand_exe_prng_43_io_out_1,
    rand_exe_prng_43_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_43 = {rand_exe_prng_43_io_out_15,rand_exe_prng_43_io_out_14,rand_exe_prng_43_io_out_13,
    rand_exe_prng_43_io_out_12,rand_exe_prng_43_io_out_11,rand_exe_prng_43_io_out_10,rand_exe_prng_43_io_out_9,
    rand_exe_prng_43_io_out_8,rand_exe_lo_43}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_44 = {rand_exe_prng_44_io_out_7,rand_exe_prng_44_io_out_6,rand_exe_prng_44_io_out_5,
    rand_exe_prng_44_io_out_4,rand_exe_prng_44_io_out_3,rand_exe_prng_44_io_out_2,rand_exe_prng_44_io_out_1,
    rand_exe_prng_44_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_44 = {rand_exe_prng_44_io_out_15,rand_exe_prng_44_io_out_14,rand_exe_prng_44_io_out_13,
    rand_exe_prng_44_io_out_12,rand_exe_prng_44_io_out_11,rand_exe_prng_44_io_out_10,rand_exe_prng_44_io_out_9,
    rand_exe_prng_44_io_out_8,rand_exe_lo_44}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_45 = {rand_exe_prng_45_io_out_7,rand_exe_prng_45_io_out_6,rand_exe_prng_45_io_out_5,
    rand_exe_prng_45_io_out_4,rand_exe_prng_45_io_out_3,rand_exe_prng_45_io_out_2,rand_exe_prng_45_io_out_1,
    rand_exe_prng_45_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_45 = {rand_exe_prng_45_io_out_15,rand_exe_prng_45_io_out_14,rand_exe_prng_45_io_out_13,
    rand_exe_prng_45_io_out_12,rand_exe_prng_45_io_out_11,rand_exe_prng_45_io_out_10,rand_exe_prng_45_io_out_9,
    rand_exe_prng_45_io_out_8,rand_exe_lo_45}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_46 = {rand_exe_prng_46_io_out_7,rand_exe_prng_46_io_out_6,rand_exe_prng_46_io_out_5,
    rand_exe_prng_46_io_out_4,rand_exe_prng_46_io_out_3,rand_exe_prng_46_io_out_2,rand_exe_prng_46_io_out_1,
    rand_exe_prng_46_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_46 = {rand_exe_prng_46_io_out_15,rand_exe_prng_46_io_out_14,rand_exe_prng_46_io_out_13,
    rand_exe_prng_46_io_out_12,rand_exe_prng_46_io_out_11,rand_exe_prng_46_io_out_10,rand_exe_prng_46_io_out_9,
    rand_exe_prng_46_io_out_8,rand_exe_lo_46}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_47 = {rand_exe_prng_47_io_out_7,rand_exe_prng_47_io_out_6,rand_exe_prng_47_io_out_5,
    rand_exe_prng_47_io_out_4,rand_exe_prng_47_io_out_3,rand_exe_prng_47_io_out_2,rand_exe_prng_47_io_out_1,
    rand_exe_prng_47_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_47 = {rand_exe_prng_47_io_out_15,rand_exe_prng_47_io_out_14,rand_exe_prng_47_io_out_13,
    rand_exe_prng_47_io_out_12,rand_exe_prng_47_io_out_11,rand_exe_prng_47_io_out_10,rand_exe_prng_47_io_out_9,
    rand_exe_prng_47_io_out_8,rand_exe_lo_47}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_48 = {rand_exe_prng_48_io_out_7,rand_exe_prng_48_io_out_6,rand_exe_prng_48_io_out_5,
    rand_exe_prng_48_io_out_4,rand_exe_prng_48_io_out_3,rand_exe_prng_48_io_out_2,rand_exe_prng_48_io_out_1,
    rand_exe_prng_48_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_48 = {rand_exe_prng_48_io_out_15,rand_exe_prng_48_io_out_14,rand_exe_prng_48_io_out_13,
    rand_exe_prng_48_io_out_12,rand_exe_prng_48_io_out_11,rand_exe_prng_48_io_out_10,rand_exe_prng_48_io_out_9,
    rand_exe_prng_48_io_out_8,rand_exe_lo_48}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_49 = {rand_exe_prng_49_io_out_7,rand_exe_prng_49_io_out_6,rand_exe_prng_49_io_out_5,
    rand_exe_prng_49_io_out_4,rand_exe_prng_49_io_out_3,rand_exe_prng_49_io_out_2,rand_exe_prng_49_io_out_1,
    rand_exe_prng_49_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_49 = {rand_exe_prng_49_io_out_15,rand_exe_prng_49_io_out_14,rand_exe_prng_49_io_out_13,
    rand_exe_prng_49_io_out_12,rand_exe_prng_49_io_out_11,rand_exe_prng_49_io_out_10,rand_exe_prng_49_io_out_9,
    rand_exe_prng_49_io_out_8,rand_exe_lo_49}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_50 = {rand_exe_prng_50_io_out_7,rand_exe_prng_50_io_out_6,rand_exe_prng_50_io_out_5,
    rand_exe_prng_50_io_out_4,rand_exe_prng_50_io_out_3,rand_exe_prng_50_io_out_2,rand_exe_prng_50_io_out_1,
    rand_exe_prng_50_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_50 = {rand_exe_prng_50_io_out_15,rand_exe_prng_50_io_out_14,rand_exe_prng_50_io_out_13,
    rand_exe_prng_50_io_out_12,rand_exe_prng_50_io_out_11,rand_exe_prng_50_io_out_10,rand_exe_prng_50_io_out_9,
    rand_exe_prng_50_io_out_8,rand_exe_lo_50}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_51 = {rand_exe_prng_51_io_out_7,rand_exe_prng_51_io_out_6,rand_exe_prng_51_io_out_5,
    rand_exe_prng_51_io_out_4,rand_exe_prng_51_io_out_3,rand_exe_prng_51_io_out_2,rand_exe_prng_51_io_out_1,
    rand_exe_prng_51_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_51 = {rand_exe_prng_51_io_out_15,rand_exe_prng_51_io_out_14,rand_exe_prng_51_io_out_13,
    rand_exe_prng_51_io_out_12,rand_exe_prng_51_io_out_11,rand_exe_prng_51_io_out_10,rand_exe_prng_51_io_out_9,
    rand_exe_prng_51_io_out_8,rand_exe_lo_51}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_52 = {rand_exe_prng_52_io_out_7,rand_exe_prng_52_io_out_6,rand_exe_prng_52_io_out_5,
    rand_exe_prng_52_io_out_4,rand_exe_prng_52_io_out_3,rand_exe_prng_52_io_out_2,rand_exe_prng_52_io_out_1,
    rand_exe_prng_52_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_52 = {rand_exe_prng_52_io_out_15,rand_exe_prng_52_io_out_14,rand_exe_prng_52_io_out_13,
    rand_exe_prng_52_io_out_12,rand_exe_prng_52_io_out_11,rand_exe_prng_52_io_out_10,rand_exe_prng_52_io_out_9,
    rand_exe_prng_52_io_out_8,rand_exe_lo_52}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_53 = {rand_exe_prng_53_io_out_7,rand_exe_prng_53_io_out_6,rand_exe_prng_53_io_out_5,
    rand_exe_prng_53_io_out_4,rand_exe_prng_53_io_out_3,rand_exe_prng_53_io_out_2,rand_exe_prng_53_io_out_1,
    rand_exe_prng_53_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_53 = {rand_exe_prng_53_io_out_15,rand_exe_prng_53_io_out_14,rand_exe_prng_53_io_out_13,
    rand_exe_prng_53_io_out_12,rand_exe_prng_53_io_out_11,rand_exe_prng_53_io_out_10,rand_exe_prng_53_io_out_9,
    rand_exe_prng_53_io_out_8,rand_exe_lo_53}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_54 = {rand_exe_prng_54_io_out_7,rand_exe_prng_54_io_out_6,rand_exe_prng_54_io_out_5,
    rand_exe_prng_54_io_out_4,rand_exe_prng_54_io_out_3,rand_exe_prng_54_io_out_2,rand_exe_prng_54_io_out_1,
    rand_exe_prng_54_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_54 = {rand_exe_prng_54_io_out_15,rand_exe_prng_54_io_out_14,rand_exe_prng_54_io_out_13,
    rand_exe_prng_54_io_out_12,rand_exe_prng_54_io_out_11,rand_exe_prng_54_io_out_10,rand_exe_prng_54_io_out_9,
    rand_exe_prng_54_io_out_8,rand_exe_lo_54}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_55 = {rand_exe_prng_55_io_out_7,rand_exe_prng_55_io_out_6,rand_exe_prng_55_io_out_5,
    rand_exe_prng_55_io_out_4,rand_exe_prng_55_io_out_3,rand_exe_prng_55_io_out_2,rand_exe_prng_55_io_out_1,
    rand_exe_prng_55_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_55 = {rand_exe_prng_55_io_out_15,rand_exe_prng_55_io_out_14,rand_exe_prng_55_io_out_13,
    rand_exe_prng_55_io_out_12,rand_exe_prng_55_io_out_11,rand_exe_prng_55_io_out_10,rand_exe_prng_55_io_out_9,
    rand_exe_prng_55_io_out_8,rand_exe_lo_55}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_56 = {rand_exe_prng_56_io_out_7,rand_exe_prng_56_io_out_6,rand_exe_prng_56_io_out_5,
    rand_exe_prng_56_io_out_4,rand_exe_prng_56_io_out_3,rand_exe_prng_56_io_out_2,rand_exe_prng_56_io_out_1,
    rand_exe_prng_56_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_56 = {rand_exe_prng_56_io_out_15,rand_exe_prng_56_io_out_14,rand_exe_prng_56_io_out_13,
    rand_exe_prng_56_io_out_12,rand_exe_prng_56_io_out_11,rand_exe_prng_56_io_out_10,rand_exe_prng_56_io_out_9,
    rand_exe_prng_56_io_out_8,rand_exe_lo_56}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_57 = {rand_exe_prng_57_io_out_7,rand_exe_prng_57_io_out_6,rand_exe_prng_57_io_out_5,
    rand_exe_prng_57_io_out_4,rand_exe_prng_57_io_out_3,rand_exe_prng_57_io_out_2,rand_exe_prng_57_io_out_1,
    rand_exe_prng_57_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_57 = {rand_exe_prng_57_io_out_15,rand_exe_prng_57_io_out_14,rand_exe_prng_57_io_out_13,
    rand_exe_prng_57_io_out_12,rand_exe_prng_57_io_out_11,rand_exe_prng_57_io_out_10,rand_exe_prng_57_io_out_9,
    rand_exe_prng_57_io_out_8,rand_exe_lo_57}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_58 = {rand_exe_prng_58_io_out_7,rand_exe_prng_58_io_out_6,rand_exe_prng_58_io_out_5,
    rand_exe_prng_58_io_out_4,rand_exe_prng_58_io_out_3,rand_exe_prng_58_io_out_2,rand_exe_prng_58_io_out_1,
    rand_exe_prng_58_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_58 = {rand_exe_prng_58_io_out_15,rand_exe_prng_58_io_out_14,rand_exe_prng_58_io_out_13,
    rand_exe_prng_58_io_out_12,rand_exe_prng_58_io_out_11,rand_exe_prng_58_io_out_10,rand_exe_prng_58_io_out_9,
    rand_exe_prng_58_io_out_8,rand_exe_lo_58}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_59 = {rand_exe_prng_59_io_out_7,rand_exe_prng_59_io_out_6,rand_exe_prng_59_io_out_5,
    rand_exe_prng_59_io_out_4,rand_exe_prng_59_io_out_3,rand_exe_prng_59_io_out_2,rand_exe_prng_59_io_out_1,
    rand_exe_prng_59_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_59 = {rand_exe_prng_59_io_out_15,rand_exe_prng_59_io_out_14,rand_exe_prng_59_io_out_13,
    rand_exe_prng_59_io_out_12,rand_exe_prng_59_io_out_11,rand_exe_prng_59_io_out_10,rand_exe_prng_59_io_out_9,
    rand_exe_prng_59_io_out_8,rand_exe_lo_59}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_60 = {rand_exe_prng_60_io_out_7,rand_exe_prng_60_io_out_6,rand_exe_prng_60_io_out_5,
    rand_exe_prng_60_io_out_4,rand_exe_prng_60_io_out_3,rand_exe_prng_60_io_out_2,rand_exe_prng_60_io_out_1,
    rand_exe_prng_60_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_60 = {rand_exe_prng_60_io_out_15,rand_exe_prng_60_io_out_14,rand_exe_prng_60_io_out_13,
    rand_exe_prng_60_io_out_12,rand_exe_prng_60_io_out_11,rand_exe_prng_60_io_out_10,rand_exe_prng_60_io_out_9,
    rand_exe_prng_60_io_out_8,rand_exe_lo_60}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_61 = {rand_exe_prng_61_io_out_7,rand_exe_prng_61_io_out_6,rand_exe_prng_61_io_out_5,
    rand_exe_prng_61_io_out_4,rand_exe_prng_61_io_out_3,rand_exe_prng_61_io_out_2,rand_exe_prng_61_io_out_1,
    rand_exe_prng_61_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_61 = {rand_exe_prng_61_io_out_15,rand_exe_prng_61_io_out_14,rand_exe_prng_61_io_out_13,
    rand_exe_prng_61_io_out_12,rand_exe_prng_61_io_out_11,rand_exe_prng_61_io_out_10,rand_exe_prng_61_io_out_9,
    rand_exe_prng_61_io_out_8,rand_exe_lo_61}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_62 = {rand_exe_prng_62_io_out_7,rand_exe_prng_62_io_out_6,rand_exe_prng_62_io_out_5,
    rand_exe_prng_62_io_out_4,rand_exe_prng_62_io_out_3,rand_exe_prng_62_io_out_2,rand_exe_prng_62_io_out_1,
    rand_exe_prng_62_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_62 = {rand_exe_prng_62_io_out_15,rand_exe_prng_62_io_out_14,rand_exe_prng_62_io_out_13,
    rand_exe_prng_62_io_out_12,rand_exe_prng_62_io_out_11,rand_exe_prng_62_io_out_10,rand_exe_prng_62_io_out_9,
    rand_exe_prng_62_io_out_8,rand_exe_lo_62}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_63 = {rand_exe_prng_63_io_out_7,rand_exe_prng_63_io_out_6,rand_exe_prng_63_io_out_5,
    rand_exe_prng_63_io_out_4,rand_exe_prng_63_io_out_3,rand_exe_prng_63_io_out_2,rand_exe_prng_63_io_out_1,
    rand_exe_prng_63_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_63 = {rand_exe_prng_63_io_out_15,rand_exe_prng_63_io_out_14,rand_exe_prng_63_io_out_13,
    rand_exe_prng_63_io_out_12,rand_exe_prng_63_io_out_11,rand_exe_prng_63_io_out_10,rand_exe_prng_63_io_out_9,
    rand_exe_prng_63_io_out_8,rand_exe_lo_63}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_64 = {rand_exe_prng_64_io_out_7,rand_exe_prng_64_io_out_6,rand_exe_prng_64_io_out_5,
    rand_exe_prng_64_io_out_4,rand_exe_prng_64_io_out_3,rand_exe_prng_64_io_out_2,rand_exe_prng_64_io_out_1,
    rand_exe_prng_64_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_64 = {rand_exe_prng_64_io_out_15,rand_exe_prng_64_io_out_14,rand_exe_prng_64_io_out_13,
    rand_exe_prng_64_io_out_12,rand_exe_prng_64_io_out_11,rand_exe_prng_64_io_out_10,rand_exe_prng_64_io_out_9,
    rand_exe_prng_64_io_out_8,rand_exe_lo_64}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_65 = {rand_exe_prng_65_io_out_7,rand_exe_prng_65_io_out_6,rand_exe_prng_65_io_out_5,
    rand_exe_prng_65_io_out_4,rand_exe_prng_65_io_out_3,rand_exe_prng_65_io_out_2,rand_exe_prng_65_io_out_1,
    rand_exe_prng_65_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_65 = {rand_exe_prng_65_io_out_15,rand_exe_prng_65_io_out_14,rand_exe_prng_65_io_out_13,
    rand_exe_prng_65_io_out_12,rand_exe_prng_65_io_out_11,rand_exe_prng_65_io_out_10,rand_exe_prng_65_io_out_9,
    rand_exe_prng_65_io_out_8,rand_exe_lo_65}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_66 = {rand_exe_prng_66_io_out_7,rand_exe_prng_66_io_out_6,rand_exe_prng_66_io_out_5,
    rand_exe_prng_66_io_out_4,rand_exe_prng_66_io_out_3,rand_exe_prng_66_io_out_2,rand_exe_prng_66_io_out_1,
    rand_exe_prng_66_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_66 = {rand_exe_prng_66_io_out_15,rand_exe_prng_66_io_out_14,rand_exe_prng_66_io_out_13,
    rand_exe_prng_66_io_out_12,rand_exe_prng_66_io_out_11,rand_exe_prng_66_io_out_10,rand_exe_prng_66_io_out_9,
    rand_exe_prng_66_io_out_8,rand_exe_lo_66}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_67 = {rand_exe_prng_67_io_out_7,rand_exe_prng_67_io_out_6,rand_exe_prng_67_io_out_5,
    rand_exe_prng_67_io_out_4,rand_exe_prng_67_io_out_3,rand_exe_prng_67_io_out_2,rand_exe_prng_67_io_out_1,
    rand_exe_prng_67_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_67 = {rand_exe_prng_67_io_out_15,rand_exe_prng_67_io_out_14,rand_exe_prng_67_io_out_13,
    rand_exe_prng_67_io_out_12,rand_exe_prng_67_io_out_11,rand_exe_prng_67_io_out_10,rand_exe_prng_67_io_out_9,
    rand_exe_prng_67_io_out_8,rand_exe_lo_67}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_68 = {rand_exe_prng_68_io_out_7,rand_exe_prng_68_io_out_6,rand_exe_prng_68_io_out_5,
    rand_exe_prng_68_io_out_4,rand_exe_prng_68_io_out_3,rand_exe_prng_68_io_out_2,rand_exe_prng_68_io_out_1,
    rand_exe_prng_68_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_68 = {rand_exe_prng_68_io_out_15,rand_exe_prng_68_io_out_14,rand_exe_prng_68_io_out_13,
    rand_exe_prng_68_io_out_12,rand_exe_prng_68_io_out_11,rand_exe_prng_68_io_out_10,rand_exe_prng_68_io_out_9,
    rand_exe_prng_68_io_out_8,rand_exe_lo_68}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_69 = {rand_exe_prng_69_io_out_7,rand_exe_prng_69_io_out_6,rand_exe_prng_69_io_out_5,
    rand_exe_prng_69_io_out_4,rand_exe_prng_69_io_out_3,rand_exe_prng_69_io_out_2,rand_exe_prng_69_io_out_1,
    rand_exe_prng_69_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_69 = {rand_exe_prng_69_io_out_15,rand_exe_prng_69_io_out_14,rand_exe_prng_69_io_out_13,
    rand_exe_prng_69_io_out_12,rand_exe_prng_69_io_out_11,rand_exe_prng_69_io_out_10,rand_exe_prng_69_io_out_9,
    rand_exe_prng_69_io_out_8,rand_exe_lo_69}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_70 = {rand_exe_prng_70_io_out_7,rand_exe_prng_70_io_out_6,rand_exe_prng_70_io_out_5,
    rand_exe_prng_70_io_out_4,rand_exe_prng_70_io_out_3,rand_exe_prng_70_io_out_2,rand_exe_prng_70_io_out_1,
    rand_exe_prng_70_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_70 = {rand_exe_prng_70_io_out_15,rand_exe_prng_70_io_out_14,rand_exe_prng_70_io_out_13,
    rand_exe_prng_70_io_out_12,rand_exe_prng_70_io_out_11,rand_exe_prng_70_io_out_10,rand_exe_prng_70_io_out_9,
    rand_exe_prng_70_io_out_8,rand_exe_lo_70}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_71 = {rand_exe_prng_71_io_out_7,rand_exe_prng_71_io_out_6,rand_exe_prng_71_io_out_5,
    rand_exe_prng_71_io_out_4,rand_exe_prng_71_io_out_3,rand_exe_prng_71_io_out_2,rand_exe_prng_71_io_out_1,
    rand_exe_prng_71_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_71 = {rand_exe_prng_71_io_out_15,rand_exe_prng_71_io_out_14,rand_exe_prng_71_io_out_13,
    rand_exe_prng_71_io_out_12,rand_exe_prng_71_io_out_11,rand_exe_prng_71_io_out_10,rand_exe_prng_71_io_out_9,
    rand_exe_prng_71_io_out_8,rand_exe_lo_71}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_72 = {rand_exe_prng_72_io_out_7,rand_exe_prng_72_io_out_6,rand_exe_prng_72_io_out_5,
    rand_exe_prng_72_io_out_4,rand_exe_prng_72_io_out_3,rand_exe_prng_72_io_out_2,rand_exe_prng_72_io_out_1,
    rand_exe_prng_72_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_72 = {rand_exe_prng_72_io_out_15,rand_exe_prng_72_io_out_14,rand_exe_prng_72_io_out_13,
    rand_exe_prng_72_io_out_12,rand_exe_prng_72_io_out_11,rand_exe_prng_72_io_out_10,rand_exe_prng_72_io_out_9,
    rand_exe_prng_72_io_out_8,rand_exe_lo_72}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_73 = {rand_exe_prng_73_io_out_7,rand_exe_prng_73_io_out_6,rand_exe_prng_73_io_out_5,
    rand_exe_prng_73_io_out_4,rand_exe_prng_73_io_out_3,rand_exe_prng_73_io_out_2,rand_exe_prng_73_io_out_1,
    rand_exe_prng_73_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_73 = {rand_exe_prng_73_io_out_15,rand_exe_prng_73_io_out_14,rand_exe_prng_73_io_out_13,
    rand_exe_prng_73_io_out_12,rand_exe_prng_73_io_out_11,rand_exe_prng_73_io_out_10,rand_exe_prng_73_io_out_9,
    rand_exe_prng_73_io_out_8,rand_exe_lo_73}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_74 = {rand_exe_prng_74_io_out_7,rand_exe_prng_74_io_out_6,rand_exe_prng_74_io_out_5,
    rand_exe_prng_74_io_out_4,rand_exe_prng_74_io_out_3,rand_exe_prng_74_io_out_2,rand_exe_prng_74_io_out_1,
    rand_exe_prng_74_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_74 = {rand_exe_prng_74_io_out_15,rand_exe_prng_74_io_out_14,rand_exe_prng_74_io_out_13,
    rand_exe_prng_74_io_out_12,rand_exe_prng_74_io_out_11,rand_exe_prng_74_io_out_10,rand_exe_prng_74_io_out_9,
    rand_exe_prng_74_io_out_8,rand_exe_lo_74}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_75 = {rand_exe_prng_75_io_out_7,rand_exe_prng_75_io_out_6,rand_exe_prng_75_io_out_5,
    rand_exe_prng_75_io_out_4,rand_exe_prng_75_io_out_3,rand_exe_prng_75_io_out_2,rand_exe_prng_75_io_out_1,
    rand_exe_prng_75_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_75 = {rand_exe_prng_75_io_out_15,rand_exe_prng_75_io_out_14,rand_exe_prng_75_io_out_13,
    rand_exe_prng_75_io_out_12,rand_exe_prng_75_io_out_11,rand_exe_prng_75_io_out_10,rand_exe_prng_75_io_out_9,
    rand_exe_prng_75_io_out_8,rand_exe_lo_75}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_76 = {rand_exe_prng_76_io_out_7,rand_exe_prng_76_io_out_6,rand_exe_prng_76_io_out_5,
    rand_exe_prng_76_io_out_4,rand_exe_prng_76_io_out_3,rand_exe_prng_76_io_out_2,rand_exe_prng_76_io_out_1,
    rand_exe_prng_76_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_76 = {rand_exe_prng_76_io_out_15,rand_exe_prng_76_io_out_14,rand_exe_prng_76_io_out_13,
    rand_exe_prng_76_io_out_12,rand_exe_prng_76_io_out_11,rand_exe_prng_76_io_out_10,rand_exe_prng_76_io_out_9,
    rand_exe_prng_76_io_out_8,rand_exe_lo_76}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_77 = {rand_exe_prng_77_io_out_7,rand_exe_prng_77_io_out_6,rand_exe_prng_77_io_out_5,
    rand_exe_prng_77_io_out_4,rand_exe_prng_77_io_out_3,rand_exe_prng_77_io_out_2,rand_exe_prng_77_io_out_1,
    rand_exe_prng_77_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_77 = {rand_exe_prng_77_io_out_15,rand_exe_prng_77_io_out_14,rand_exe_prng_77_io_out_13,
    rand_exe_prng_77_io_out_12,rand_exe_prng_77_io_out_11,rand_exe_prng_77_io_out_10,rand_exe_prng_77_io_out_9,
    rand_exe_prng_77_io_out_8,rand_exe_lo_77}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_78 = {rand_exe_prng_78_io_out_7,rand_exe_prng_78_io_out_6,rand_exe_prng_78_io_out_5,
    rand_exe_prng_78_io_out_4,rand_exe_prng_78_io_out_3,rand_exe_prng_78_io_out_2,rand_exe_prng_78_io_out_1,
    rand_exe_prng_78_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_78 = {rand_exe_prng_78_io_out_15,rand_exe_prng_78_io_out_14,rand_exe_prng_78_io_out_13,
    rand_exe_prng_78_io_out_12,rand_exe_prng_78_io_out_11,rand_exe_prng_78_io_out_10,rand_exe_prng_78_io_out_9,
    rand_exe_prng_78_io_out_8,rand_exe_lo_78}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_79 = {rand_exe_prng_79_io_out_7,rand_exe_prng_79_io_out_6,rand_exe_prng_79_io_out_5,
    rand_exe_prng_79_io_out_4,rand_exe_prng_79_io_out_3,rand_exe_prng_79_io_out_2,rand_exe_prng_79_io_out_1,
    rand_exe_prng_79_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_79 = {rand_exe_prng_79_io_out_15,rand_exe_prng_79_io_out_14,rand_exe_prng_79_io_out_13,
    rand_exe_prng_79_io_out_12,rand_exe_prng_79_io_out_11,rand_exe_prng_79_io_out_10,rand_exe_prng_79_io_out_9,
    rand_exe_prng_79_io_out_8,rand_exe_lo_79}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_80 = {rand_exe_prng_80_io_out_7,rand_exe_prng_80_io_out_6,rand_exe_prng_80_io_out_5,
    rand_exe_prng_80_io_out_4,rand_exe_prng_80_io_out_3,rand_exe_prng_80_io_out_2,rand_exe_prng_80_io_out_1,
    rand_exe_prng_80_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_80 = {rand_exe_prng_80_io_out_15,rand_exe_prng_80_io_out_14,rand_exe_prng_80_io_out_13,
    rand_exe_prng_80_io_out_12,rand_exe_prng_80_io_out_11,rand_exe_prng_80_io_out_10,rand_exe_prng_80_io_out_9,
    rand_exe_prng_80_io_out_8,rand_exe_lo_80}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_81 = {rand_exe_prng_81_io_out_7,rand_exe_prng_81_io_out_6,rand_exe_prng_81_io_out_5,
    rand_exe_prng_81_io_out_4,rand_exe_prng_81_io_out_3,rand_exe_prng_81_io_out_2,rand_exe_prng_81_io_out_1,
    rand_exe_prng_81_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_81 = {rand_exe_prng_81_io_out_15,rand_exe_prng_81_io_out_14,rand_exe_prng_81_io_out_13,
    rand_exe_prng_81_io_out_12,rand_exe_prng_81_io_out_11,rand_exe_prng_81_io_out_10,rand_exe_prng_81_io_out_9,
    rand_exe_prng_81_io_out_8,rand_exe_lo_81}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_82 = {rand_exe_prng_82_io_out_7,rand_exe_prng_82_io_out_6,rand_exe_prng_82_io_out_5,
    rand_exe_prng_82_io_out_4,rand_exe_prng_82_io_out_3,rand_exe_prng_82_io_out_2,rand_exe_prng_82_io_out_1,
    rand_exe_prng_82_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_82 = {rand_exe_prng_82_io_out_15,rand_exe_prng_82_io_out_14,rand_exe_prng_82_io_out_13,
    rand_exe_prng_82_io_out_12,rand_exe_prng_82_io_out_11,rand_exe_prng_82_io_out_10,rand_exe_prng_82_io_out_9,
    rand_exe_prng_82_io_out_8,rand_exe_lo_82}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_83 = {rand_exe_prng_83_io_out_7,rand_exe_prng_83_io_out_6,rand_exe_prng_83_io_out_5,
    rand_exe_prng_83_io_out_4,rand_exe_prng_83_io_out_3,rand_exe_prng_83_io_out_2,rand_exe_prng_83_io_out_1,
    rand_exe_prng_83_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_83 = {rand_exe_prng_83_io_out_15,rand_exe_prng_83_io_out_14,rand_exe_prng_83_io_out_13,
    rand_exe_prng_83_io_out_12,rand_exe_prng_83_io_out_11,rand_exe_prng_83_io_out_10,rand_exe_prng_83_io_out_9,
    rand_exe_prng_83_io_out_8,rand_exe_lo_83}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_84 = {rand_exe_prng_84_io_out_7,rand_exe_prng_84_io_out_6,rand_exe_prng_84_io_out_5,
    rand_exe_prng_84_io_out_4,rand_exe_prng_84_io_out_3,rand_exe_prng_84_io_out_2,rand_exe_prng_84_io_out_1,
    rand_exe_prng_84_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_84 = {rand_exe_prng_84_io_out_15,rand_exe_prng_84_io_out_14,rand_exe_prng_84_io_out_13,
    rand_exe_prng_84_io_out_12,rand_exe_prng_84_io_out_11,rand_exe_prng_84_io_out_10,rand_exe_prng_84_io_out_9,
    rand_exe_prng_84_io_out_8,rand_exe_lo_84}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_85 = {rand_exe_prng_85_io_out_7,rand_exe_prng_85_io_out_6,rand_exe_prng_85_io_out_5,
    rand_exe_prng_85_io_out_4,rand_exe_prng_85_io_out_3,rand_exe_prng_85_io_out_2,rand_exe_prng_85_io_out_1,
    rand_exe_prng_85_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_85 = {rand_exe_prng_85_io_out_15,rand_exe_prng_85_io_out_14,rand_exe_prng_85_io_out_13,
    rand_exe_prng_85_io_out_12,rand_exe_prng_85_io_out_11,rand_exe_prng_85_io_out_10,rand_exe_prng_85_io_out_9,
    rand_exe_prng_85_io_out_8,rand_exe_lo_85}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_86 = {rand_exe_prng_86_io_out_7,rand_exe_prng_86_io_out_6,rand_exe_prng_86_io_out_5,
    rand_exe_prng_86_io_out_4,rand_exe_prng_86_io_out_3,rand_exe_prng_86_io_out_2,rand_exe_prng_86_io_out_1,
    rand_exe_prng_86_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_86 = {rand_exe_prng_86_io_out_15,rand_exe_prng_86_io_out_14,rand_exe_prng_86_io_out_13,
    rand_exe_prng_86_io_out_12,rand_exe_prng_86_io_out_11,rand_exe_prng_86_io_out_10,rand_exe_prng_86_io_out_9,
    rand_exe_prng_86_io_out_8,rand_exe_lo_86}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_87 = {rand_exe_prng_87_io_out_7,rand_exe_prng_87_io_out_6,rand_exe_prng_87_io_out_5,
    rand_exe_prng_87_io_out_4,rand_exe_prng_87_io_out_3,rand_exe_prng_87_io_out_2,rand_exe_prng_87_io_out_1,
    rand_exe_prng_87_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_87 = {rand_exe_prng_87_io_out_15,rand_exe_prng_87_io_out_14,rand_exe_prng_87_io_out_13,
    rand_exe_prng_87_io_out_12,rand_exe_prng_87_io_out_11,rand_exe_prng_87_io_out_10,rand_exe_prng_87_io_out_9,
    rand_exe_prng_87_io_out_8,rand_exe_lo_87}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_88 = {rand_exe_prng_88_io_out_7,rand_exe_prng_88_io_out_6,rand_exe_prng_88_io_out_5,
    rand_exe_prng_88_io_out_4,rand_exe_prng_88_io_out_3,rand_exe_prng_88_io_out_2,rand_exe_prng_88_io_out_1,
    rand_exe_prng_88_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_88 = {rand_exe_prng_88_io_out_15,rand_exe_prng_88_io_out_14,rand_exe_prng_88_io_out_13,
    rand_exe_prng_88_io_out_12,rand_exe_prng_88_io_out_11,rand_exe_prng_88_io_out_10,rand_exe_prng_88_io_out_9,
    rand_exe_prng_88_io_out_8,rand_exe_lo_88}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_89 = {rand_exe_prng_89_io_out_7,rand_exe_prng_89_io_out_6,rand_exe_prng_89_io_out_5,
    rand_exe_prng_89_io_out_4,rand_exe_prng_89_io_out_3,rand_exe_prng_89_io_out_2,rand_exe_prng_89_io_out_1,
    rand_exe_prng_89_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_89 = {rand_exe_prng_89_io_out_15,rand_exe_prng_89_io_out_14,rand_exe_prng_89_io_out_13,
    rand_exe_prng_89_io_out_12,rand_exe_prng_89_io_out_11,rand_exe_prng_89_io_out_10,rand_exe_prng_89_io_out_9,
    rand_exe_prng_89_io_out_8,rand_exe_lo_89}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_90 = {rand_exe_prng_90_io_out_7,rand_exe_prng_90_io_out_6,rand_exe_prng_90_io_out_5,
    rand_exe_prng_90_io_out_4,rand_exe_prng_90_io_out_3,rand_exe_prng_90_io_out_2,rand_exe_prng_90_io_out_1,
    rand_exe_prng_90_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_90 = {rand_exe_prng_90_io_out_15,rand_exe_prng_90_io_out_14,rand_exe_prng_90_io_out_13,
    rand_exe_prng_90_io_out_12,rand_exe_prng_90_io_out_11,rand_exe_prng_90_io_out_10,rand_exe_prng_90_io_out_9,
    rand_exe_prng_90_io_out_8,rand_exe_lo_90}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_91 = {rand_exe_prng_91_io_out_7,rand_exe_prng_91_io_out_6,rand_exe_prng_91_io_out_5,
    rand_exe_prng_91_io_out_4,rand_exe_prng_91_io_out_3,rand_exe_prng_91_io_out_2,rand_exe_prng_91_io_out_1,
    rand_exe_prng_91_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_91 = {rand_exe_prng_91_io_out_15,rand_exe_prng_91_io_out_14,rand_exe_prng_91_io_out_13,
    rand_exe_prng_91_io_out_12,rand_exe_prng_91_io_out_11,rand_exe_prng_91_io_out_10,rand_exe_prng_91_io_out_9,
    rand_exe_prng_91_io_out_8,rand_exe_lo_91}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_92 = {rand_exe_prng_92_io_out_7,rand_exe_prng_92_io_out_6,rand_exe_prng_92_io_out_5,
    rand_exe_prng_92_io_out_4,rand_exe_prng_92_io_out_3,rand_exe_prng_92_io_out_2,rand_exe_prng_92_io_out_1,
    rand_exe_prng_92_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_92 = {rand_exe_prng_92_io_out_15,rand_exe_prng_92_io_out_14,rand_exe_prng_92_io_out_13,
    rand_exe_prng_92_io_out_12,rand_exe_prng_92_io_out_11,rand_exe_prng_92_io_out_10,rand_exe_prng_92_io_out_9,
    rand_exe_prng_92_io_out_8,rand_exe_lo_92}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_93 = {rand_exe_prng_93_io_out_7,rand_exe_prng_93_io_out_6,rand_exe_prng_93_io_out_5,
    rand_exe_prng_93_io_out_4,rand_exe_prng_93_io_out_3,rand_exe_prng_93_io_out_2,rand_exe_prng_93_io_out_1,
    rand_exe_prng_93_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_93 = {rand_exe_prng_93_io_out_15,rand_exe_prng_93_io_out_14,rand_exe_prng_93_io_out_13,
    rand_exe_prng_93_io_out_12,rand_exe_prng_93_io_out_11,rand_exe_prng_93_io_out_10,rand_exe_prng_93_io_out_9,
    rand_exe_prng_93_io_out_8,rand_exe_lo_93}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_94 = {rand_exe_prng_94_io_out_7,rand_exe_prng_94_io_out_6,rand_exe_prng_94_io_out_5,
    rand_exe_prng_94_io_out_4,rand_exe_prng_94_io_out_3,rand_exe_prng_94_io_out_2,rand_exe_prng_94_io_out_1,
    rand_exe_prng_94_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_94 = {rand_exe_prng_94_io_out_15,rand_exe_prng_94_io_out_14,rand_exe_prng_94_io_out_13,
    rand_exe_prng_94_io_out_12,rand_exe_prng_94_io_out_11,rand_exe_prng_94_io_out_10,rand_exe_prng_94_io_out_9,
    rand_exe_prng_94_io_out_8,rand_exe_lo_94}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_95 = {rand_exe_prng_95_io_out_7,rand_exe_prng_95_io_out_6,rand_exe_prng_95_io_out_5,
    rand_exe_prng_95_io_out_4,rand_exe_prng_95_io_out_3,rand_exe_prng_95_io_out_2,rand_exe_prng_95_io_out_1,
    rand_exe_prng_95_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_95 = {rand_exe_prng_95_io_out_15,rand_exe_prng_95_io_out_14,rand_exe_prng_95_io_out_13,
    rand_exe_prng_95_io_out_12,rand_exe_prng_95_io_out_11,rand_exe_prng_95_io_out_10,rand_exe_prng_95_io_out_9,
    rand_exe_prng_95_io_out_8,rand_exe_lo_95}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_96 = {rand_exe_prng_96_io_out_7,rand_exe_prng_96_io_out_6,rand_exe_prng_96_io_out_5,
    rand_exe_prng_96_io_out_4,rand_exe_prng_96_io_out_3,rand_exe_prng_96_io_out_2,rand_exe_prng_96_io_out_1,
    rand_exe_prng_96_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_96 = {rand_exe_prng_96_io_out_15,rand_exe_prng_96_io_out_14,rand_exe_prng_96_io_out_13,
    rand_exe_prng_96_io_out_12,rand_exe_prng_96_io_out_11,rand_exe_prng_96_io_out_10,rand_exe_prng_96_io_out_9,
    rand_exe_prng_96_io_out_8,rand_exe_lo_96}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_97 = {rand_exe_prng_97_io_out_7,rand_exe_prng_97_io_out_6,rand_exe_prng_97_io_out_5,
    rand_exe_prng_97_io_out_4,rand_exe_prng_97_io_out_3,rand_exe_prng_97_io_out_2,rand_exe_prng_97_io_out_1,
    rand_exe_prng_97_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_97 = {rand_exe_prng_97_io_out_15,rand_exe_prng_97_io_out_14,rand_exe_prng_97_io_out_13,
    rand_exe_prng_97_io_out_12,rand_exe_prng_97_io_out_11,rand_exe_prng_97_io_out_10,rand_exe_prng_97_io_out_9,
    rand_exe_prng_97_io_out_8,rand_exe_lo_97}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_98 = {rand_exe_prng_98_io_out_7,rand_exe_prng_98_io_out_6,rand_exe_prng_98_io_out_5,
    rand_exe_prng_98_io_out_4,rand_exe_prng_98_io_out_3,rand_exe_prng_98_io_out_2,rand_exe_prng_98_io_out_1,
    rand_exe_prng_98_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_98 = {rand_exe_prng_98_io_out_15,rand_exe_prng_98_io_out_14,rand_exe_prng_98_io_out_13,
    rand_exe_prng_98_io_out_12,rand_exe_prng_98_io_out_11,rand_exe_prng_98_io_out_10,rand_exe_prng_98_io_out_9,
    rand_exe_prng_98_io_out_8,rand_exe_lo_98}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_99 = {rand_exe_prng_99_io_out_7,rand_exe_prng_99_io_out_6,rand_exe_prng_99_io_out_5,
    rand_exe_prng_99_io_out_4,rand_exe_prng_99_io_out_3,rand_exe_prng_99_io_out_2,rand_exe_prng_99_io_out_1,
    rand_exe_prng_99_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_99 = {rand_exe_prng_99_io_out_15,rand_exe_prng_99_io_out_14,rand_exe_prng_99_io_out_13,
    rand_exe_prng_99_io_out_12,rand_exe_prng_99_io_out_11,rand_exe_prng_99_io_out_10,rand_exe_prng_99_io_out_9,
    rand_exe_prng_99_io_out_8,rand_exe_lo_99}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_100 = {rand_exe_prng_100_io_out_7,rand_exe_prng_100_io_out_6,rand_exe_prng_100_io_out_5,
    rand_exe_prng_100_io_out_4,rand_exe_prng_100_io_out_3,rand_exe_prng_100_io_out_2,rand_exe_prng_100_io_out_1,
    rand_exe_prng_100_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_100 = {rand_exe_prng_100_io_out_15,rand_exe_prng_100_io_out_14,rand_exe_prng_100_io_out_13,
    rand_exe_prng_100_io_out_12,rand_exe_prng_100_io_out_11,rand_exe_prng_100_io_out_10,rand_exe_prng_100_io_out_9,
    rand_exe_prng_100_io_out_8,rand_exe_lo_100}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_101 = {rand_exe_prng_101_io_out_7,rand_exe_prng_101_io_out_6,rand_exe_prng_101_io_out_5,
    rand_exe_prng_101_io_out_4,rand_exe_prng_101_io_out_3,rand_exe_prng_101_io_out_2,rand_exe_prng_101_io_out_1,
    rand_exe_prng_101_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_101 = {rand_exe_prng_101_io_out_15,rand_exe_prng_101_io_out_14,rand_exe_prng_101_io_out_13,
    rand_exe_prng_101_io_out_12,rand_exe_prng_101_io_out_11,rand_exe_prng_101_io_out_10,rand_exe_prng_101_io_out_9,
    rand_exe_prng_101_io_out_8,rand_exe_lo_101}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_102 = {rand_exe_prng_102_io_out_7,rand_exe_prng_102_io_out_6,rand_exe_prng_102_io_out_5,
    rand_exe_prng_102_io_out_4,rand_exe_prng_102_io_out_3,rand_exe_prng_102_io_out_2,rand_exe_prng_102_io_out_1,
    rand_exe_prng_102_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_102 = {rand_exe_prng_102_io_out_15,rand_exe_prng_102_io_out_14,rand_exe_prng_102_io_out_13,
    rand_exe_prng_102_io_out_12,rand_exe_prng_102_io_out_11,rand_exe_prng_102_io_out_10,rand_exe_prng_102_io_out_9,
    rand_exe_prng_102_io_out_8,rand_exe_lo_102}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_103 = {rand_exe_prng_103_io_out_7,rand_exe_prng_103_io_out_6,rand_exe_prng_103_io_out_5,
    rand_exe_prng_103_io_out_4,rand_exe_prng_103_io_out_3,rand_exe_prng_103_io_out_2,rand_exe_prng_103_io_out_1,
    rand_exe_prng_103_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_103 = {rand_exe_prng_103_io_out_15,rand_exe_prng_103_io_out_14,rand_exe_prng_103_io_out_13,
    rand_exe_prng_103_io_out_12,rand_exe_prng_103_io_out_11,rand_exe_prng_103_io_out_10,rand_exe_prng_103_io_out_9,
    rand_exe_prng_103_io_out_8,rand_exe_lo_103}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_104 = {rand_exe_prng_104_io_out_7,rand_exe_prng_104_io_out_6,rand_exe_prng_104_io_out_5,
    rand_exe_prng_104_io_out_4,rand_exe_prng_104_io_out_3,rand_exe_prng_104_io_out_2,rand_exe_prng_104_io_out_1,
    rand_exe_prng_104_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_104 = {rand_exe_prng_104_io_out_15,rand_exe_prng_104_io_out_14,rand_exe_prng_104_io_out_13,
    rand_exe_prng_104_io_out_12,rand_exe_prng_104_io_out_11,rand_exe_prng_104_io_out_10,rand_exe_prng_104_io_out_9,
    rand_exe_prng_104_io_out_8,rand_exe_lo_104}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_105 = {rand_exe_prng_105_io_out_7,rand_exe_prng_105_io_out_6,rand_exe_prng_105_io_out_5,
    rand_exe_prng_105_io_out_4,rand_exe_prng_105_io_out_3,rand_exe_prng_105_io_out_2,rand_exe_prng_105_io_out_1,
    rand_exe_prng_105_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_105 = {rand_exe_prng_105_io_out_15,rand_exe_prng_105_io_out_14,rand_exe_prng_105_io_out_13,
    rand_exe_prng_105_io_out_12,rand_exe_prng_105_io_out_11,rand_exe_prng_105_io_out_10,rand_exe_prng_105_io_out_9,
    rand_exe_prng_105_io_out_8,rand_exe_lo_105}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_106 = {rand_exe_prng_106_io_out_7,rand_exe_prng_106_io_out_6,rand_exe_prng_106_io_out_5,
    rand_exe_prng_106_io_out_4,rand_exe_prng_106_io_out_3,rand_exe_prng_106_io_out_2,rand_exe_prng_106_io_out_1,
    rand_exe_prng_106_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_106 = {rand_exe_prng_106_io_out_15,rand_exe_prng_106_io_out_14,rand_exe_prng_106_io_out_13,
    rand_exe_prng_106_io_out_12,rand_exe_prng_106_io_out_11,rand_exe_prng_106_io_out_10,rand_exe_prng_106_io_out_9,
    rand_exe_prng_106_io_out_8,rand_exe_lo_106}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_107 = {rand_exe_prng_107_io_out_7,rand_exe_prng_107_io_out_6,rand_exe_prng_107_io_out_5,
    rand_exe_prng_107_io_out_4,rand_exe_prng_107_io_out_3,rand_exe_prng_107_io_out_2,rand_exe_prng_107_io_out_1,
    rand_exe_prng_107_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_107 = {rand_exe_prng_107_io_out_15,rand_exe_prng_107_io_out_14,rand_exe_prng_107_io_out_13,
    rand_exe_prng_107_io_out_12,rand_exe_prng_107_io_out_11,rand_exe_prng_107_io_out_10,rand_exe_prng_107_io_out_9,
    rand_exe_prng_107_io_out_8,rand_exe_lo_107}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_108 = {rand_exe_prng_108_io_out_7,rand_exe_prng_108_io_out_6,rand_exe_prng_108_io_out_5,
    rand_exe_prng_108_io_out_4,rand_exe_prng_108_io_out_3,rand_exe_prng_108_io_out_2,rand_exe_prng_108_io_out_1,
    rand_exe_prng_108_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_108 = {rand_exe_prng_108_io_out_15,rand_exe_prng_108_io_out_14,rand_exe_prng_108_io_out_13,
    rand_exe_prng_108_io_out_12,rand_exe_prng_108_io_out_11,rand_exe_prng_108_io_out_10,rand_exe_prng_108_io_out_9,
    rand_exe_prng_108_io_out_8,rand_exe_lo_108}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_109 = {rand_exe_prng_109_io_out_7,rand_exe_prng_109_io_out_6,rand_exe_prng_109_io_out_5,
    rand_exe_prng_109_io_out_4,rand_exe_prng_109_io_out_3,rand_exe_prng_109_io_out_2,rand_exe_prng_109_io_out_1,
    rand_exe_prng_109_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_109 = {rand_exe_prng_109_io_out_15,rand_exe_prng_109_io_out_14,rand_exe_prng_109_io_out_13,
    rand_exe_prng_109_io_out_12,rand_exe_prng_109_io_out_11,rand_exe_prng_109_io_out_10,rand_exe_prng_109_io_out_9,
    rand_exe_prng_109_io_out_8,rand_exe_lo_109}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_110 = {rand_exe_prng_110_io_out_7,rand_exe_prng_110_io_out_6,rand_exe_prng_110_io_out_5,
    rand_exe_prng_110_io_out_4,rand_exe_prng_110_io_out_3,rand_exe_prng_110_io_out_2,rand_exe_prng_110_io_out_1,
    rand_exe_prng_110_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_110 = {rand_exe_prng_110_io_out_15,rand_exe_prng_110_io_out_14,rand_exe_prng_110_io_out_13,
    rand_exe_prng_110_io_out_12,rand_exe_prng_110_io_out_11,rand_exe_prng_110_io_out_10,rand_exe_prng_110_io_out_9,
    rand_exe_prng_110_io_out_8,rand_exe_lo_110}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_111 = {rand_exe_prng_111_io_out_7,rand_exe_prng_111_io_out_6,rand_exe_prng_111_io_out_5,
    rand_exe_prng_111_io_out_4,rand_exe_prng_111_io_out_3,rand_exe_prng_111_io_out_2,rand_exe_prng_111_io_out_1,
    rand_exe_prng_111_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_111 = {rand_exe_prng_111_io_out_15,rand_exe_prng_111_io_out_14,rand_exe_prng_111_io_out_13,
    rand_exe_prng_111_io_out_12,rand_exe_prng_111_io_out_11,rand_exe_prng_111_io_out_10,rand_exe_prng_111_io_out_9,
    rand_exe_prng_111_io_out_8,rand_exe_lo_111}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_112 = {rand_exe_prng_112_io_out_7,rand_exe_prng_112_io_out_6,rand_exe_prng_112_io_out_5,
    rand_exe_prng_112_io_out_4,rand_exe_prng_112_io_out_3,rand_exe_prng_112_io_out_2,rand_exe_prng_112_io_out_1,
    rand_exe_prng_112_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_112 = {rand_exe_prng_112_io_out_15,rand_exe_prng_112_io_out_14,rand_exe_prng_112_io_out_13,
    rand_exe_prng_112_io_out_12,rand_exe_prng_112_io_out_11,rand_exe_prng_112_io_out_10,rand_exe_prng_112_io_out_9,
    rand_exe_prng_112_io_out_8,rand_exe_lo_112}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_113 = {rand_exe_prng_113_io_out_7,rand_exe_prng_113_io_out_6,rand_exe_prng_113_io_out_5,
    rand_exe_prng_113_io_out_4,rand_exe_prng_113_io_out_3,rand_exe_prng_113_io_out_2,rand_exe_prng_113_io_out_1,
    rand_exe_prng_113_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_113 = {rand_exe_prng_113_io_out_15,rand_exe_prng_113_io_out_14,rand_exe_prng_113_io_out_13,
    rand_exe_prng_113_io_out_12,rand_exe_prng_113_io_out_11,rand_exe_prng_113_io_out_10,rand_exe_prng_113_io_out_9,
    rand_exe_prng_113_io_out_8,rand_exe_lo_113}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_114 = {rand_exe_prng_114_io_out_7,rand_exe_prng_114_io_out_6,rand_exe_prng_114_io_out_5,
    rand_exe_prng_114_io_out_4,rand_exe_prng_114_io_out_3,rand_exe_prng_114_io_out_2,rand_exe_prng_114_io_out_1,
    rand_exe_prng_114_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_114 = {rand_exe_prng_114_io_out_15,rand_exe_prng_114_io_out_14,rand_exe_prng_114_io_out_13,
    rand_exe_prng_114_io_out_12,rand_exe_prng_114_io_out_11,rand_exe_prng_114_io_out_10,rand_exe_prng_114_io_out_9,
    rand_exe_prng_114_io_out_8,rand_exe_lo_114}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_115 = {rand_exe_prng_115_io_out_7,rand_exe_prng_115_io_out_6,rand_exe_prng_115_io_out_5,
    rand_exe_prng_115_io_out_4,rand_exe_prng_115_io_out_3,rand_exe_prng_115_io_out_2,rand_exe_prng_115_io_out_1,
    rand_exe_prng_115_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_115 = {rand_exe_prng_115_io_out_15,rand_exe_prng_115_io_out_14,rand_exe_prng_115_io_out_13,
    rand_exe_prng_115_io_out_12,rand_exe_prng_115_io_out_11,rand_exe_prng_115_io_out_10,rand_exe_prng_115_io_out_9,
    rand_exe_prng_115_io_out_8,rand_exe_lo_115}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_116 = {rand_exe_prng_116_io_out_7,rand_exe_prng_116_io_out_6,rand_exe_prng_116_io_out_5,
    rand_exe_prng_116_io_out_4,rand_exe_prng_116_io_out_3,rand_exe_prng_116_io_out_2,rand_exe_prng_116_io_out_1,
    rand_exe_prng_116_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_116 = {rand_exe_prng_116_io_out_15,rand_exe_prng_116_io_out_14,rand_exe_prng_116_io_out_13,
    rand_exe_prng_116_io_out_12,rand_exe_prng_116_io_out_11,rand_exe_prng_116_io_out_10,rand_exe_prng_116_io_out_9,
    rand_exe_prng_116_io_out_8,rand_exe_lo_116}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_117 = {rand_exe_prng_117_io_out_7,rand_exe_prng_117_io_out_6,rand_exe_prng_117_io_out_5,
    rand_exe_prng_117_io_out_4,rand_exe_prng_117_io_out_3,rand_exe_prng_117_io_out_2,rand_exe_prng_117_io_out_1,
    rand_exe_prng_117_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_117 = {rand_exe_prng_117_io_out_15,rand_exe_prng_117_io_out_14,rand_exe_prng_117_io_out_13,
    rand_exe_prng_117_io_out_12,rand_exe_prng_117_io_out_11,rand_exe_prng_117_io_out_10,rand_exe_prng_117_io_out_9,
    rand_exe_prng_117_io_out_8,rand_exe_lo_117}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_118 = {rand_exe_prng_118_io_out_7,rand_exe_prng_118_io_out_6,rand_exe_prng_118_io_out_5,
    rand_exe_prng_118_io_out_4,rand_exe_prng_118_io_out_3,rand_exe_prng_118_io_out_2,rand_exe_prng_118_io_out_1,
    rand_exe_prng_118_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_118 = {rand_exe_prng_118_io_out_15,rand_exe_prng_118_io_out_14,rand_exe_prng_118_io_out_13,
    rand_exe_prng_118_io_out_12,rand_exe_prng_118_io_out_11,rand_exe_prng_118_io_out_10,rand_exe_prng_118_io_out_9,
    rand_exe_prng_118_io_out_8,rand_exe_lo_118}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_119 = {rand_exe_prng_119_io_out_7,rand_exe_prng_119_io_out_6,rand_exe_prng_119_io_out_5,
    rand_exe_prng_119_io_out_4,rand_exe_prng_119_io_out_3,rand_exe_prng_119_io_out_2,rand_exe_prng_119_io_out_1,
    rand_exe_prng_119_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_119 = {rand_exe_prng_119_io_out_15,rand_exe_prng_119_io_out_14,rand_exe_prng_119_io_out_13,
    rand_exe_prng_119_io_out_12,rand_exe_prng_119_io_out_11,rand_exe_prng_119_io_out_10,rand_exe_prng_119_io_out_9,
    rand_exe_prng_119_io_out_8,rand_exe_lo_119}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_120 = {rand_exe_prng_120_io_out_7,rand_exe_prng_120_io_out_6,rand_exe_prng_120_io_out_5,
    rand_exe_prng_120_io_out_4,rand_exe_prng_120_io_out_3,rand_exe_prng_120_io_out_2,rand_exe_prng_120_io_out_1,
    rand_exe_prng_120_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_120 = {rand_exe_prng_120_io_out_15,rand_exe_prng_120_io_out_14,rand_exe_prng_120_io_out_13,
    rand_exe_prng_120_io_out_12,rand_exe_prng_120_io_out_11,rand_exe_prng_120_io_out_10,rand_exe_prng_120_io_out_9,
    rand_exe_prng_120_io_out_8,rand_exe_lo_120}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_121 = {rand_exe_prng_121_io_out_7,rand_exe_prng_121_io_out_6,rand_exe_prng_121_io_out_5,
    rand_exe_prng_121_io_out_4,rand_exe_prng_121_io_out_3,rand_exe_prng_121_io_out_2,rand_exe_prng_121_io_out_1,
    rand_exe_prng_121_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_121 = {rand_exe_prng_121_io_out_15,rand_exe_prng_121_io_out_14,rand_exe_prng_121_io_out_13,
    rand_exe_prng_121_io_out_12,rand_exe_prng_121_io_out_11,rand_exe_prng_121_io_out_10,rand_exe_prng_121_io_out_9,
    rand_exe_prng_121_io_out_8,rand_exe_lo_121}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_122 = {rand_exe_prng_122_io_out_7,rand_exe_prng_122_io_out_6,rand_exe_prng_122_io_out_5,
    rand_exe_prng_122_io_out_4,rand_exe_prng_122_io_out_3,rand_exe_prng_122_io_out_2,rand_exe_prng_122_io_out_1,
    rand_exe_prng_122_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_122 = {rand_exe_prng_122_io_out_15,rand_exe_prng_122_io_out_14,rand_exe_prng_122_io_out_13,
    rand_exe_prng_122_io_out_12,rand_exe_prng_122_io_out_11,rand_exe_prng_122_io_out_10,rand_exe_prng_122_io_out_9,
    rand_exe_prng_122_io_out_8,rand_exe_lo_122}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_123 = {rand_exe_prng_123_io_out_7,rand_exe_prng_123_io_out_6,rand_exe_prng_123_io_out_5,
    rand_exe_prng_123_io_out_4,rand_exe_prng_123_io_out_3,rand_exe_prng_123_io_out_2,rand_exe_prng_123_io_out_1,
    rand_exe_prng_123_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_123 = {rand_exe_prng_123_io_out_15,rand_exe_prng_123_io_out_14,rand_exe_prng_123_io_out_13,
    rand_exe_prng_123_io_out_12,rand_exe_prng_123_io_out_11,rand_exe_prng_123_io_out_10,rand_exe_prng_123_io_out_9,
    rand_exe_prng_123_io_out_8,rand_exe_lo_123}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_124 = {rand_exe_prng_124_io_out_7,rand_exe_prng_124_io_out_6,rand_exe_prng_124_io_out_5,
    rand_exe_prng_124_io_out_4,rand_exe_prng_124_io_out_3,rand_exe_prng_124_io_out_2,rand_exe_prng_124_io_out_1,
    rand_exe_prng_124_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_124 = {rand_exe_prng_124_io_out_15,rand_exe_prng_124_io_out_14,rand_exe_prng_124_io_out_13,
    rand_exe_prng_124_io_out_12,rand_exe_prng_124_io_out_11,rand_exe_prng_124_io_out_10,rand_exe_prng_124_io_out_9,
    rand_exe_prng_124_io_out_8,rand_exe_lo_124}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_125 = {rand_exe_prng_125_io_out_7,rand_exe_prng_125_io_out_6,rand_exe_prng_125_io_out_5,
    rand_exe_prng_125_io_out_4,rand_exe_prng_125_io_out_3,rand_exe_prng_125_io_out_2,rand_exe_prng_125_io_out_1,
    rand_exe_prng_125_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_125 = {rand_exe_prng_125_io_out_15,rand_exe_prng_125_io_out_14,rand_exe_prng_125_io_out_13,
    rand_exe_prng_125_io_out_12,rand_exe_prng_125_io_out_11,rand_exe_prng_125_io_out_10,rand_exe_prng_125_io_out_9,
    rand_exe_prng_125_io_out_8,rand_exe_lo_125}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_126 = {rand_exe_prng_126_io_out_7,rand_exe_prng_126_io_out_6,rand_exe_prng_126_io_out_5,
    rand_exe_prng_126_io_out_4,rand_exe_prng_126_io_out_3,rand_exe_prng_126_io_out_2,rand_exe_prng_126_io_out_1,
    rand_exe_prng_126_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_126 = {rand_exe_prng_126_io_out_15,rand_exe_prng_126_io_out_14,rand_exe_prng_126_io_out_13,
    rand_exe_prng_126_io_out_12,rand_exe_prng_126_io_out_11,rand_exe_prng_126_io_out_10,rand_exe_prng_126_io_out_9,
    rand_exe_prng_126_io_out_8,rand_exe_lo_126}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_127 = {rand_exe_prng_127_io_out_7,rand_exe_prng_127_io_out_6,rand_exe_prng_127_io_out_5,
    rand_exe_prng_127_io_out_4,rand_exe_prng_127_io_out_3,rand_exe_prng_127_io_out_2,rand_exe_prng_127_io_out_1,
    rand_exe_prng_127_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_127 = {rand_exe_prng_127_io_out_15,rand_exe_prng_127_io_out_14,rand_exe_prng_127_io_out_13,
    rand_exe_prng_127_io_out_12,rand_exe_prng_127_io_out_11,rand_exe_prng_127_io_out_10,rand_exe_prng_127_io_out_9,
    rand_exe_prng_127_io_out_8,rand_exe_lo_127}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_128 = {rand_exe_prng_128_io_out_7,rand_exe_prng_128_io_out_6,rand_exe_prng_128_io_out_5,
    rand_exe_prng_128_io_out_4,rand_exe_prng_128_io_out_3,rand_exe_prng_128_io_out_2,rand_exe_prng_128_io_out_1,
    rand_exe_prng_128_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_128 = {rand_exe_prng_128_io_out_15,rand_exe_prng_128_io_out_14,rand_exe_prng_128_io_out_13,
    rand_exe_prng_128_io_out_12,rand_exe_prng_128_io_out_11,rand_exe_prng_128_io_out_10,rand_exe_prng_128_io_out_9,
    rand_exe_prng_128_io_out_8,rand_exe_lo_128}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_129 = {rand_exe_prng_129_io_out_7,rand_exe_prng_129_io_out_6,rand_exe_prng_129_io_out_5,
    rand_exe_prng_129_io_out_4,rand_exe_prng_129_io_out_3,rand_exe_prng_129_io_out_2,rand_exe_prng_129_io_out_1,
    rand_exe_prng_129_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_129 = {rand_exe_prng_129_io_out_15,rand_exe_prng_129_io_out_14,rand_exe_prng_129_io_out_13,
    rand_exe_prng_129_io_out_12,rand_exe_prng_129_io_out_11,rand_exe_prng_129_io_out_10,rand_exe_prng_129_io_out_9,
    rand_exe_prng_129_io_out_8,rand_exe_lo_129}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_130 = {rand_exe_prng_130_io_out_7,rand_exe_prng_130_io_out_6,rand_exe_prng_130_io_out_5,
    rand_exe_prng_130_io_out_4,rand_exe_prng_130_io_out_3,rand_exe_prng_130_io_out_2,rand_exe_prng_130_io_out_1,
    rand_exe_prng_130_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_130 = {rand_exe_prng_130_io_out_15,rand_exe_prng_130_io_out_14,rand_exe_prng_130_io_out_13,
    rand_exe_prng_130_io_out_12,rand_exe_prng_130_io_out_11,rand_exe_prng_130_io_out_10,rand_exe_prng_130_io_out_9,
    rand_exe_prng_130_io_out_8,rand_exe_lo_130}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_131 = {rand_exe_prng_131_io_out_7,rand_exe_prng_131_io_out_6,rand_exe_prng_131_io_out_5,
    rand_exe_prng_131_io_out_4,rand_exe_prng_131_io_out_3,rand_exe_prng_131_io_out_2,rand_exe_prng_131_io_out_1,
    rand_exe_prng_131_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_131 = {rand_exe_prng_131_io_out_15,rand_exe_prng_131_io_out_14,rand_exe_prng_131_io_out_13,
    rand_exe_prng_131_io_out_12,rand_exe_prng_131_io_out_11,rand_exe_prng_131_io_out_10,rand_exe_prng_131_io_out_9,
    rand_exe_prng_131_io_out_8,rand_exe_lo_131}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_132 = {rand_exe_prng_132_io_out_7,rand_exe_prng_132_io_out_6,rand_exe_prng_132_io_out_5,
    rand_exe_prng_132_io_out_4,rand_exe_prng_132_io_out_3,rand_exe_prng_132_io_out_2,rand_exe_prng_132_io_out_1,
    rand_exe_prng_132_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_132 = {rand_exe_prng_132_io_out_15,rand_exe_prng_132_io_out_14,rand_exe_prng_132_io_out_13,
    rand_exe_prng_132_io_out_12,rand_exe_prng_132_io_out_11,rand_exe_prng_132_io_out_10,rand_exe_prng_132_io_out_9,
    rand_exe_prng_132_io_out_8,rand_exe_lo_132}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_133 = {rand_exe_prng_133_io_out_7,rand_exe_prng_133_io_out_6,rand_exe_prng_133_io_out_5,
    rand_exe_prng_133_io_out_4,rand_exe_prng_133_io_out_3,rand_exe_prng_133_io_out_2,rand_exe_prng_133_io_out_1,
    rand_exe_prng_133_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_133 = {rand_exe_prng_133_io_out_15,rand_exe_prng_133_io_out_14,rand_exe_prng_133_io_out_13,
    rand_exe_prng_133_io_out_12,rand_exe_prng_133_io_out_11,rand_exe_prng_133_io_out_10,rand_exe_prng_133_io_out_9,
    rand_exe_prng_133_io_out_8,rand_exe_lo_133}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_134 = {rand_exe_prng_134_io_out_7,rand_exe_prng_134_io_out_6,rand_exe_prng_134_io_out_5,
    rand_exe_prng_134_io_out_4,rand_exe_prng_134_io_out_3,rand_exe_prng_134_io_out_2,rand_exe_prng_134_io_out_1,
    rand_exe_prng_134_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_134 = {rand_exe_prng_134_io_out_15,rand_exe_prng_134_io_out_14,rand_exe_prng_134_io_out_13,
    rand_exe_prng_134_io_out_12,rand_exe_prng_134_io_out_11,rand_exe_prng_134_io_out_10,rand_exe_prng_134_io_out_9,
    rand_exe_prng_134_io_out_8,rand_exe_lo_134}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_135 = {rand_exe_prng_135_io_out_7,rand_exe_prng_135_io_out_6,rand_exe_prng_135_io_out_5,
    rand_exe_prng_135_io_out_4,rand_exe_prng_135_io_out_3,rand_exe_prng_135_io_out_2,rand_exe_prng_135_io_out_1,
    rand_exe_prng_135_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_135 = {rand_exe_prng_135_io_out_15,rand_exe_prng_135_io_out_14,rand_exe_prng_135_io_out_13,
    rand_exe_prng_135_io_out_12,rand_exe_prng_135_io_out_11,rand_exe_prng_135_io_out_10,rand_exe_prng_135_io_out_9,
    rand_exe_prng_135_io_out_8,rand_exe_lo_135}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_136 = {rand_exe_prng_136_io_out_7,rand_exe_prng_136_io_out_6,rand_exe_prng_136_io_out_5,
    rand_exe_prng_136_io_out_4,rand_exe_prng_136_io_out_3,rand_exe_prng_136_io_out_2,rand_exe_prng_136_io_out_1,
    rand_exe_prng_136_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_136 = {rand_exe_prng_136_io_out_15,rand_exe_prng_136_io_out_14,rand_exe_prng_136_io_out_13,
    rand_exe_prng_136_io_out_12,rand_exe_prng_136_io_out_11,rand_exe_prng_136_io_out_10,rand_exe_prng_136_io_out_9,
    rand_exe_prng_136_io_out_8,rand_exe_lo_136}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_137 = {rand_exe_prng_137_io_out_7,rand_exe_prng_137_io_out_6,rand_exe_prng_137_io_out_5,
    rand_exe_prng_137_io_out_4,rand_exe_prng_137_io_out_3,rand_exe_prng_137_io_out_2,rand_exe_prng_137_io_out_1,
    rand_exe_prng_137_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_137 = {rand_exe_prng_137_io_out_15,rand_exe_prng_137_io_out_14,rand_exe_prng_137_io_out_13,
    rand_exe_prng_137_io_out_12,rand_exe_prng_137_io_out_11,rand_exe_prng_137_io_out_10,rand_exe_prng_137_io_out_9,
    rand_exe_prng_137_io_out_8,rand_exe_lo_137}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_138 = {rand_exe_prng_138_io_out_7,rand_exe_prng_138_io_out_6,rand_exe_prng_138_io_out_5,
    rand_exe_prng_138_io_out_4,rand_exe_prng_138_io_out_3,rand_exe_prng_138_io_out_2,rand_exe_prng_138_io_out_1,
    rand_exe_prng_138_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_138 = {rand_exe_prng_138_io_out_15,rand_exe_prng_138_io_out_14,rand_exe_prng_138_io_out_13,
    rand_exe_prng_138_io_out_12,rand_exe_prng_138_io_out_11,rand_exe_prng_138_io_out_10,rand_exe_prng_138_io_out_9,
    rand_exe_prng_138_io_out_8,rand_exe_lo_138}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_139 = {rand_exe_prng_139_io_out_7,rand_exe_prng_139_io_out_6,rand_exe_prng_139_io_out_5,
    rand_exe_prng_139_io_out_4,rand_exe_prng_139_io_out_3,rand_exe_prng_139_io_out_2,rand_exe_prng_139_io_out_1,
    rand_exe_prng_139_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_139 = {rand_exe_prng_139_io_out_15,rand_exe_prng_139_io_out_14,rand_exe_prng_139_io_out_13,
    rand_exe_prng_139_io_out_12,rand_exe_prng_139_io_out_11,rand_exe_prng_139_io_out_10,rand_exe_prng_139_io_out_9,
    rand_exe_prng_139_io_out_8,rand_exe_lo_139}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_140 = {rand_exe_prng_140_io_out_7,rand_exe_prng_140_io_out_6,rand_exe_prng_140_io_out_5,
    rand_exe_prng_140_io_out_4,rand_exe_prng_140_io_out_3,rand_exe_prng_140_io_out_2,rand_exe_prng_140_io_out_1,
    rand_exe_prng_140_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_140 = {rand_exe_prng_140_io_out_15,rand_exe_prng_140_io_out_14,rand_exe_prng_140_io_out_13,
    rand_exe_prng_140_io_out_12,rand_exe_prng_140_io_out_11,rand_exe_prng_140_io_out_10,rand_exe_prng_140_io_out_9,
    rand_exe_prng_140_io_out_8,rand_exe_lo_140}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_141 = {rand_exe_prng_141_io_out_7,rand_exe_prng_141_io_out_6,rand_exe_prng_141_io_out_5,
    rand_exe_prng_141_io_out_4,rand_exe_prng_141_io_out_3,rand_exe_prng_141_io_out_2,rand_exe_prng_141_io_out_1,
    rand_exe_prng_141_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_141 = {rand_exe_prng_141_io_out_15,rand_exe_prng_141_io_out_14,rand_exe_prng_141_io_out_13,
    rand_exe_prng_141_io_out_12,rand_exe_prng_141_io_out_11,rand_exe_prng_141_io_out_10,rand_exe_prng_141_io_out_9,
    rand_exe_prng_141_io_out_8,rand_exe_lo_141}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_142 = {rand_exe_prng_142_io_out_7,rand_exe_prng_142_io_out_6,rand_exe_prng_142_io_out_5,
    rand_exe_prng_142_io_out_4,rand_exe_prng_142_io_out_3,rand_exe_prng_142_io_out_2,rand_exe_prng_142_io_out_1,
    rand_exe_prng_142_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_142 = {rand_exe_prng_142_io_out_15,rand_exe_prng_142_io_out_14,rand_exe_prng_142_io_out_13,
    rand_exe_prng_142_io_out_12,rand_exe_prng_142_io_out_11,rand_exe_prng_142_io_out_10,rand_exe_prng_142_io_out_9,
    rand_exe_prng_142_io_out_8,rand_exe_lo_142}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_143 = {rand_exe_prng_143_io_out_7,rand_exe_prng_143_io_out_6,rand_exe_prng_143_io_out_5,
    rand_exe_prng_143_io_out_4,rand_exe_prng_143_io_out_3,rand_exe_prng_143_io_out_2,rand_exe_prng_143_io_out_1,
    rand_exe_prng_143_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_143 = {rand_exe_prng_143_io_out_15,rand_exe_prng_143_io_out_14,rand_exe_prng_143_io_out_13,
    rand_exe_prng_143_io_out_12,rand_exe_prng_143_io_out_11,rand_exe_prng_143_io_out_10,rand_exe_prng_143_io_out_9,
    rand_exe_prng_143_io_out_8,rand_exe_lo_143}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_144 = {rand_exe_prng_144_io_out_7,rand_exe_prng_144_io_out_6,rand_exe_prng_144_io_out_5,
    rand_exe_prng_144_io_out_4,rand_exe_prng_144_io_out_3,rand_exe_prng_144_io_out_2,rand_exe_prng_144_io_out_1,
    rand_exe_prng_144_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_144 = {rand_exe_prng_144_io_out_15,rand_exe_prng_144_io_out_14,rand_exe_prng_144_io_out_13,
    rand_exe_prng_144_io_out_12,rand_exe_prng_144_io_out_11,rand_exe_prng_144_io_out_10,rand_exe_prng_144_io_out_9,
    rand_exe_prng_144_io_out_8,rand_exe_lo_144}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_145 = {rand_exe_prng_145_io_out_7,rand_exe_prng_145_io_out_6,rand_exe_prng_145_io_out_5,
    rand_exe_prng_145_io_out_4,rand_exe_prng_145_io_out_3,rand_exe_prng_145_io_out_2,rand_exe_prng_145_io_out_1,
    rand_exe_prng_145_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_145 = {rand_exe_prng_145_io_out_15,rand_exe_prng_145_io_out_14,rand_exe_prng_145_io_out_13,
    rand_exe_prng_145_io_out_12,rand_exe_prng_145_io_out_11,rand_exe_prng_145_io_out_10,rand_exe_prng_145_io_out_9,
    rand_exe_prng_145_io_out_8,rand_exe_lo_145}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_146 = {rand_exe_prng_146_io_out_7,rand_exe_prng_146_io_out_6,rand_exe_prng_146_io_out_5,
    rand_exe_prng_146_io_out_4,rand_exe_prng_146_io_out_3,rand_exe_prng_146_io_out_2,rand_exe_prng_146_io_out_1,
    rand_exe_prng_146_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_146 = {rand_exe_prng_146_io_out_15,rand_exe_prng_146_io_out_14,rand_exe_prng_146_io_out_13,
    rand_exe_prng_146_io_out_12,rand_exe_prng_146_io_out_11,rand_exe_prng_146_io_out_10,rand_exe_prng_146_io_out_9,
    rand_exe_prng_146_io_out_8,rand_exe_lo_146}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_147 = {rand_exe_prng_147_io_out_7,rand_exe_prng_147_io_out_6,rand_exe_prng_147_io_out_5,
    rand_exe_prng_147_io_out_4,rand_exe_prng_147_io_out_3,rand_exe_prng_147_io_out_2,rand_exe_prng_147_io_out_1,
    rand_exe_prng_147_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_147 = {rand_exe_prng_147_io_out_15,rand_exe_prng_147_io_out_14,rand_exe_prng_147_io_out_13,
    rand_exe_prng_147_io_out_12,rand_exe_prng_147_io_out_11,rand_exe_prng_147_io_out_10,rand_exe_prng_147_io_out_9,
    rand_exe_prng_147_io_out_8,rand_exe_lo_147}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_148 = {rand_exe_prng_148_io_out_7,rand_exe_prng_148_io_out_6,rand_exe_prng_148_io_out_5,
    rand_exe_prng_148_io_out_4,rand_exe_prng_148_io_out_3,rand_exe_prng_148_io_out_2,rand_exe_prng_148_io_out_1,
    rand_exe_prng_148_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_148 = {rand_exe_prng_148_io_out_15,rand_exe_prng_148_io_out_14,rand_exe_prng_148_io_out_13,
    rand_exe_prng_148_io_out_12,rand_exe_prng_148_io_out_11,rand_exe_prng_148_io_out_10,rand_exe_prng_148_io_out_9,
    rand_exe_prng_148_io_out_8,rand_exe_lo_148}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_149 = {rand_exe_prng_149_io_out_7,rand_exe_prng_149_io_out_6,rand_exe_prng_149_io_out_5,
    rand_exe_prng_149_io_out_4,rand_exe_prng_149_io_out_3,rand_exe_prng_149_io_out_2,rand_exe_prng_149_io_out_1,
    rand_exe_prng_149_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_149 = {rand_exe_prng_149_io_out_15,rand_exe_prng_149_io_out_14,rand_exe_prng_149_io_out_13,
    rand_exe_prng_149_io_out_12,rand_exe_prng_149_io_out_11,rand_exe_prng_149_io_out_10,rand_exe_prng_149_io_out_9,
    rand_exe_prng_149_io_out_8,rand_exe_lo_149}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_150 = {rand_exe_prng_150_io_out_7,rand_exe_prng_150_io_out_6,rand_exe_prng_150_io_out_5,
    rand_exe_prng_150_io_out_4,rand_exe_prng_150_io_out_3,rand_exe_prng_150_io_out_2,rand_exe_prng_150_io_out_1,
    rand_exe_prng_150_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_150 = {rand_exe_prng_150_io_out_15,rand_exe_prng_150_io_out_14,rand_exe_prng_150_io_out_13,
    rand_exe_prng_150_io_out_12,rand_exe_prng_150_io_out_11,rand_exe_prng_150_io_out_10,rand_exe_prng_150_io_out_9,
    rand_exe_prng_150_io_out_8,rand_exe_lo_150}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_151 = {rand_exe_prng_151_io_out_7,rand_exe_prng_151_io_out_6,rand_exe_prng_151_io_out_5,
    rand_exe_prng_151_io_out_4,rand_exe_prng_151_io_out_3,rand_exe_prng_151_io_out_2,rand_exe_prng_151_io_out_1,
    rand_exe_prng_151_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_151 = {rand_exe_prng_151_io_out_15,rand_exe_prng_151_io_out_14,rand_exe_prng_151_io_out_13,
    rand_exe_prng_151_io_out_12,rand_exe_prng_151_io_out_11,rand_exe_prng_151_io_out_10,rand_exe_prng_151_io_out_9,
    rand_exe_prng_151_io_out_8,rand_exe_lo_151}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_152 = {rand_exe_prng_152_io_out_7,rand_exe_prng_152_io_out_6,rand_exe_prng_152_io_out_5,
    rand_exe_prng_152_io_out_4,rand_exe_prng_152_io_out_3,rand_exe_prng_152_io_out_2,rand_exe_prng_152_io_out_1,
    rand_exe_prng_152_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_152 = {rand_exe_prng_152_io_out_15,rand_exe_prng_152_io_out_14,rand_exe_prng_152_io_out_13,
    rand_exe_prng_152_io_out_12,rand_exe_prng_152_io_out_11,rand_exe_prng_152_io_out_10,rand_exe_prng_152_io_out_9,
    rand_exe_prng_152_io_out_8,rand_exe_lo_152}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_153 = {rand_exe_prng_153_io_out_7,rand_exe_prng_153_io_out_6,rand_exe_prng_153_io_out_5,
    rand_exe_prng_153_io_out_4,rand_exe_prng_153_io_out_3,rand_exe_prng_153_io_out_2,rand_exe_prng_153_io_out_1,
    rand_exe_prng_153_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_153 = {rand_exe_prng_153_io_out_15,rand_exe_prng_153_io_out_14,rand_exe_prng_153_io_out_13,
    rand_exe_prng_153_io_out_12,rand_exe_prng_153_io_out_11,rand_exe_prng_153_io_out_10,rand_exe_prng_153_io_out_9,
    rand_exe_prng_153_io_out_8,rand_exe_lo_153}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_154 = {rand_exe_prng_154_io_out_7,rand_exe_prng_154_io_out_6,rand_exe_prng_154_io_out_5,
    rand_exe_prng_154_io_out_4,rand_exe_prng_154_io_out_3,rand_exe_prng_154_io_out_2,rand_exe_prng_154_io_out_1,
    rand_exe_prng_154_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_154 = {rand_exe_prng_154_io_out_15,rand_exe_prng_154_io_out_14,rand_exe_prng_154_io_out_13,
    rand_exe_prng_154_io_out_12,rand_exe_prng_154_io_out_11,rand_exe_prng_154_io_out_10,rand_exe_prng_154_io_out_9,
    rand_exe_prng_154_io_out_8,rand_exe_lo_154}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_155 = {rand_exe_prng_155_io_out_7,rand_exe_prng_155_io_out_6,rand_exe_prng_155_io_out_5,
    rand_exe_prng_155_io_out_4,rand_exe_prng_155_io_out_3,rand_exe_prng_155_io_out_2,rand_exe_prng_155_io_out_1,
    rand_exe_prng_155_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_155 = {rand_exe_prng_155_io_out_15,rand_exe_prng_155_io_out_14,rand_exe_prng_155_io_out_13,
    rand_exe_prng_155_io_out_12,rand_exe_prng_155_io_out_11,rand_exe_prng_155_io_out_10,rand_exe_prng_155_io_out_9,
    rand_exe_prng_155_io_out_8,rand_exe_lo_155}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_156 = {rand_exe_prng_156_io_out_7,rand_exe_prng_156_io_out_6,rand_exe_prng_156_io_out_5,
    rand_exe_prng_156_io_out_4,rand_exe_prng_156_io_out_3,rand_exe_prng_156_io_out_2,rand_exe_prng_156_io_out_1,
    rand_exe_prng_156_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_156 = {rand_exe_prng_156_io_out_15,rand_exe_prng_156_io_out_14,rand_exe_prng_156_io_out_13,
    rand_exe_prng_156_io_out_12,rand_exe_prng_156_io_out_11,rand_exe_prng_156_io_out_10,rand_exe_prng_156_io_out_9,
    rand_exe_prng_156_io_out_8,rand_exe_lo_156}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_157 = {rand_exe_prng_157_io_out_7,rand_exe_prng_157_io_out_6,rand_exe_prng_157_io_out_5,
    rand_exe_prng_157_io_out_4,rand_exe_prng_157_io_out_3,rand_exe_prng_157_io_out_2,rand_exe_prng_157_io_out_1,
    rand_exe_prng_157_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_157 = {rand_exe_prng_157_io_out_15,rand_exe_prng_157_io_out_14,rand_exe_prng_157_io_out_13,
    rand_exe_prng_157_io_out_12,rand_exe_prng_157_io_out_11,rand_exe_prng_157_io_out_10,rand_exe_prng_157_io_out_9,
    rand_exe_prng_157_io_out_8,rand_exe_lo_157}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_158 = {rand_exe_prng_158_io_out_7,rand_exe_prng_158_io_out_6,rand_exe_prng_158_io_out_5,
    rand_exe_prng_158_io_out_4,rand_exe_prng_158_io_out_3,rand_exe_prng_158_io_out_2,rand_exe_prng_158_io_out_1,
    rand_exe_prng_158_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_158 = {rand_exe_prng_158_io_out_15,rand_exe_prng_158_io_out_14,rand_exe_prng_158_io_out_13,
    rand_exe_prng_158_io_out_12,rand_exe_prng_158_io_out_11,rand_exe_prng_158_io_out_10,rand_exe_prng_158_io_out_9,
    rand_exe_prng_158_io_out_8,rand_exe_lo_158}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_159 = {rand_exe_prng_159_io_out_7,rand_exe_prng_159_io_out_6,rand_exe_prng_159_io_out_5,
    rand_exe_prng_159_io_out_4,rand_exe_prng_159_io_out_3,rand_exe_prng_159_io_out_2,rand_exe_prng_159_io_out_1,
    rand_exe_prng_159_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_159 = {rand_exe_prng_159_io_out_15,rand_exe_prng_159_io_out_14,rand_exe_prng_159_io_out_13,
    rand_exe_prng_159_io_out_12,rand_exe_prng_159_io_out_11,rand_exe_prng_159_io_out_10,rand_exe_prng_159_io_out_9,
    rand_exe_prng_159_io_out_8,rand_exe_lo_159}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_160 = {rand_exe_prng_160_io_out_7,rand_exe_prng_160_io_out_6,rand_exe_prng_160_io_out_5,
    rand_exe_prng_160_io_out_4,rand_exe_prng_160_io_out_3,rand_exe_prng_160_io_out_2,rand_exe_prng_160_io_out_1,
    rand_exe_prng_160_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_160 = {rand_exe_prng_160_io_out_15,rand_exe_prng_160_io_out_14,rand_exe_prng_160_io_out_13,
    rand_exe_prng_160_io_out_12,rand_exe_prng_160_io_out_11,rand_exe_prng_160_io_out_10,rand_exe_prng_160_io_out_9,
    rand_exe_prng_160_io_out_8,rand_exe_lo_160}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_161 = {rand_exe_prng_161_io_out_7,rand_exe_prng_161_io_out_6,rand_exe_prng_161_io_out_5,
    rand_exe_prng_161_io_out_4,rand_exe_prng_161_io_out_3,rand_exe_prng_161_io_out_2,rand_exe_prng_161_io_out_1,
    rand_exe_prng_161_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_161 = {rand_exe_prng_161_io_out_15,rand_exe_prng_161_io_out_14,rand_exe_prng_161_io_out_13,
    rand_exe_prng_161_io_out_12,rand_exe_prng_161_io_out_11,rand_exe_prng_161_io_out_10,rand_exe_prng_161_io_out_9,
    rand_exe_prng_161_io_out_8,rand_exe_lo_161}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_162 = {rand_exe_prng_162_io_out_7,rand_exe_prng_162_io_out_6,rand_exe_prng_162_io_out_5,
    rand_exe_prng_162_io_out_4,rand_exe_prng_162_io_out_3,rand_exe_prng_162_io_out_2,rand_exe_prng_162_io_out_1,
    rand_exe_prng_162_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_162 = {rand_exe_prng_162_io_out_15,rand_exe_prng_162_io_out_14,rand_exe_prng_162_io_out_13,
    rand_exe_prng_162_io_out_12,rand_exe_prng_162_io_out_11,rand_exe_prng_162_io_out_10,rand_exe_prng_162_io_out_9,
    rand_exe_prng_162_io_out_8,rand_exe_lo_162}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_163 = {rand_exe_prng_163_io_out_7,rand_exe_prng_163_io_out_6,rand_exe_prng_163_io_out_5,
    rand_exe_prng_163_io_out_4,rand_exe_prng_163_io_out_3,rand_exe_prng_163_io_out_2,rand_exe_prng_163_io_out_1,
    rand_exe_prng_163_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_163 = {rand_exe_prng_163_io_out_15,rand_exe_prng_163_io_out_14,rand_exe_prng_163_io_out_13,
    rand_exe_prng_163_io_out_12,rand_exe_prng_163_io_out_11,rand_exe_prng_163_io_out_10,rand_exe_prng_163_io_out_9,
    rand_exe_prng_163_io_out_8,rand_exe_lo_163}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_164 = {rand_exe_prng_164_io_out_7,rand_exe_prng_164_io_out_6,rand_exe_prng_164_io_out_5,
    rand_exe_prng_164_io_out_4,rand_exe_prng_164_io_out_3,rand_exe_prng_164_io_out_2,rand_exe_prng_164_io_out_1,
    rand_exe_prng_164_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_164 = {rand_exe_prng_164_io_out_15,rand_exe_prng_164_io_out_14,rand_exe_prng_164_io_out_13,
    rand_exe_prng_164_io_out_12,rand_exe_prng_164_io_out_11,rand_exe_prng_164_io_out_10,rand_exe_prng_164_io_out_9,
    rand_exe_prng_164_io_out_8,rand_exe_lo_164}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_165 = {rand_exe_prng_165_io_out_7,rand_exe_prng_165_io_out_6,rand_exe_prng_165_io_out_5,
    rand_exe_prng_165_io_out_4,rand_exe_prng_165_io_out_3,rand_exe_prng_165_io_out_2,rand_exe_prng_165_io_out_1,
    rand_exe_prng_165_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_165 = {rand_exe_prng_165_io_out_15,rand_exe_prng_165_io_out_14,rand_exe_prng_165_io_out_13,
    rand_exe_prng_165_io_out_12,rand_exe_prng_165_io_out_11,rand_exe_prng_165_io_out_10,rand_exe_prng_165_io_out_9,
    rand_exe_prng_165_io_out_8,rand_exe_lo_165}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_166 = {rand_exe_prng_166_io_out_7,rand_exe_prng_166_io_out_6,rand_exe_prng_166_io_out_5,
    rand_exe_prng_166_io_out_4,rand_exe_prng_166_io_out_3,rand_exe_prng_166_io_out_2,rand_exe_prng_166_io_out_1,
    rand_exe_prng_166_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_166 = {rand_exe_prng_166_io_out_15,rand_exe_prng_166_io_out_14,rand_exe_prng_166_io_out_13,
    rand_exe_prng_166_io_out_12,rand_exe_prng_166_io_out_11,rand_exe_prng_166_io_out_10,rand_exe_prng_166_io_out_9,
    rand_exe_prng_166_io_out_8,rand_exe_lo_166}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_167 = {rand_exe_prng_167_io_out_7,rand_exe_prng_167_io_out_6,rand_exe_prng_167_io_out_5,
    rand_exe_prng_167_io_out_4,rand_exe_prng_167_io_out_3,rand_exe_prng_167_io_out_2,rand_exe_prng_167_io_out_1,
    rand_exe_prng_167_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_167 = {rand_exe_prng_167_io_out_15,rand_exe_prng_167_io_out_14,rand_exe_prng_167_io_out_13,
    rand_exe_prng_167_io_out_12,rand_exe_prng_167_io_out_11,rand_exe_prng_167_io_out_10,rand_exe_prng_167_io_out_9,
    rand_exe_prng_167_io_out_8,rand_exe_lo_167}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_168 = {rand_exe_prng_168_io_out_7,rand_exe_prng_168_io_out_6,rand_exe_prng_168_io_out_5,
    rand_exe_prng_168_io_out_4,rand_exe_prng_168_io_out_3,rand_exe_prng_168_io_out_2,rand_exe_prng_168_io_out_1,
    rand_exe_prng_168_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_168 = {rand_exe_prng_168_io_out_15,rand_exe_prng_168_io_out_14,rand_exe_prng_168_io_out_13,
    rand_exe_prng_168_io_out_12,rand_exe_prng_168_io_out_11,rand_exe_prng_168_io_out_10,rand_exe_prng_168_io_out_9,
    rand_exe_prng_168_io_out_8,rand_exe_lo_168}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_169 = {rand_exe_prng_169_io_out_7,rand_exe_prng_169_io_out_6,rand_exe_prng_169_io_out_5,
    rand_exe_prng_169_io_out_4,rand_exe_prng_169_io_out_3,rand_exe_prng_169_io_out_2,rand_exe_prng_169_io_out_1,
    rand_exe_prng_169_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_169 = {rand_exe_prng_169_io_out_15,rand_exe_prng_169_io_out_14,rand_exe_prng_169_io_out_13,
    rand_exe_prng_169_io_out_12,rand_exe_prng_169_io_out_11,rand_exe_prng_169_io_out_10,rand_exe_prng_169_io_out_9,
    rand_exe_prng_169_io_out_8,rand_exe_lo_169}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_170 = {rand_exe_prng_170_io_out_7,rand_exe_prng_170_io_out_6,rand_exe_prng_170_io_out_5,
    rand_exe_prng_170_io_out_4,rand_exe_prng_170_io_out_3,rand_exe_prng_170_io_out_2,rand_exe_prng_170_io_out_1,
    rand_exe_prng_170_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_170 = {rand_exe_prng_170_io_out_15,rand_exe_prng_170_io_out_14,rand_exe_prng_170_io_out_13,
    rand_exe_prng_170_io_out_12,rand_exe_prng_170_io_out_11,rand_exe_prng_170_io_out_10,rand_exe_prng_170_io_out_9,
    rand_exe_prng_170_io_out_8,rand_exe_lo_170}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_171 = {rand_exe_prng_171_io_out_7,rand_exe_prng_171_io_out_6,rand_exe_prng_171_io_out_5,
    rand_exe_prng_171_io_out_4,rand_exe_prng_171_io_out_3,rand_exe_prng_171_io_out_2,rand_exe_prng_171_io_out_1,
    rand_exe_prng_171_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_171 = {rand_exe_prng_171_io_out_15,rand_exe_prng_171_io_out_14,rand_exe_prng_171_io_out_13,
    rand_exe_prng_171_io_out_12,rand_exe_prng_171_io_out_11,rand_exe_prng_171_io_out_10,rand_exe_prng_171_io_out_9,
    rand_exe_prng_171_io_out_8,rand_exe_lo_171}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_172 = {rand_exe_prng_172_io_out_7,rand_exe_prng_172_io_out_6,rand_exe_prng_172_io_out_5,
    rand_exe_prng_172_io_out_4,rand_exe_prng_172_io_out_3,rand_exe_prng_172_io_out_2,rand_exe_prng_172_io_out_1,
    rand_exe_prng_172_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_172 = {rand_exe_prng_172_io_out_15,rand_exe_prng_172_io_out_14,rand_exe_prng_172_io_out_13,
    rand_exe_prng_172_io_out_12,rand_exe_prng_172_io_out_11,rand_exe_prng_172_io_out_10,rand_exe_prng_172_io_out_9,
    rand_exe_prng_172_io_out_8,rand_exe_lo_172}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_173 = {rand_exe_prng_173_io_out_7,rand_exe_prng_173_io_out_6,rand_exe_prng_173_io_out_5,
    rand_exe_prng_173_io_out_4,rand_exe_prng_173_io_out_3,rand_exe_prng_173_io_out_2,rand_exe_prng_173_io_out_1,
    rand_exe_prng_173_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_173 = {rand_exe_prng_173_io_out_15,rand_exe_prng_173_io_out_14,rand_exe_prng_173_io_out_13,
    rand_exe_prng_173_io_out_12,rand_exe_prng_173_io_out_11,rand_exe_prng_173_io_out_10,rand_exe_prng_173_io_out_9,
    rand_exe_prng_173_io_out_8,rand_exe_lo_173}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_174 = {rand_exe_prng_174_io_out_7,rand_exe_prng_174_io_out_6,rand_exe_prng_174_io_out_5,
    rand_exe_prng_174_io_out_4,rand_exe_prng_174_io_out_3,rand_exe_prng_174_io_out_2,rand_exe_prng_174_io_out_1,
    rand_exe_prng_174_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_174 = {rand_exe_prng_174_io_out_15,rand_exe_prng_174_io_out_14,rand_exe_prng_174_io_out_13,
    rand_exe_prng_174_io_out_12,rand_exe_prng_174_io_out_11,rand_exe_prng_174_io_out_10,rand_exe_prng_174_io_out_9,
    rand_exe_prng_174_io_out_8,rand_exe_lo_174}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_175 = {rand_exe_prng_175_io_out_7,rand_exe_prng_175_io_out_6,rand_exe_prng_175_io_out_5,
    rand_exe_prng_175_io_out_4,rand_exe_prng_175_io_out_3,rand_exe_prng_175_io_out_2,rand_exe_prng_175_io_out_1,
    rand_exe_prng_175_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_175 = {rand_exe_prng_175_io_out_15,rand_exe_prng_175_io_out_14,rand_exe_prng_175_io_out_13,
    rand_exe_prng_175_io_out_12,rand_exe_prng_175_io_out_11,rand_exe_prng_175_io_out_10,rand_exe_prng_175_io_out_9,
    rand_exe_prng_175_io_out_8,rand_exe_lo_175}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_176 = {rand_exe_prng_176_io_out_7,rand_exe_prng_176_io_out_6,rand_exe_prng_176_io_out_5,
    rand_exe_prng_176_io_out_4,rand_exe_prng_176_io_out_3,rand_exe_prng_176_io_out_2,rand_exe_prng_176_io_out_1,
    rand_exe_prng_176_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_176 = {rand_exe_prng_176_io_out_15,rand_exe_prng_176_io_out_14,rand_exe_prng_176_io_out_13,
    rand_exe_prng_176_io_out_12,rand_exe_prng_176_io_out_11,rand_exe_prng_176_io_out_10,rand_exe_prng_176_io_out_9,
    rand_exe_prng_176_io_out_8,rand_exe_lo_176}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_177 = {rand_exe_prng_177_io_out_7,rand_exe_prng_177_io_out_6,rand_exe_prng_177_io_out_5,
    rand_exe_prng_177_io_out_4,rand_exe_prng_177_io_out_3,rand_exe_prng_177_io_out_2,rand_exe_prng_177_io_out_1,
    rand_exe_prng_177_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_177 = {rand_exe_prng_177_io_out_15,rand_exe_prng_177_io_out_14,rand_exe_prng_177_io_out_13,
    rand_exe_prng_177_io_out_12,rand_exe_prng_177_io_out_11,rand_exe_prng_177_io_out_10,rand_exe_prng_177_io_out_9,
    rand_exe_prng_177_io_out_8,rand_exe_lo_177}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_178 = {rand_exe_prng_178_io_out_7,rand_exe_prng_178_io_out_6,rand_exe_prng_178_io_out_5,
    rand_exe_prng_178_io_out_4,rand_exe_prng_178_io_out_3,rand_exe_prng_178_io_out_2,rand_exe_prng_178_io_out_1,
    rand_exe_prng_178_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_178 = {rand_exe_prng_178_io_out_15,rand_exe_prng_178_io_out_14,rand_exe_prng_178_io_out_13,
    rand_exe_prng_178_io_out_12,rand_exe_prng_178_io_out_11,rand_exe_prng_178_io_out_10,rand_exe_prng_178_io_out_9,
    rand_exe_prng_178_io_out_8,rand_exe_lo_178}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_179 = {rand_exe_prng_179_io_out_7,rand_exe_prng_179_io_out_6,rand_exe_prng_179_io_out_5,
    rand_exe_prng_179_io_out_4,rand_exe_prng_179_io_out_3,rand_exe_prng_179_io_out_2,rand_exe_prng_179_io_out_1,
    rand_exe_prng_179_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_179 = {rand_exe_prng_179_io_out_15,rand_exe_prng_179_io_out_14,rand_exe_prng_179_io_out_13,
    rand_exe_prng_179_io_out_12,rand_exe_prng_179_io_out_11,rand_exe_prng_179_io_out_10,rand_exe_prng_179_io_out_9,
    rand_exe_prng_179_io_out_8,rand_exe_lo_179}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_180 = {rand_exe_prng_180_io_out_7,rand_exe_prng_180_io_out_6,rand_exe_prng_180_io_out_5,
    rand_exe_prng_180_io_out_4,rand_exe_prng_180_io_out_3,rand_exe_prng_180_io_out_2,rand_exe_prng_180_io_out_1,
    rand_exe_prng_180_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_180 = {rand_exe_prng_180_io_out_15,rand_exe_prng_180_io_out_14,rand_exe_prng_180_io_out_13,
    rand_exe_prng_180_io_out_12,rand_exe_prng_180_io_out_11,rand_exe_prng_180_io_out_10,rand_exe_prng_180_io_out_9,
    rand_exe_prng_180_io_out_8,rand_exe_lo_180}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_181 = {rand_exe_prng_181_io_out_7,rand_exe_prng_181_io_out_6,rand_exe_prng_181_io_out_5,
    rand_exe_prng_181_io_out_4,rand_exe_prng_181_io_out_3,rand_exe_prng_181_io_out_2,rand_exe_prng_181_io_out_1,
    rand_exe_prng_181_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_181 = {rand_exe_prng_181_io_out_15,rand_exe_prng_181_io_out_14,rand_exe_prng_181_io_out_13,
    rand_exe_prng_181_io_out_12,rand_exe_prng_181_io_out_11,rand_exe_prng_181_io_out_10,rand_exe_prng_181_io_out_9,
    rand_exe_prng_181_io_out_8,rand_exe_lo_181}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_182 = {rand_exe_prng_182_io_out_7,rand_exe_prng_182_io_out_6,rand_exe_prng_182_io_out_5,
    rand_exe_prng_182_io_out_4,rand_exe_prng_182_io_out_3,rand_exe_prng_182_io_out_2,rand_exe_prng_182_io_out_1,
    rand_exe_prng_182_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_182 = {rand_exe_prng_182_io_out_15,rand_exe_prng_182_io_out_14,rand_exe_prng_182_io_out_13,
    rand_exe_prng_182_io_out_12,rand_exe_prng_182_io_out_11,rand_exe_prng_182_io_out_10,rand_exe_prng_182_io_out_9,
    rand_exe_prng_182_io_out_8,rand_exe_lo_182}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_183 = {rand_exe_prng_183_io_out_7,rand_exe_prng_183_io_out_6,rand_exe_prng_183_io_out_5,
    rand_exe_prng_183_io_out_4,rand_exe_prng_183_io_out_3,rand_exe_prng_183_io_out_2,rand_exe_prng_183_io_out_1,
    rand_exe_prng_183_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_183 = {rand_exe_prng_183_io_out_15,rand_exe_prng_183_io_out_14,rand_exe_prng_183_io_out_13,
    rand_exe_prng_183_io_out_12,rand_exe_prng_183_io_out_11,rand_exe_prng_183_io_out_10,rand_exe_prng_183_io_out_9,
    rand_exe_prng_183_io_out_8,rand_exe_lo_183}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_184 = {rand_exe_prng_184_io_out_7,rand_exe_prng_184_io_out_6,rand_exe_prng_184_io_out_5,
    rand_exe_prng_184_io_out_4,rand_exe_prng_184_io_out_3,rand_exe_prng_184_io_out_2,rand_exe_prng_184_io_out_1,
    rand_exe_prng_184_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_184 = {rand_exe_prng_184_io_out_15,rand_exe_prng_184_io_out_14,rand_exe_prng_184_io_out_13,
    rand_exe_prng_184_io_out_12,rand_exe_prng_184_io_out_11,rand_exe_prng_184_io_out_10,rand_exe_prng_184_io_out_9,
    rand_exe_prng_184_io_out_8,rand_exe_lo_184}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_185 = {rand_exe_prng_185_io_out_7,rand_exe_prng_185_io_out_6,rand_exe_prng_185_io_out_5,
    rand_exe_prng_185_io_out_4,rand_exe_prng_185_io_out_3,rand_exe_prng_185_io_out_2,rand_exe_prng_185_io_out_1,
    rand_exe_prng_185_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_185 = {rand_exe_prng_185_io_out_15,rand_exe_prng_185_io_out_14,rand_exe_prng_185_io_out_13,
    rand_exe_prng_185_io_out_12,rand_exe_prng_185_io_out_11,rand_exe_prng_185_io_out_10,rand_exe_prng_185_io_out_9,
    rand_exe_prng_185_io_out_8,rand_exe_lo_185}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_186 = {rand_exe_prng_186_io_out_7,rand_exe_prng_186_io_out_6,rand_exe_prng_186_io_out_5,
    rand_exe_prng_186_io_out_4,rand_exe_prng_186_io_out_3,rand_exe_prng_186_io_out_2,rand_exe_prng_186_io_out_1,
    rand_exe_prng_186_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_186 = {rand_exe_prng_186_io_out_15,rand_exe_prng_186_io_out_14,rand_exe_prng_186_io_out_13,
    rand_exe_prng_186_io_out_12,rand_exe_prng_186_io_out_11,rand_exe_prng_186_io_out_10,rand_exe_prng_186_io_out_9,
    rand_exe_prng_186_io_out_8,rand_exe_lo_186}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_187 = {rand_exe_prng_187_io_out_7,rand_exe_prng_187_io_out_6,rand_exe_prng_187_io_out_5,
    rand_exe_prng_187_io_out_4,rand_exe_prng_187_io_out_3,rand_exe_prng_187_io_out_2,rand_exe_prng_187_io_out_1,
    rand_exe_prng_187_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_187 = {rand_exe_prng_187_io_out_15,rand_exe_prng_187_io_out_14,rand_exe_prng_187_io_out_13,
    rand_exe_prng_187_io_out_12,rand_exe_prng_187_io_out_11,rand_exe_prng_187_io_out_10,rand_exe_prng_187_io_out_9,
    rand_exe_prng_187_io_out_8,rand_exe_lo_187}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_188 = {rand_exe_prng_188_io_out_7,rand_exe_prng_188_io_out_6,rand_exe_prng_188_io_out_5,
    rand_exe_prng_188_io_out_4,rand_exe_prng_188_io_out_3,rand_exe_prng_188_io_out_2,rand_exe_prng_188_io_out_1,
    rand_exe_prng_188_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_188 = {rand_exe_prng_188_io_out_15,rand_exe_prng_188_io_out_14,rand_exe_prng_188_io_out_13,
    rand_exe_prng_188_io_out_12,rand_exe_prng_188_io_out_11,rand_exe_prng_188_io_out_10,rand_exe_prng_188_io_out_9,
    rand_exe_prng_188_io_out_8,rand_exe_lo_188}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_189 = {rand_exe_prng_189_io_out_7,rand_exe_prng_189_io_out_6,rand_exe_prng_189_io_out_5,
    rand_exe_prng_189_io_out_4,rand_exe_prng_189_io_out_3,rand_exe_prng_189_io_out_2,rand_exe_prng_189_io_out_1,
    rand_exe_prng_189_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_189 = {rand_exe_prng_189_io_out_15,rand_exe_prng_189_io_out_14,rand_exe_prng_189_io_out_13,
    rand_exe_prng_189_io_out_12,rand_exe_prng_189_io_out_11,rand_exe_prng_189_io_out_10,rand_exe_prng_189_io_out_9,
    rand_exe_prng_189_io_out_8,rand_exe_lo_189}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_190 = {rand_exe_prng_190_io_out_7,rand_exe_prng_190_io_out_6,rand_exe_prng_190_io_out_5,
    rand_exe_prng_190_io_out_4,rand_exe_prng_190_io_out_3,rand_exe_prng_190_io_out_2,rand_exe_prng_190_io_out_1,
    rand_exe_prng_190_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_190 = {rand_exe_prng_190_io_out_15,rand_exe_prng_190_io_out_14,rand_exe_prng_190_io_out_13,
    rand_exe_prng_190_io_out_12,rand_exe_prng_190_io_out_11,rand_exe_prng_190_io_out_10,rand_exe_prng_190_io_out_9,
    rand_exe_prng_190_io_out_8,rand_exe_lo_190}; // @[PRNG.scala 86:17]
  wire [7:0] rand_exe_lo_191 = {rand_exe_prng_191_io_out_7,rand_exe_prng_191_io_out_6,rand_exe_prng_191_io_out_5,
    rand_exe_prng_191_io_out_4,rand_exe_prng_191_io_out_3,rand_exe_prng_191_io_out_2,rand_exe_prng_191_io_out_1,
    rand_exe_prng_191_io_out_0}; // @[PRNG.scala 86:17]
  wire [15:0] rand_191 = {rand_exe_prng_191_io_out_15,rand_exe_prng_191_io_out_14,rand_exe_prng_191_io_out_13,
    rand_exe_prng_191_io_out_12,rand_exe_prng_191_io_out_11,rand_exe_prng_191_io_out_10,rand_exe_prng_191_io_out_9,
    rand_exe_prng_191_io_out_8,rand_exe_lo_191}; // @[PRNG.scala 86:17]
  MaxPeriodFibonacciLFSR rand_exe_prng ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_clock),
    .reset(rand_exe_prng_reset),
    .io_out_0(rand_exe_prng_io_out_0),
    .io_out_1(rand_exe_prng_io_out_1),
    .io_out_2(rand_exe_prng_io_out_2),
    .io_out_3(rand_exe_prng_io_out_3),
    .io_out_4(rand_exe_prng_io_out_4),
    .io_out_5(rand_exe_prng_io_out_5),
    .io_out_6(rand_exe_prng_io_out_6),
    .io_out_7(rand_exe_prng_io_out_7),
    .io_out_8(rand_exe_prng_io_out_8),
    .io_out_9(rand_exe_prng_io_out_9),
    .io_out_10(rand_exe_prng_io_out_10),
    .io_out_11(rand_exe_prng_io_out_11),
    .io_out_12(rand_exe_prng_io_out_12),
    .io_out_13(rand_exe_prng_io_out_13),
    .io_out_14(rand_exe_prng_io_out_14),
    .io_out_15(rand_exe_prng_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_1 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_1_clock),
    .reset(rand_exe_prng_1_reset),
    .io_out_0(rand_exe_prng_1_io_out_0),
    .io_out_1(rand_exe_prng_1_io_out_1),
    .io_out_2(rand_exe_prng_1_io_out_2),
    .io_out_3(rand_exe_prng_1_io_out_3),
    .io_out_4(rand_exe_prng_1_io_out_4),
    .io_out_5(rand_exe_prng_1_io_out_5),
    .io_out_6(rand_exe_prng_1_io_out_6),
    .io_out_7(rand_exe_prng_1_io_out_7),
    .io_out_8(rand_exe_prng_1_io_out_8),
    .io_out_9(rand_exe_prng_1_io_out_9),
    .io_out_10(rand_exe_prng_1_io_out_10),
    .io_out_11(rand_exe_prng_1_io_out_11),
    .io_out_12(rand_exe_prng_1_io_out_12),
    .io_out_13(rand_exe_prng_1_io_out_13),
    .io_out_14(rand_exe_prng_1_io_out_14),
    .io_out_15(rand_exe_prng_1_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_2 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_2_clock),
    .reset(rand_exe_prng_2_reset),
    .io_out_0(rand_exe_prng_2_io_out_0),
    .io_out_1(rand_exe_prng_2_io_out_1),
    .io_out_2(rand_exe_prng_2_io_out_2),
    .io_out_3(rand_exe_prng_2_io_out_3),
    .io_out_4(rand_exe_prng_2_io_out_4),
    .io_out_5(rand_exe_prng_2_io_out_5),
    .io_out_6(rand_exe_prng_2_io_out_6),
    .io_out_7(rand_exe_prng_2_io_out_7),
    .io_out_8(rand_exe_prng_2_io_out_8),
    .io_out_9(rand_exe_prng_2_io_out_9),
    .io_out_10(rand_exe_prng_2_io_out_10),
    .io_out_11(rand_exe_prng_2_io_out_11),
    .io_out_12(rand_exe_prng_2_io_out_12),
    .io_out_13(rand_exe_prng_2_io_out_13),
    .io_out_14(rand_exe_prng_2_io_out_14),
    .io_out_15(rand_exe_prng_2_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_3 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_3_clock),
    .reset(rand_exe_prng_3_reset),
    .io_out_0(rand_exe_prng_3_io_out_0),
    .io_out_1(rand_exe_prng_3_io_out_1),
    .io_out_2(rand_exe_prng_3_io_out_2),
    .io_out_3(rand_exe_prng_3_io_out_3),
    .io_out_4(rand_exe_prng_3_io_out_4),
    .io_out_5(rand_exe_prng_3_io_out_5),
    .io_out_6(rand_exe_prng_3_io_out_6),
    .io_out_7(rand_exe_prng_3_io_out_7),
    .io_out_8(rand_exe_prng_3_io_out_8),
    .io_out_9(rand_exe_prng_3_io_out_9),
    .io_out_10(rand_exe_prng_3_io_out_10),
    .io_out_11(rand_exe_prng_3_io_out_11),
    .io_out_12(rand_exe_prng_3_io_out_12),
    .io_out_13(rand_exe_prng_3_io_out_13),
    .io_out_14(rand_exe_prng_3_io_out_14),
    .io_out_15(rand_exe_prng_3_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_4 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_4_clock),
    .reset(rand_exe_prng_4_reset),
    .io_out_0(rand_exe_prng_4_io_out_0),
    .io_out_1(rand_exe_prng_4_io_out_1),
    .io_out_2(rand_exe_prng_4_io_out_2),
    .io_out_3(rand_exe_prng_4_io_out_3),
    .io_out_4(rand_exe_prng_4_io_out_4),
    .io_out_5(rand_exe_prng_4_io_out_5),
    .io_out_6(rand_exe_prng_4_io_out_6),
    .io_out_7(rand_exe_prng_4_io_out_7),
    .io_out_8(rand_exe_prng_4_io_out_8),
    .io_out_9(rand_exe_prng_4_io_out_9),
    .io_out_10(rand_exe_prng_4_io_out_10),
    .io_out_11(rand_exe_prng_4_io_out_11),
    .io_out_12(rand_exe_prng_4_io_out_12),
    .io_out_13(rand_exe_prng_4_io_out_13),
    .io_out_14(rand_exe_prng_4_io_out_14),
    .io_out_15(rand_exe_prng_4_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_5 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_5_clock),
    .reset(rand_exe_prng_5_reset),
    .io_out_0(rand_exe_prng_5_io_out_0),
    .io_out_1(rand_exe_prng_5_io_out_1),
    .io_out_2(rand_exe_prng_5_io_out_2),
    .io_out_3(rand_exe_prng_5_io_out_3),
    .io_out_4(rand_exe_prng_5_io_out_4),
    .io_out_5(rand_exe_prng_5_io_out_5),
    .io_out_6(rand_exe_prng_5_io_out_6),
    .io_out_7(rand_exe_prng_5_io_out_7),
    .io_out_8(rand_exe_prng_5_io_out_8),
    .io_out_9(rand_exe_prng_5_io_out_9),
    .io_out_10(rand_exe_prng_5_io_out_10),
    .io_out_11(rand_exe_prng_5_io_out_11),
    .io_out_12(rand_exe_prng_5_io_out_12),
    .io_out_13(rand_exe_prng_5_io_out_13),
    .io_out_14(rand_exe_prng_5_io_out_14),
    .io_out_15(rand_exe_prng_5_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_6 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_6_clock),
    .reset(rand_exe_prng_6_reset),
    .io_out_0(rand_exe_prng_6_io_out_0),
    .io_out_1(rand_exe_prng_6_io_out_1),
    .io_out_2(rand_exe_prng_6_io_out_2),
    .io_out_3(rand_exe_prng_6_io_out_3),
    .io_out_4(rand_exe_prng_6_io_out_4),
    .io_out_5(rand_exe_prng_6_io_out_5),
    .io_out_6(rand_exe_prng_6_io_out_6),
    .io_out_7(rand_exe_prng_6_io_out_7),
    .io_out_8(rand_exe_prng_6_io_out_8),
    .io_out_9(rand_exe_prng_6_io_out_9),
    .io_out_10(rand_exe_prng_6_io_out_10),
    .io_out_11(rand_exe_prng_6_io_out_11),
    .io_out_12(rand_exe_prng_6_io_out_12),
    .io_out_13(rand_exe_prng_6_io_out_13),
    .io_out_14(rand_exe_prng_6_io_out_14),
    .io_out_15(rand_exe_prng_6_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_7 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_7_clock),
    .reset(rand_exe_prng_7_reset),
    .io_out_0(rand_exe_prng_7_io_out_0),
    .io_out_1(rand_exe_prng_7_io_out_1),
    .io_out_2(rand_exe_prng_7_io_out_2),
    .io_out_3(rand_exe_prng_7_io_out_3),
    .io_out_4(rand_exe_prng_7_io_out_4),
    .io_out_5(rand_exe_prng_7_io_out_5),
    .io_out_6(rand_exe_prng_7_io_out_6),
    .io_out_7(rand_exe_prng_7_io_out_7),
    .io_out_8(rand_exe_prng_7_io_out_8),
    .io_out_9(rand_exe_prng_7_io_out_9),
    .io_out_10(rand_exe_prng_7_io_out_10),
    .io_out_11(rand_exe_prng_7_io_out_11),
    .io_out_12(rand_exe_prng_7_io_out_12),
    .io_out_13(rand_exe_prng_7_io_out_13),
    .io_out_14(rand_exe_prng_7_io_out_14),
    .io_out_15(rand_exe_prng_7_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_8 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_8_clock),
    .reset(rand_exe_prng_8_reset),
    .io_out_0(rand_exe_prng_8_io_out_0),
    .io_out_1(rand_exe_prng_8_io_out_1),
    .io_out_2(rand_exe_prng_8_io_out_2),
    .io_out_3(rand_exe_prng_8_io_out_3),
    .io_out_4(rand_exe_prng_8_io_out_4),
    .io_out_5(rand_exe_prng_8_io_out_5),
    .io_out_6(rand_exe_prng_8_io_out_6),
    .io_out_7(rand_exe_prng_8_io_out_7),
    .io_out_8(rand_exe_prng_8_io_out_8),
    .io_out_9(rand_exe_prng_8_io_out_9),
    .io_out_10(rand_exe_prng_8_io_out_10),
    .io_out_11(rand_exe_prng_8_io_out_11),
    .io_out_12(rand_exe_prng_8_io_out_12),
    .io_out_13(rand_exe_prng_8_io_out_13),
    .io_out_14(rand_exe_prng_8_io_out_14),
    .io_out_15(rand_exe_prng_8_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_9 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_9_clock),
    .reset(rand_exe_prng_9_reset),
    .io_out_0(rand_exe_prng_9_io_out_0),
    .io_out_1(rand_exe_prng_9_io_out_1),
    .io_out_2(rand_exe_prng_9_io_out_2),
    .io_out_3(rand_exe_prng_9_io_out_3),
    .io_out_4(rand_exe_prng_9_io_out_4),
    .io_out_5(rand_exe_prng_9_io_out_5),
    .io_out_6(rand_exe_prng_9_io_out_6),
    .io_out_7(rand_exe_prng_9_io_out_7),
    .io_out_8(rand_exe_prng_9_io_out_8),
    .io_out_9(rand_exe_prng_9_io_out_9),
    .io_out_10(rand_exe_prng_9_io_out_10),
    .io_out_11(rand_exe_prng_9_io_out_11),
    .io_out_12(rand_exe_prng_9_io_out_12),
    .io_out_13(rand_exe_prng_9_io_out_13),
    .io_out_14(rand_exe_prng_9_io_out_14),
    .io_out_15(rand_exe_prng_9_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_10 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_10_clock),
    .reset(rand_exe_prng_10_reset),
    .io_out_0(rand_exe_prng_10_io_out_0),
    .io_out_1(rand_exe_prng_10_io_out_1),
    .io_out_2(rand_exe_prng_10_io_out_2),
    .io_out_3(rand_exe_prng_10_io_out_3),
    .io_out_4(rand_exe_prng_10_io_out_4),
    .io_out_5(rand_exe_prng_10_io_out_5),
    .io_out_6(rand_exe_prng_10_io_out_6),
    .io_out_7(rand_exe_prng_10_io_out_7),
    .io_out_8(rand_exe_prng_10_io_out_8),
    .io_out_9(rand_exe_prng_10_io_out_9),
    .io_out_10(rand_exe_prng_10_io_out_10),
    .io_out_11(rand_exe_prng_10_io_out_11),
    .io_out_12(rand_exe_prng_10_io_out_12),
    .io_out_13(rand_exe_prng_10_io_out_13),
    .io_out_14(rand_exe_prng_10_io_out_14),
    .io_out_15(rand_exe_prng_10_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_11 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_11_clock),
    .reset(rand_exe_prng_11_reset),
    .io_out_0(rand_exe_prng_11_io_out_0),
    .io_out_1(rand_exe_prng_11_io_out_1),
    .io_out_2(rand_exe_prng_11_io_out_2),
    .io_out_3(rand_exe_prng_11_io_out_3),
    .io_out_4(rand_exe_prng_11_io_out_4),
    .io_out_5(rand_exe_prng_11_io_out_5),
    .io_out_6(rand_exe_prng_11_io_out_6),
    .io_out_7(rand_exe_prng_11_io_out_7),
    .io_out_8(rand_exe_prng_11_io_out_8),
    .io_out_9(rand_exe_prng_11_io_out_9),
    .io_out_10(rand_exe_prng_11_io_out_10),
    .io_out_11(rand_exe_prng_11_io_out_11),
    .io_out_12(rand_exe_prng_11_io_out_12),
    .io_out_13(rand_exe_prng_11_io_out_13),
    .io_out_14(rand_exe_prng_11_io_out_14),
    .io_out_15(rand_exe_prng_11_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_12 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_12_clock),
    .reset(rand_exe_prng_12_reset),
    .io_out_0(rand_exe_prng_12_io_out_0),
    .io_out_1(rand_exe_prng_12_io_out_1),
    .io_out_2(rand_exe_prng_12_io_out_2),
    .io_out_3(rand_exe_prng_12_io_out_3),
    .io_out_4(rand_exe_prng_12_io_out_4),
    .io_out_5(rand_exe_prng_12_io_out_5),
    .io_out_6(rand_exe_prng_12_io_out_6),
    .io_out_7(rand_exe_prng_12_io_out_7),
    .io_out_8(rand_exe_prng_12_io_out_8),
    .io_out_9(rand_exe_prng_12_io_out_9),
    .io_out_10(rand_exe_prng_12_io_out_10),
    .io_out_11(rand_exe_prng_12_io_out_11),
    .io_out_12(rand_exe_prng_12_io_out_12),
    .io_out_13(rand_exe_prng_12_io_out_13),
    .io_out_14(rand_exe_prng_12_io_out_14),
    .io_out_15(rand_exe_prng_12_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_13 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_13_clock),
    .reset(rand_exe_prng_13_reset),
    .io_out_0(rand_exe_prng_13_io_out_0),
    .io_out_1(rand_exe_prng_13_io_out_1),
    .io_out_2(rand_exe_prng_13_io_out_2),
    .io_out_3(rand_exe_prng_13_io_out_3),
    .io_out_4(rand_exe_prng_13_io_out_4),
    .io_out_5(rand_exe_prng_13_io_out_5),
    .io_out_6(rand_exe_prng_13_io_out_6),
    .io_out_7(rand_exe_prng_13_io_out_7),
    .io_out_8(rand_exe_prng_13_io_out_8),
    .io_out_9(rand_exe_prng_13_io_out_9),
    .io_out_10(rand_exe_prng_13_io_out_10),
    .io_out_11(rand_exe_prng_13_io_out_11),
    .io_out_12(rand_exe_prng_13_io_out_12),
    .io_out_13(rand_exe_prng_13_io_out_13),
    .io_out_14(rand_exe_prng_13_io_out_14),
    .io_out_15(rand_exe_prng_13_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_14 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_14_clock),
    .reset(rand_exe_prng_14_reset),
    .io_out_0(rand_exe_prng_14_io_out_0),
    .io_out_1(rand_exe_prng_14_io_out_1),
    .io_out_2(rand_exe_prng_14_io_out_2),
    .io_out_3(rand_exe_prng_14_io_out_3),
    .io_out_4(rand_exe_prng_14_io_out_4),
    .io_out_5(rand_exe_prng_14_io_out_5),
    .io_out_6(rand_exe_prng_14_io_out_6),
    .io_out_7(rand_exe_prng_14_io_out_7),
    .io_out_8(rand_exe_prng_14_io_out_8),
    .io_out_9(rand_exe_prng_14_io_out_9),
    .io_out_10(rand_exe_prng_14_io_out_10),
    .io_out_11(rand_exe_prng_14_io_out_11),
    .io_out_12(rand_exe_prng_14_io_out_12),
    .io_out_13(rand_exe_prng_14_io_out_13),
    .io_out_14(rand_exe_prng_14_io_out_14),
    .io_out_15(rand_exe_prng_14_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_15 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_15_clock),
    .reset(rand_exe_prng_15_reset),
    .io_out_0(rand_exe_prng_15_io_out_0),
    .io_out_1(rand_exe_prng_15_io_out_1),
    .io_out_2(rand_exe_prng_15_io_out_2),
    .io_out_3(rand_exe_prng_15_io_out_3),
    .io_out_4(rand_exe_prng_15_io_out_4),
    .io_out_5(rand_exe_prng_15_io_out_5),
    .io_out_6(rand_exe_prng_15_io_out_6),
    .io_out_7(rand_exe_prng_15_io_out_7),
    .io_out_8(rand_exe_prng_15_io_out_8),
    .io_out_9(rand_exe_prng_15_io_out_9),
    .io_out_10(rand_exe_prng_15_io_out_10),
    .io_out_11(rand_exe_prng_15_io_out_11),
    .io_out_12(rand_exe_prng_15_io_out_12),
    .io_out_13(rand_exe_prng_15_io_out_13),
    .io_out_14(rand_exe_prng_15_io_out_14),
    .io_out_15(rand_exe_prng_15_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_16 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_16_clock),
    .reset(rand_exe_prng_16_reset),
    .io_out_0(rand_exe_prng_16_io_out_0),
    .io_out_1(rand_exe_prng_16_io_out_1),
    .io_out_2(rand_exe_prng_16_io_out_2),
    .io_out_3(rand_exe_prng_16_io_out_3),
    .io_out_4(rand_exe_prng_16_io_out_4),
    .io_out_5(rand_exe_prng_16_io_out_5),
    .io_out_6(rand_exe_prng_16_io_out_6),
    .io_out_7(rand_exe_prng_16_io_out_7),
    .io_out_8(rand_exe_prng_16_io_out_8),
    .io_out_9(rand_exe_prng_16_io_out_9),
    .io_out_10(rand_exe_prng_16_io_out_10),
    .io_out_11(rand_exe_prng_16_io_out_11),
    .io_out_12(rand_exe_prng_16_io_out_12),
    .io_out_13(rand_exe_prng_16_io_out_13),
    .io_out_14(rand_exe_prng_16_io_out_14),
    .io_out_15(rand_exe_prng_16_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_17 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_17_clock),
    .reset(rand_exe_prng_17_reset),
    .io_out_0(rand_exe_prng_17_io_out_0),
    .io_out_1(rand_exe_prng_17_io_out_1),
    .io_out_2(rand_exe_prng_17_io_out_2),
    .io_out_3(rand_exe_prng_17_io_out_3),
    .io_out_4(rand_exe_prng_17_io_out_4),
    .io_out_5(rand_exe_prng_17_io_out_5),
    .io_out_6(rand_exe_prng_17_io_out_6),
    .io_out_7(rand_exe_prng_17_io_out_7),
    .io_out_8(rand_exe_prng_17_io_out_8),
    .io_out_9(rand_exe_prng_17_io_out_9),
    .io_out_10(rand_exe_prng_17_io_out_10),
    .io_out_11(rand_exe_prng_17_io_out_11),
    .io_out_12(rand_exe_prng_17_io_out_12),
    .io_out_13(rand_exe_prng_17_io_out_13),
    .io_out_14(rand_exe_prng_17_io_out_14),
    .io_out_15(rand_exe_prng_17_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_18 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_18_clock),
    .reset(rand_exe_prng_18_reset),
    .io_out_0(rand_exe_prng_18_io_out_0),
    .io_out_1(rand_exe_prng_18_io_out_1),
    .io_out_2(rand_exe_prng_18_io_out_2),
    .io_out_3(rand_exe_prng_18_io_out_3),
    .io_out_4(rand_exe_prng_18_io_out_4),
    .io_out_5(rand_exe_prng_18_io_out_5),
    .io_out_6(rand_exe_prng_18_io_out_6),
    .io_out_7(rand_exe_prng_18_io_out_7),
    .io_out_8(rand_exe_prng_18_io_out_8),
    .io_out_9(rand_exe_prng_18_io_out_9),
    .io_out_10(rand_exe_prng_18_io_out_10),
    .io_out_11(rand_exe_prng_18_io_out_11),
    .io_out_12(rand_exe_prng_18_io_out_12),
    .io_out_13(rand_exe_prng_18_io_out_13),
    .io_out_14(rand_exe_prng_18_io_out_14),
    .io_out_15(rand_exe_prng_18_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_19 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_19_clock),
    .reset(rand_exe_prng_19_reset),
    .io_out_0(rand_exe_prng_19_io_out_0),
    .io_out_1(rand_exe_prng_19_io_out_1),
    .io_out_2(rand_exe_prng_19_io_out_2),
    .io_out_3(rand_exe_prng_19_io_out_3),
    .io_out_4(rand_exe_prng_19_io_out_4),
    .io_out_5(rand_exe_prng_19_io_out_5),
    .io_out_6(rand_exe_prng_19_io_out_6),
    .io_out_7(rand_exe_prng_19_io_out_7),
    .io_out_8(rand_exe_prng_19_io_out_8),
    .io_out_9(rand_exe_prng_19_io_out_9),
    .io_out_10(rand_exe_prng_19_io_out_10),
    .io_out_11(rand_exe_prng_19_io_out_11),
    .io_out_12(rand_exe_prng_19_io_out_12),
    .io_out_13(rand_exe_prng_19_io_out_13),
    .io_out_14(rand_exe_prng_19_io_out_14),
    .io_out_15(rand_exe_prng_19_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_20 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_20_clock),
    .reset(rand_exe_prng_20_reset),
    .io_out_0(rand_exe_prng_20_io_out_0),
    .io_out_1(rand_exe_prng_20_io_out_1),
    .io_out_2(rand_exe_prng_20_io_out_2),
    .io_out_3(rand_exe_prng_20_io_out_3),
    .io_out_4(rand_exe_prng_20_io_out_4),
    .io_out_5(rand_exe_prng_20_io_out_5),
    .io_out_6(rand_exe_prng_20_io_out_6),
    .io_out_7(rand_exe_prng_20_io_out_7),
    .io_out_8(rand_exe_prng_20_io_out_8),
    .io_out_9(rand_exe_prng_20_io_out_9),
    .io_out_10(rand_exe_prng_20_io_out_10),
    .io_out_11(rand_exe_prng_20_io_out_11),
    .io_out_12(rand_exe_prng_20_io_out_12),
    .io_out_13(rand_exe_prng_20_io_out_13),
    .io_out_14(rand_exe_prng_20_io_out_14),
    .io_out_15(rand_exe_prng_20_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_21 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_21_clock),
    .reset(rand_exe_prng_21_reset),
    .io_out_0(rand_exe_prng_21_io_out_0),
    .io_out_1(rand_exe_prng_21_io_out_1),
    .io_out_2(rand_exe_prng_21_io_out_2),
    .io_out_3(rand_exe_prng_21_io_out_3),
    .io_out_4(rand_exe_prng_21_io_out_4),
    .io_out_5(rand_exe_prng_21_io_out_5),
    .io_out_6(rand_exe_prng_21_io_out_6),
    .io_out_7(rand_exe_prng_21_io_out_7),
    .io_out_8(rand_exe_prng_21_io_out_8),
    .io_out_9(rand_exe_prng_21_io_out_9),
    .io_out_10(rand_exe_prng_21_io_out_10),
    .io_out_11(rand_exe_prng_21_io_out_11),
    .io_out_12(rand_exe_prng_21_io_out_12),
    .io_out_13(rand_exe_prng_21_io_out_13),
    .io_out_14(rand_exe_prng_21_io_out_14),
    .io_out_15(rand_exe_prng_21_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_22 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_22_clock),
    .reset(rand_exe_prng_22_reset),
    .io_out_0(rand_exe_prng_22_io_out_0),
    .io_out_1(rand_exe_prng_22_io_out_1),
    .io_out_2(rand_exe_prng_22_io_out_2),
    .io_out_3(rand_exe_prng_22_io_out_3),
    .io_out_4(rand_exe_prng_22_io_out_4),
    .io_out_5(rand_exe_prng_22_io_out_5),
    .io_out_6(rand_exe_prng_22_io_out_6),
    .io_out_7(rand_exe_prng_22_io_out_7),
    .io_out_8(rand_exe_prng_22_io_out_8),
    .io_out_9(rand_exe_prng_22_io_out_9),
    .io_out_10(rand_exe_prng_22_io_out_10),
    .io_out_11(rand_exe_prng_22_io_out_11),
    .io_out_12(rand_exe_prng_22_io_out_12),
    .io_out_13(rand_exe_prng_22_io_out_13),
    .io_out_14(rand_exe_prng_22_io_out_14),
    .io_out_15(rand_exe_prng_22_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_23 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_23_clock),
    .reset(rand_exe_prng_23_reset),
    .io_out_0(rand_exe_prng_23_io_out_0),
    .io_out_1(rand_exe_prng_23_io_out_1),
    .io_out_2(rand_exe_prng_23_io_out_2),
    .io_out_3(rand_exe_prng_23_io_out_3),
    .io_out_4(rand_exe_prng_23_io_out_4),
    .io_out_5(rand_exe_prng_23_io_out_5),
    .io_out_6(rand_exe_prng_23_io_out_6),
    .io_out_7(rand_exe_prng_23_io_out_7),
    .io_out_8(rand_exe_prng_23_io_out_8),
    .io_out_9(rand_exe_prng_23_io_out_9),
    .io_out_10(rand_exe_prng_23_io_out_10),
    .io_out_11(rand_exe_prng_23_io_out_11),
    .io_out_12(rand_exe_prng_23_io_out_12),
    .io_out_13(rand_exe_prng_23_io_out_13),
    .io_out_14(rand_exe_prng_23_io_out_14),
    .io_out_15(rand_exe_prng_23_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_24 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_24_clock),
    .reset(rand_exe_prng_24_reset),
    .io_out_0(rand_exe_prng_24_io_out_0),
    .io_out_1(rand_exe_prng_24_io_out_1),
    .io_out_2(rand_exe_prng_24_io_out_2),
    .io_out_3(rand_exe_prng_24_io_out_3),
    .io_out_4(rand_exe_prng_24_io_out_4),
    .io_out_5(rand_exe_prng_24_io_out_5),
    .io_out_6(rand_exe_prng_24_io_out_6),
    .io_out_7(rand_exe_prng_24_io_out_7),
    .io_out_8(rand_exe_prng_24_io_out_8),
    .io_out_9(rand_exe_prng_24_io_out_9),
    .io_out_10(rand_exe_prng_24_io_out_10),
    .io_out_11(rand_exe_prng_24_io_out_11),
    .io_out_12(rand_exe_prng_24_io_out_12),
    .io_out_13(rand_exe_prng_24_io_out_13),
    .io_out_14(rand_exe_prng_24_io_out_14),
    .io_out_15(rand_exe_prng_24_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_25 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_25_clock),
    .reset(rand_exe_prng_25_reset),
    .io_out_0(rand_exe_prng_25_io_out_0),
    .io_out_1(rand_exe_prng_25_io_out_1),
    .io_out_2(rand_exe_prng_25_io_out_2),
    .io_out_3(rand_exe_prng_25_io_out_3),
    .io_out_4(rand_exe_prng_25_io_out_4),
    .io_out_5(rand_exe_prng_25_io_out_5),
    .io_out_6(rand_exe_prng_25_io_out_6),
    .io_out_7(rand_exe_prng_25_io_out_7),
    .io_out_8(rand_exe_prng_25_io_out_8),
    .io_out_9(rand_exe_prng_25_io_out_9),
    .io_out_10(rand_exe_prng_25_io_out_10),
    .io_out_11(rand_exe_prng_25_io_out_11),
    .io_out_12(rand_exe_prng_25_io_out_12),
    .io_out_13(rand_exe_prng_25_io_out_13),
    .io_out_14(rand_exe_prng_25_io_out_14),
    .io_out_15(rand_exe_prng_25_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_26 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_26_clock),
    .reset(rand_exe_prng_26_reset),
    .io_out_0(rand_exe_prng_26_io_out_0),
    .io_out_1(rand_exe_prng_26_io_out_1),
    .io_out_2(rand_exe_prng_26_io_out_2),
    .io_out_3(rand_exe_prng_26_io_out_3),
    .io_out_4(rand_exe_prng_26_io_out_4),
    .io_out_5(rand_exe_prng_26_io_out_5),
    .io_out_6(rand_exe_prng_26_io_out_6),
    .io_out_7(rand_exe_prng_26_io_out_7),
    .io_out_8(rand_exe_prng_26_io_out_8),
    .io_out_9(rand_exe_prng_26_io_out_9),
    .io_out_10(rand_exe_prng_26_io_out_10),
    .io_out_11(rand_exe_prng_26_io_out_11),
    .io_out_12(rand_exe_prng_26_io_out_12),
    .io_out_13(rand_exe_prng_26_io_out_13),
    .io_out_14(rand_exe_prng_26_io_out_14),
    .io_out_15(rand_exe_prng_26_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_27 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_27_clock),
    .reset(rand_exe_prng_27_reset),
    .io_out_0(rand_exe_prng_27_io_out_0),
    .io_out_1(rand_exe_prng_27_io_out_1),
    .io_out_2(rand_exe_prng_27_io_out_2),
    .io_out_3(rand_exe_prng_27_io_out_3),
    .io_out_4(rand_exe_prng_27_io_out_4),
    .io_out_5(rand_exe_prng_27_io_out_5),
    .io_out_6(rand_exe_prng_27_io_out_6),
    .io_out_7(rand_exe_prng_27_io_out_7),
    .io_out_8(rand_exe_prng_27_io_out_8),
    .io_out_9(rand_exe_prng_27_io_out_9),
    .io_out_10(rand_exe_prng_27_io_out_10),
    .io_out_11(rand_exe_prng_27_io_out_11),
    .io_out_12(rand_exe_prng_27_io_out_12),
    .io_out_13(rand_exe_prng_27_io_out_13),
    .io_out_14(rand_exe_prng_27_io_out_14),
    .io_out_15(rand_exe_prng_27_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_28 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_28_clock),
    .reset(rand_exe_prng_28_reset),
    .io_out_0(rand_exe_prng_28_io_out_0),
    .io_out_1(rand_exe_prng_28_io_out_1),
    .io_out_2(rand_exe_prng_28_io_out_2),
    .io_out_3(rand_exe_prng_28_io_out_3),
    .io_out_4(rand_exe_prng_28_io_out_4),
    .io_out_5(rand_exe_prng_28_io_out_5),
    .io_out_6(rand_exe_prng_28_io_out_6),
    .io_out_7(rand_exe_prng_28_io_out_7),
    .io_out_8(rand_exe_prng_28_io_out_8),
    .io_out_9(rand_exe_prng_28_io_out_9),
    .io_out_10(rand_exe_prng_28_io_out_10),
    .io_out_11(rand_exe_prng_28_io_out_11),
    .io_out_12(rand_exe_prng_28_io_out_12),
    .io_out_13(rand_exe_prng_28_io_out_13),
    .io_out_14(rand_exe_prng_28_io_out_14),
    .io_out_15(rand_exe_prng_28_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_29 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_29_clock),
    .reset(rand_exe_prng_29_reset),
    .io_out_0(rand_exe_prng_29_io_out_0),
    .io_out_1(rand_exe_prng_29_io_out_1),
    .io_out_2(rand_exe_prng_29_io_out_2),
    .io_out_3(rand_exe_prng_29_io_out_3),
    .io_out_4(rand_exe_prng_29_io_out_4),
    .io_out_5(rand_exe_prng_29_io_out_5),
    .io_out_6(rand_exe_prng_29_io_out_6),
    .io_out_7(rand_exe_prng_29_io_out_7),
    .io_out_8(rand_exe_prng_29_io_out_8),
    .io_out_9(rand_exe_prng_29_io_out_9),
    .io_out_10(rand_exe_prng_29_io_out_10),
    .io_out_11(rand_exe_prng_29_io_out_11),
    .io_out_12(rand_exe_prng_29_io_out_12),
    .io_out_13(rand_exe_prng_29_io_out_13),
    .io_out_14(rand_exe_prng_29_io_out_14),
    .io_out_15(rand_exe_prng_29_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_30 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_30_clock),
    .reset(rand_exe_prng_30_reset),
    .io_out_0(rand_exe_prng_30_io_out_0),
    .io_out_1(rand_exe_prng_30_io_out_1),
    .io_out_2(rand_exe_prng_30_io_out_2),
    .io_out_3(rand_exe_prng_30_io_out_3),
    .io_out_4(rand_exe_prng_30_io_out_4),
    .io_out_5(rand_exe_prng_30_io_out_5),
    .io_out_6(rand_exe_prng_30_io_out_6),
    .io_out_7(rand_exe_prng_30_io_out_7),
    .io_out_8(rand_exe_prng_30_io_out_8),
    .io_out_9(rand_exe_prng_30_io_out_9),
    .io_out_10(rand_exe_prng_30_io_out_10),
    .io_out_11(rand_exe_prng_30_io_out_11),
    .io_out_12(rand_exe_prng_30_io_out_12),
    .io_out_13(rand_exe_prng_30_io_out_13),
    .io_out_14(rand_exe_prng_30_io_out_14),
    .io_out_15(rand_exe_prng_30_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_31 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_31_clock),
    .reset(rand_exe_prng_31_reset),
    .io_out_0(rand_exe_prng_31_io_out_0),
    .io_out_1(rand_exe_prng_31_io_out_1),
    .io_out_2(rand_exe_prng_31_io_out_2),
    .io_out_3(rand_exe_prng_31_io_out_3),
    .io_out_4(rand_exe_prng_31_io_out_4),
    .io_out_5(rand_exe_prng_31_io_out_5),
    .io_out_6(rand_exe_prng_31_io_out_6),
    .io_out_7(rand_exe_prng_31_io_out_7),
    .io_out_8(rand_exe_prng_31_io_out_8),
    .io_out_9(rand_exe_prng_31_io_out_9),
    .io_out_10(rand_exe_prng_31_io_out_10),
    .io_out_11(rand_exe_prng_31_io_out_11),
    .io_out_12(rand_exe_prng_31_io_out_12),
    .io_out_13(rand_exe_prng_31_io_out_13),
    .io_out_14(rand_exe_prng_31_io_out_14),
    .io_out_15(rand_exe_prng_31_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_32 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_32_clock),
    .reset(rand_exe_prng_32_reset),
    .io_out_0(rand_exe_prng_32_io_out_0),
    .io_out_1(rand_exe_prng_32_io_out_1),
    .io_out_2(rand_exe_prng_32_io_out_2),
    .io_out_3(rand_exe_prng_32_io_out_3),
    .io_out_4(rand_exe_prng_32_io_out_4),
    .io_out_5(rand_exe_prng_32_io_out_5),
    .io_out_6(rand_exe_prng_32_io_out_6),
    .io_out_7(rand_exe_prng_32_io_out_7),
    .io_out_8(rand_exe_prng_32_io_out_8),
    .io_out_9(rand_exe_prng_32_io_out_9),
    .io_out_10(rand_exe_prng_32_io_out_10),
    .io_out_11(rand_exe_prng_32_io_out_11),
    .io_out_12(rand_exe_prng_32_io_out_12),
    .io_out_13(rand_exe_prng_32_io_out_13),
    .io_out_14(rand_exe_prng_32_io_out_14),
    .io_out_15(rand_exe_prng_32_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_33 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_33_clock),
    .reset(rand_exe_prng_33_reset),
    .io_out_0(rand_exe_prng_33_io_out_0),
    .io_out_1(rand_exe_prng_33_io_out_1),
    .io_out_2(rand_exe_prng_33_io_out_2),
    .io_out_3(rand_exe_prng_33_io_out_3),
    .io_out_4(rand_exe_prng_33_io_out_4),
    .io_out_5(rand_exe_prng_33_io_out_5),
    .io_out_6(rand_exe_prng_33_io_out_6),
    .io_out_7(rand_exe_prng_33_io_out_7),
    .io_out_8(rand_exe_prng_33_io_out_8),
    .io_out_9(rand_exe_prng_33_io_out_9),
    .io_out_10(rand_exe_prng_33_io_out_10),
    .io_out_11(rand_exe_prng_33_io_out_11),
    .io_out_12(rand_exe_prng_33_io_out_12),
    .io_out_13(rand_exe_prng_33_io_out_13),
    .io_out_14(rand_exe_prng_33_io_out_14),
    .io_out_15(rand_exe_prng_33_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_34 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_34_clock),
    .reset(rand_exe_prng_34_reset),
    .io_out_0(rand_exe_prng_34_io_out_0),
    .io_out_1(rand_exe_prng_34_io_out_1),
    .io_out_2(rand_exe_prng_34_io_out_2),
    .io_out_3(rand_exe_prng_34_io_out_3),
    .io_out_4(rand_exe_prng_34_io_out_4),
    .io_out_5(rand_exe_prng_34_io_out_5),
    .io_out_6(rand_exe_prng_34_io_out_6),
    .io_out_7(rand_exe_prng_34_io_out_7),
    .io_out_8(rand_exe_prng_34_io_out_8),
    .io_out_9(rand_exe_prng_34_io_out_9),
    .io_out_10(rand_exe_prng_34_io_out_10),
    .io_out_11(rand_exe_prng_34_io_out_11),
    .io_out_12(rand_exe_prng_34_io_out_12),
    .io_out_13(rand_exe_prng_34_io_out_13),
    .io_out_14(rand_exe_prng_34_io_out_14),
    .io_out_15(rand_exe_prng_34_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_35 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_35_clock),
    .reset(rand_exe_prng_35_reset),
    .io_out_0(rand_exe_prng_35_io_out_0),
    .io_out_1(rand_exe_prng_35_io_out_1),
    .io_out_2(rand_exe_prng_35_io_out_2),
    .io_out_3(rand_exe_prng_35_io_out_3),
    .io_out_4(rand_exe_prng_35_io_out_4),
    .io_out_5(rand_exe_prng_35_io_out_5),
    .io_out_6(rand_exe_prng_35_io_out_6),
    .io_out_7(rand_exe_prng_35_io_out_7),
    .io_out_8(rand_exe_prng_35_io_out_8),
    .io_out_9(rand_exe_prng_35_io_out_9),
    .io_out_10(rand_exe_prng_35_io_out_10),
    .io_out_11(rand_exe_prng_35_io_out_11),
    .io_out_12(rand_exe_prng_35_io_out_12),
    .io_out_13(rand_exe_prng_35_io_out_13),
    .io_out_14(rand_exe_prng_35_io_out_14),
    .io_out_15(rand_exe_prng_35_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_36 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_36_clock),
    .reset(rand_exe_prng_36_reset),
    .io_out_0(rand_exe_prng_36_io_out_0),
    .io_out_1(rand_exe_prng_36_io_out_1),
    .io_out_2(rand_exe_prng_36_io_out_2),
    .io_out_3(rand_exe_prng_36_io_out_3),
    .io_out_4(rand_exe_prng_36_io_out_4),
    .io_out_5(rand_exe_prng_36_io_out_5),
    .io_out_6(rand_exe_prng_36_io_out_6),
    .io_out_7(rand_exe_prng_36_io_out_7),
    .io_out_8(rand_exe_prng_36_io_out_8),
    .io_out_9(rand_exe_prng_36_io_out_9),
    .io_out_10(rand_exe_prng_36_io_out_10),
    .io_out_11(rand_exe_prng_36_io_out_11),
    .io_out_12(rand_exe_prng_36_io_out_12),
    .io_out_13(rand_exe_prng_36_io_out_13),
    .io_out_14(rand_exe_prng_36_io_out_14),
    .io_out_15(rand_exe_prng_36_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_37 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_37_clock),
    .reset(rand_exe_prng_37_reset),
    .io_out_0(rand_exe_prng_37_io_out_0),
    .io_out_1(rand_exe_prng_37_io_out_1),
    .io_out_2(rand_exe_prng_37_io_out_2),
    .io_out_3(rand_exe_prng_37_io_out_3),
    .io_out_4(rand_exe_prng_37_io_out_4),
    .io_out_5(rand_exe_prng_37_io_out_5),
    .io_out_6(rand_exe_prng_37_io_out_6),
    .io_out_7(rand_exe_prng_37_io_out_7),
    .io_out_8(rand_exe_prng_37_io_out_8),
    .io_out_9(rand_exe_prng_37_io_out_9),
    .io_out_10(rand_exe_prng_37_io_out_10),
    .io_out_11(rand_exe_prng_37_io_out_11),
    .io_out_12(rand_exe_prng_37_io_out_12),
    .io_out_13(rand_exe_prng_37_io_out_13),
    .io_out_14(rand_exe_prng_37_io_out_14),
    .io_out_15(rand_exe_prng_37_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_38 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_38_clock),
    .reset(rand_exe_prng_38_reset),
    .io_out_0(rand_exe_prng_38_io_out_0),
    .io_out_1(rand_exe_prng_38_io_out_1),
    .io_out_2(rand_exe_prng_38_io_out_2),
    .io_out_3(rand_exe_prng_38_io_out_3),
    .io_out_4(rand_exe_prng_38_io_out_4),
    .io_out_5(rand_exe_prng_38_io_out_5),
    .io_out_6(rand_exe_prng_38_io_out_6),
    .io_out_7(rand_exe_prng_38_io_out_7),
    .io_out_8(rand_exe_prng_38_io_out_8),
    .io_out_9(rand_exe_prng_38_io_out_9),
    .io_out_10(rand_exe_prng_38_io_out_10),
    .io_out_11(rand_exe_prng_38_io_out_11),
    .io_out_12(rand_exe_prng_38_io_out_12),
    .io_out_13(rand_exe_prng_38_io_out_13),
    .io_out_14(rand_exe_prng_38_io_out_14),
    .io_out_15(rand_exe_prng_38_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_39 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_39_clock),
    .reset(rand_exe_prng_39_reset),
    .io_out_0(rand_exe_prng_39_io_out_0),
    .io_out_1(rand_exe_prng_39_io_out_1),
    .io_out_2(rand_exe_prng_39_io_out_2),
    .io_out_3(rand_exe_prng_39_io_out_3),
    .io_out_4(rand_exe_prng_39_io_out_4),
    .io_out_5(rand_exe_prng_39_io_out_5),
    .io_out_6(rand_exe_prng_39_io_out_6),
    .io_out_7(rand_exe_prng_39_io_out_7),
    .io_out_8(rand_exe_prng_39_io_out_8),
    .io_out_9(rand_exe_prng_39_io_out_9),
    .io_out_10(rand_exe_prng_39_io_out_10),
    .io_out_11(rand_exe_prng_39_io_out_11),
    .io_out_12(rand_exe_prng_39_io_out_12),
    .io_out_13(rand_exe_prng_39_io_out_13),
    .io_out_14(rand_exe_prng_39_io_out_14),
    .io_out_15(rand_exe_prng_39_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_40 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_40_clock),
    .reset(rand_exe_prng_40_reset),
    .io_out_0(rand_exe_prng_40_io_out_0),
    .io_out_1(rand_exe_prng_40_io_out_1),
    .io_out_2(rand_exe_prng_40_io_out_2),
    .io_out_3(rand_exe_prng_40_io_out_3),
    .io_out_4(rand_exe_prng_40_io_out_4),
    .io_out_5(rand_exe_prng_40_io_out_5),
    .io_out_6(rand_exe_prng_40_io_out_6),
    .io_out_7(rand_exe_prng_40_io_out_7),
    .io_out_8(rand_exe_prng_40_io_out_8),
    .io_out_9(rand_exe_prng_40_io_out_9),
    .io_out_10(rand_exe_prng_40_io_out_10),
    .io_out_11(rand_exe_prng_40_io_out_11),
    .io_out_12(rand_exe_prng_40_io_out_12),
    .io_out_13(rand_exe_prng_40_io_out_13),
    .io_out_14(rand_exe_prng_40_io_out_14),
    .io_out_15(rand_exe_prng_40_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_41 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_41_clock),
    .reset(rand_exe_prng_41_reset),
    .io_out_0(rand_exe_prng_41_io_out_0),
    .io_out_1(rand_exe_prng_41_io_out_1),
    .io_out_2(rand_exe_prng_41_io_out_2),
    .io_out_3(rand_exe_prng_41_io_out_3),
    .io_out_4(rand_exe_prng_41_io_out_4),
    .io_out_5(rand_exe_prng_41_io_out_5),
    .io_out_6(rand_exe_prng_41_io_out_6),
    .io_out_7(rand_exe_prng_41_io_out_7),
    .io_out_8(rand_exe_prng_41_io_out_8),
    .io_out_9(rand_exe_prng_41_io_out_9),
    .io_out_10(rand_exe_prng_41_io_out_10),
    .io_out_11(rand_exe_prng_41_io_out_11),
    .io_out_12(rand_exe_prng_41_io_out_12),
    .io_out_13(rand_exe_prng_41_io_out_13),
    .io_out_14(rand_exe_prng_41_io_out_14),
    .io_out_15(rand_exe_prng_41_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_42 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_42_clock),
    .reset(rand_exe_prng_42_reset),
    .io_out_0(rand_exe_prng_42_io_out_0),
    .io_out_1(rand_exe_prng_42_io_out_1),
    .io_out_2(rand_exe_prng_42_io_out_2),
    .io_out_3(rand_exe_prng_42_io_out_3),
    .io_out_4(rand_exe_prng_42_io_out_4),
    .io_out_5(rand_exe_prng_42_io_out_5),
    .io_out_6(rand_exe_prng_42_io_out_6),
    .io_out_7(rand_exe_prng_42_io_out_7),
    .io_out_8(rand_exe_prng_42_io_out_8),
    .io_out_9(rand_exe_prng_42_io_out_9),
    .io_out_10(rand_exe_prng_42_io_out_10),
    .io_out_11(rand_exe_prng_42_io_out_11),
    .io_out_12(rand_exe_prng_42_io_out_12),
    .io_out_13(rand_exe_prng_42_io_out_13),
    .io_out_14(rand_exe_prng_42_io_out_14),
    .io_out_15(rand_exe_prng_42_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_43 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_43_clock),
    .reset(rand_exe_prng_43_reset),
    .io_out_0(rand_exe_prng_43_io_out_0),
    .io_out_1(rand_exe_prng_43_io_out_1),
    .io_out_2(rand_exe_prng_43_io_out_2),
    .io_out_3(rand_exe_prng_43_io_out_3),
    .io_out_4(rand_exe_prng_43_io_out_4),
    .io_out_5(rand_exe_prng_43_io_out_5),
    .io_out_6(rand_exe_prng_43_io_out_6),
    .io_out_7(rand_exe_prng_43_io_out_7),
    .io_out_8(rand_exe_prng_43_io_out_8),
    .io_out_9(rand_exe_prng_43_io_out_9),
    .io_out_10(rand_exe_prng_43_io_out_10),
    .io_out_11(rand_exe_prng_43_io_out_11),
    .io_out_12(rand_exe_prng_43_io_out_12),
    .io_out_13(rand_exe_prng_43_io_out_13),
    .io_out_14(rand_exe_prng_43_io_out_14),
    .io_out_15(rand_exe_prng_43_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_44 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_44_clock),
    .reset(rand_exe_prng_44_reset),
    .io_out_0(rand_exe_prng_44_io_out_0),
    .io_out_1(rand_exe_prng_44_io_out_1),
    .io_out_2(rand_exe_prng_44_io_out_2),
    .io_out_3(rand_exe_prng_44_io_out_3),
    .io_out_4(rand_exe_prng_44_io_out_4),
    .io_out_5(rand_exe_prng_44_io_out_5),
    .io_out_6(rand_exe_prng_44_io_out_6),
    .io_out_7(rand_exe_prng_44_io_out_7),
    .io_out_8(rand_exe_prng_44_io_out_8),
    .io_out_9(rand_exe_prng_44_io_out_9),
    .io_out_10(rand_exe_prng_44_io_out_10),
    .io_out_11(rand_exe_prng_44_io_out_11),
    .io_out_12(rand_exe_prng_44_io_out_12),
    .io_out_13(rand_exe_prng_44_io_out_13),
    .io_out_14(rand_exe_prng_44_io_out_14),
    .io_out_15(rand_exe_prng_44_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_45 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_45_clock),
    .reset(rand_exe_prng_45_reset),
    .io_out_0(rand_exe_prng_45_io_out_0),
    .io_out_1(rand_exe_prng_45_io_out_1),
    .io_out_2(rand_exe_prng_45_io_out_2),
    .io_out_3(rand_exe_prng_45_io_out_3),
    .io_out_4(rand_exe_prng_45_io_out_4),
    .io_out_5(rand_exe_prng_45_io_out_5),
    .io_out_6(rand_exe_prng_45_io_out_6),
    .io_out_7(rand_exe_prng_45_io_out_7),
    .io_out_8(rand_exe_prng_45_io_out_8),
    .io_out_9(rand_exe_prng_45_io_out_9),
    .io_out_10(rand_exe_prng_45_io_out_10),
    .io_out_11(rand_exe_prng_45_io_out_11),
    .io_out_12(rand_exe_prng_45_io_out_12),
    .io_out_13(rand_exe_prng_45_io_out_13),
    .io_out_14(rand_exe_prng_45_io_out_14),
    .io_out_15(rand_exe_prng_45_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_46 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_46_clock),
    .reset(rand_exe_prng_46_reset),
    .io_out_0(rand_exe_prng_46_io_out_0),
    .io_out_1(rand_exe_prng_46_io_out_1),
    .io_out_2(rand_exe_prng_46_io_out_2),
    .io_out_3(rand_exe_prng_46_io_out_3),
    .io_out_4(rand_exe_prng_46_io_out_4),
    .io_out_5(rand_exe_prng_46_io_out_5),
    .io_out_6(rand_exe_prng_46_io_out_6),
    .io_out_7(rand_exe_prng_46_io_out_7),
    .io_out_8(rand_exe_prng_46_io_out_8),
    .io_out_9(rand_exe_prng_46_io_out_9),
    .io_out_10(rand_exe_prng_46_io_out_10),
    .io_out_11(rand_exe_prng_46_io_out_11),
    .io_out_12(rand_exe_prng_46_io_out_12),
    .io_out_13(rand_exe_prng_46_io_out_13),
    .io_out_14(rand_exe_prng_46_io_out_14),
    .io_out_15(rand_exe_prng_46_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_47 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_47_clock),
    .reset(rand_exe_prng_47_reset),
    .io_out_0(rand_exe_prng_47_io_out_0),
    .io_out_1(rand_exe_prng_47_io_out_1),
    .io_out_2(rand_exe_prng_47_io_out_2),
    .io_out_3(rand_exe_prng_47_io_out_3),
    .io_out_4(rand_exe_prng_47_io_out_4),
    .io_out_5(rand_exe_prng_47_io_out_5),
    .io_out_6(rand_exe_prng_47_io_out_6),
    .io_out_7(rand_exe_prng_47_io_out_7),
    .io_out_8(rand_exe_prng_47_io_out_8),
    .io_out_9(rand_exe_prng_47_io_out_9),
    .io_out_10(rand_exe_prng_47_io_out_10),
    .io_out_11(rand_exe_prng_47_io_out_11),
    .io_out_12(rand_exe_prng_47_io_out_12),
    .io_out_13(rand_exe_prng_47_io_out_13),
    .io_out_14(rand_exe_prng_47_io_out_14),
    .io_out_15(rand_exe_prng_47_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_48 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_48_clock),
    .reset(rand_exe_prng_48_reset),
    .io_out_0(rand_exe_prng_48_io_out_0),
    .io_out_1(rand_exe_prng_48_io_out_1),
    .io_out_2(rand_exe_prng_48_io_out_2),
    .io_out_3(rand_exe_prng_48_io_out_3),
    .io_out_4(rand_exe_prng_48_io_out_4),
    .io_out_5(rand_exe_prng_48_io_out_5),
    .io_out_6(rand_exe_prng_48_io_out_6),
    .io_out_7(rand_exe_prng_48_io_out_7),
    .io_out_8(rand_exe_prng_48_io_out_8),
    .io_out_9(rand_exe_prng_48_io_out_9),
    .io_out_10(rand_exe_prng_48_io_out_10),
    .io_out_11(rand_exe_prng_48_io_out_11),
    .io_out_12(rand_exe_prng_48_io_out_12),
    .io_out_13(rand_exe_prng_48_io_out_13),
    .io_out_14(rand_exe_prng_48_io_out_14),
    .io_out_15(rand_exe_prng_48_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_49 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_49_clock),
    .reset(rand_exe_prng_49_reset),
    .io_out_0(rand_exe_prng_49_io_out_0),
    .io_out_1(rand_exe_prng_49_io_out_1),
    .io_out_2(rand_exe_prng_49_io_out_2),
    .io_out_3(rand_exe_prng_49_io_out_3),
    .io_out_4(rand_exe_prng_49_io_out_4),
    .io_out_5(rand_exe_prng_49_io_out_5),
    .io_out_6(rand_exe_prng_49_io_out_6),
    .io_out_7(rand_exe_prng_49_io_out_7),
    .io_out_8(rand_exe_prng_49_io_out_8),
    .io_out_9(rand_exe_prng_49_io_out_9),
    .io_out_10(rand_exe_prng_49_io_out_10),
    .io_out_11(rand_exe_prng_49_io_out_11),
    .io_out_12(rand_exe_prng_49_io_out_12),
    .io_out_13(rand_exe_prng_49_io_out_13),
    .io_out_14(rand_exe_prng_49_io_out_14),
    .io_out_15(rand_exe_prng_49_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_50 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_50_clock),
    .reset(rand_exe_prng_50_reset),
    .io_out_0(rand_exe_prng_50_io_out_0),
    .io_out_1(rand_exe_prng_50_io_out_1),
    .io_out_2(rand_exe_prng_50_io_out_2),
    .io_out_3(rand_exe_prng_50_io_out_3),
    .io_out_4(rand_exe_prng_50_io_out_4),
    .io_out_5(rand_exe_prng_50_io_out_5),
    .io_out_6(rand_exe_prng_50_io_out_6),
    .io_out_7(rand_exe_prng_50_io_out_7),
    .io_out_8(rand_exe_prng_50_io_out_8),
    .io_out_9(rand_exe_prng_50_io_out_9),
    .io_out_10(rand_exe_prng_50_io_out_10),
    .io_out_11(rand_exe_prng_50_io_out_11),
    .io_out_12(rand_exe_prng_50_io_out_12),
    .io_out_13(rand_exe_prng_50_io_out_13),
    .io_out_14(rand_exe_prng_50_io_out_14),
    .io_out_15(rand_exe_prng_50_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_51 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_51_clock),
    .reset(rand_exe_prng_51_reset),
    .io_out_0(rand_exe_prng_51_io_out_0),
    .io_out_1(rand_exe_prng_51_io_out_1),
    .io_out_2(rand_exe_prng_51_io_out_2),
    .io_out_3(rand_exe_prng_51_io_out_3),
    .io_out_4(rand_exe_prng_51_io_out_4),
    .io_out_5(rand_exe_prng_51_io_out_5),
    .io_out_6(rand_exe_prng_51_io_out_6),
    .io_out_7(rand_exe_prng_51_io_out_7),
    .io_out_8(rand_exe_prng_51_io_out_8),
    .io_out_9(rand_exe_prng_51_io_out_9),
    .io_out_10(rand_exe_prng_51_io_out_10),
    .io_out_11(rand_exe_prng_51_io_out_11),
    .io_out_12(rand_exe_prng_51_io_out_12),
    .io_out_13(rand_exe_prng_51_io_out_13),
    .io_out_14(rand_exe_prng_51_io_out_14),
    .io_out_15(rand_exe_prng_51_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_52 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_52_clock),
    .reset(rand_exe_prng_52_reset),
    .io_out_0(rand_exe_prng_52_io_out_0),
    .io_out_1(rand_exe_prng_52_io_out_1),
    .io_out_2(rand_exe_prng_52_io_out_2),
    .io_out_3(rand_exe_prng_52_io_out_3),
    .io_out_4(rand_exe_prng_52_io_out_4),
    .io_out_5(rand_exe_prng_52_io_out_5),
    .io_out_6(rand_exe_prng_52_io_out_6),
    .io_out_7(rand_exe_prng_52_io_out_7),
    .io_out_8(rand_exe_prng_52_io_out_8),
    .io_out_9(rand_exe_prng_52_io_out_9),
    .io_out_10(rand_exe_prng_52_io_out_10),
    .io_out_11(rand_exe_prng_52_io_out_11),
    .io_out_12(rand_exe_prng_52_io_out_12),
    .io_out_13(rand_exe_prng_52_io_out_13),
    .io_out_14(rand_exe_prng_52_io_out_14),
    .io_out_15(rand_exe_prng_52_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_53 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_53_clock),
    .reset(rand_exe_prng_53_reset),
    .io_out_0(rand_exe_prng_53_io_out_0),
    .io_out_1(rand_exe_prng_53_io_out_1),
    .io_out_2(rand_exe_prng_53_io_out_2),
    .io_out_3(rand_exe_prng_53_io_out_3),
    .io_out_4(rand_exe_prng_53_io_out_4),
    .io_out_5(rand_exe_prng_53_io_out_5),
    .io_out_6(rand_exe_prng_53_io_out_6),
    .io_out_7(rand_exe_prng_53_io_out_7),
    .io_out_8(rand_exe_prng_53_io_out_8),
    .io_out_9(rand_exe_prng_53_io_out_9),
    .io_out_10(rand_exe_prng_53_io_out_10),
    .io_out_11(rand_exe_prng_53_io_out_11),
    .io_out_12(rand_exe_prng_53_io_out_12),
    .io_out_13(rand_exe_prng_53_io_out_13),
    .io_out_14(rand_exe_prng_53_io_out_14),
    .io_out_15(rand_exe_prng_53_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_54 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_54_clock),
    .reset(rand_exe_prng_54_reset),
    .io_out_0(rand_exe_prng_54_io_out_0),
    .io_out_1(rand_exe_prng_54_io_out_1),
    .io_out_2(rand_exe_prng_54_io_out_2),
    .io_out_3(rand_exe_prng_54_io_out_3),
    .io_out_4(rand_exe_prng_54_io_out_4),
    .io_out_5(rand_exe_prng_54_io_out_5),
    .io_out_6(rand_exe_prng_54_io_out_6),
    .io_out_7(rand_exe_prng_54_io_out_7),
    .io_out_8(rand_exe_prng_54_io_out_8),
    .io_out_9(rand_exe_prng_54_io_out_9),
    .io_out_10(rand_exe_prng_54_io_out_10),
    .io_out_11(rand_exe_prng_54_io_out_11),
    .io_out_12(rand_exe_prng_54_io_out_12),
    .io_out_13(rand_exe_prng_54_io_out_13),
    .io_out_14(rand_exe_prng_54_io_out_14),
    .io_out_15(rand_exe_prng_54_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_55 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_55_clock),
    .reset(rand_exe_prng_55_reset),
    .io_out_0(rand_exe_prng_55_io_out_0),
    .io_out_1(rand_exe_prng_55_io_out_1),
    .io_out_2(rand_exe_prng_55_io_out_2),
    .io_out_3(rand_exe_prng_55_io_out_3),
    .io_out_4(rand_exe_prng_55_io_out_4),
    .io_out_5(rand_exe_prng_55_io_out_5),
    .io_out_6(rand_exe_prng_55_io_out_6),
    .io_out_7(rand_exe_prng_55_io_out_7),
    .io_out_8(rand_exe_prng_55_io_out_8),
    .io_out_9(rand_exe_prng_55_io_out_9),
    .io_out_10(rand_exe_prng_55_io_out_10),
    .io_out_11(rand_exe_prng_55_io_out_11),
    .io_out_12(rand_exe_prng_55_io_out_12),
    .io_out_13(rand_exe_prng_55_io_out_13),
    .io_out_14(rand_exe_prng_55_io_out_14),
    .io_out_15(rand_exe_prng_55_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_56 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_56_clock),
    .reset(rand_exe_prng_56_reset),
    .io_out_0(rand_exe_prng_56_io_out_0),
    .io_out_1(rand_exe_prng_56_io_out_1),
    .io_out_2(rand_exe_prng_56_io_out_2),
    .io_out_3(rand_exe_prng_56_io_out_3),
    .io_out_4(rand_exe_prng_56_io_out_4),
    .io_out_5(rand_exe_prng_56_io_out_5),
    .io_out_6(rand_exe_prng_56_io_out_6),
    .io_out_7(rand_exe_prng_56_io_out_7),
    .io_out_8(rand_exe_prng_56_io_out_8),
    .io_out_9(rand_exe_prng_56_io_out_9),
    .io_out_10(rand_exe_prng_56_io_out_10),
    .io_out_11(rand_exe_prng_56_io_out_11),
    .io_out_12(rand_exe_prng_56_io_out_12),
    .io_out_13(rand_exe_prng_56_io_out_13),
    .io_out_14(rand_exe_prng_56_io_out_14),
    .io_out_15(rand_exe_prng_56_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_57 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_57_clock),
    .reset(rand_exe_prng_57_reset),
    .io_out_0(rand_exe_prng_57_io_out_0),
    .io_out_1(rand_exe_prng_57_io_out_1),
    .io_out_2(rand_exe_prng_57_io_out_2),
    .io_out_3(rand_exe_prng_57_io_out_3),
    .io_out_4(rand_exe_prng_57_io_out_4),
    .io_out_5(rand_exe_prng_57_io_out_5),
    .io_out_6(rand_exe_prng_57_io_out_6),
    .io_out_7(rand_exe_prng_57_io_out_7),
    .io_out_8(rand_exe_prng_57_io_out_8),
    .io_out_9(rand_exe_prng_57_io_out_9),
    .io_out_10(rand_exe_prng_57_io_out_10),
    .io_out_11(rand_exe_prng_57_io_out_11),
    .io_out_12(rand_exe_prng_57_io_out_12),
    .io_out_13(rand_exe_prng_57_io_out_13),
    .io_out_14(rand_exe_prng_57_io_out_14),
    .io_out_15(rand_exe_prng_57_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_58 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_58_clock),
    .reset(rand_exe_prng_58_reset),
    .io_out_0(rand_exe_prng_58_io_out_0),
    .io_out_1(rand_exe_prng_58_io_out_1),
    .io_out_2(rand_exe_prng_58_io_out_2),
    .io_out_3(rand_exe_prng_58_io_out_3),
    .io_out_4(rand_exe_prng_58_io_out_4),
    .io_out_5(rand_exe_prng_58_io_out_5),
    .io_out_6(rand_exe_prng_58_io_out_6),
    .io_out_7(rand_exe_prng_58_io_out_7),
    .io_out_8(rand_exe_prng_58_io_out_8),
    .io_out_9(rand_exe_prng_58_io_out_9),
    .io_out_10(rand_exe_prng_58_io_out_10),
    .io_out_11(rand_exe_prng_58_io_out_11),
    .io_out_12(rand_exe_prng_58_io_out_12),
    .io_out_13(rand_exe_prng_58_io_out_13),
    .io_out_14(rand_exe_prng_58_io_out_14),
    .io_out_15(rand_exe_prng_58_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_59 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_59_clock),
    .reset(rand_exe_prng_59_reset),
    .io_out_0(rand_exe_prng_59_io_out_0),
    .io_out_1(rand_exe_prng_59_io_out_1),
    .io_out_2(rand_exe_prng_59_io_out_2),
    .io_out_3(rand_exe_prng_59_io_out_3),
    .io_out_4(rand_exe_prng_59_io_out_4),
    .io_out_5(rand_exe_prng_59_io_out_5),
    .io_out_6(rand_exe_prng_59_io_out_6),
    .io_out_7(rand_exe_prng_59_io_out_7),
    .io_out_8(rand_exe_prng_59_io_out_8),
    .io_out_9(rand_exe_prng_59_io_out_9),
    .io_out_10(rand_exe_prng_59_io_out_10),
    .io_out_11(rand_exe_prng_59_io_out_11),
    .io_out_12(rand_exe_prng_59_io_out_12),
    .io_out_13(rand_exe_prng_59_io_out_13),
    .io_out_14(rand_exe_prng_59_io_out_14),
    .io_out_15(rand_exe_prng_59_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_60 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_60_clock),
    .reset(rand_exe_prng_60_reset),
    .io_out_0(rand_exe_prng_60_io_out_0),
    .io_out_1(rand_exe_prng_60_io_out_1),
    .io_out_2(rand_exe_prng_60_io_out_2),
    .io_out_3(rand_exe_prng_60_io_out_3),
    .io_out_4(rand_exe_prng_60_io_out_4),
    .io_out_5(rand_exe_prng_60_io_out_5),
    .io_out_6(rand_exe_prng_60_io_out_6),
    .io_out_7(rand_exe_prng_60_io_out_7),
    .io_out_8(rand_exe_prng_60_io_out_8),
    .io_out_9(rand_exe_prng_60_io_out_9),
    .io_out_10(rand_exe_prng_60_io_out_10),
    .io_out_11(rand_exe_prng_60_io_out_11),
    .io_out_12(rand_exe_prng_60_io_out_12),
    .io_out_13(rand_exe_prng_60_io_out_13),
    .io_out_14(rand_exe_prng_60_io_out_14),
    .io_out_15(rand_exe_prng_60_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_61 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_61_clock),
    .reset(rand_exe_prng_61_reset),
    .io_out_0(rand_exe_prng_61_io_out_0),
    .io_out_1(rand_exe_prng_61_io_out_1),
    .io_out_2(rand_exe_prng_61_io_out_2),
    .io_out_3(rand_exe_prng_61_io_out_3),
    .io_out_4(rand_exe_prng_61_io_out_4),
    .io_out_5(rand_exe_prng_61_io_out_5),
    .io_out_6(rand_exe_prng_61_io_out_6),
    .io_out_7(rand_exe_prng_61_io_out_7),
    .io_out_8(rand_exe_prng_61_io_out_8),
    .io_out_9(rand_exe_prng_61_io_out_9),
    .io_out_10(rand_exe_prng_61_io_out_10),
    .io_out_11(rand_exe_prng_61_io_out_11),
    .io_out_12(rand_exe_prng_61_io_out_12),
    .io_out_13(rand_exe_prng_61_io_out_13),
    .io_out_14(rand_exe_prng_61_io_out_14),
    .io_out_15(rand_exe_prng_61_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_62 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_62_clock),
    .reset(rand_exe_prng_62_reset),
    .io_out_0(rand_exe_prng_62_io_out_0),
    .io_out_1(rand_exe_prng_62_io_out_1),
    .io_out_2(rand_exe_prng_62_io_out_2),
    .io_out_3(rand_exe_prng_62_io_out_3),
    .io_out_4(rand_exe_prng_62_io_out_4),
    .io_out_5(rand_exe_prng_62_io_out_5),
    .io_out_6(rand_exe_prng_62_io_out_6),
    .io_out_7(rand_exe_prng_62_io_out_7),
    .io_out_8(rand_exe_prng_62_io_out_8),
    .io_out_9(rand_exe_prng_62_io_out_9),
    .io_out_10(rand_exe_prng_62_io_out_10),
    .io_out_11(rand_exe_prng_62_io_out_11),
    .io_out_12(rand_exe_prng_62_io_out_12),
    .io_out_13(rand_exe_prng_62_io_out_13),
    .io_out_14(rand_exe_prng_62_io_out_14),
    .io_out_15(rand_exe_prng_62_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_63 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_63_clock),
    .reset(rand_exe_prng_63_reset),
    .io_out_0(rand_exe_prng_63_io_out_0),
    .io_out_1(rand_exe_prng_63_io_out_1),
    .io_out_2(rand_exe_prng_63_io_out_2),
    .io_out_3(rand_exe_prng_63_io_out_3),
    .io_out_4(rand_exe_prng_63_io_out_4),
    .io_out_5(rand_exe_prng_63_io_out_5),
    .io_out_6(rand_exe_prng_63_io_out_6),
    .io_out_7(rand_exe_prng_63_io_out_7),
    .io_out_8(rand_exe_prng_63_io_out_8),
    .io_out_9(rand_exe_prng_63_io_out_9),
    .io_out_10(rand_exe_prng_63_io_out_10),
    .io_out_11(rand_exe_prng_63_io_out_11),
    .io_out_12(rand_exe_prng_63_io_out_12),
    .io_out_13(rand_exe_prng_63_io_out_13),
    .io_out_14(rand_exe_prng_63_io_out_14),
    .io_out_15(rand_exe_prng_63_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_64 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_64_clock),
    .reset(rand_exe_prng_64_reset),
    .io_out_0(rand_exe_prng_64_io_out_0),
    .io_out_1(rand_exe_prng_64_io_out_1),
    .io_out_2(rand_exe_prng_64_io_out_2),
    .io_out_3(rand_exe_prng_64_io_out_3),
    .io_out_4(rand_exe_prng_64_io_out_4),
    .io_out_5(rand_exe_prng_64_io_out_5),
    .io_out_6(rand_exe_prng_64_io_out_6),
    .io_out_7(rand_exe_prng_64_io_out_7),
    .io_out_8(rand_exe_prng_64_io_out_8),
    .io_out_9(rand_exe_prng_64_io_out_9),
    .io_out_10(rand_exe_prng_64_io_out_10),
    .io_out_11(rand_exe_prng_64_io_out_11),
    .io_out_12(rand_exe_prng_64_io_out_12),
    .io_out_13(rand_exe_prng_64_io_out_13),
    .io_out_14(rand_exe_prng_64_io_out_14),
    .io_out_15(rand_exe_prng_64_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_65 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_65_clock),
    .reset(rand_exe_prng_65_reset),
    .io_out_0(rand_exe_prng_65_io_out_0),
    .io_out_1(rand_exe_prng_65_io_out_1),
    .io_out_2(rand_exe_prng_65_io_out_2),
    .io_out_3(rand_exe_prng_65_io_out_3),
    .io_out_4(rand_exe_prng_65_io_out_4),
    .io_out_5(rand_exe_prng_65_io_out_5),
    .io_out_6(rand_exe_prng_65_io_out_6),
    .io_out_7(rand_exe_prng_65_io_out_7),
    .io_out_8(rand_exe_prng_65_io_out_8),
    .io_out_9(rand_exe_prng_65_io_out_9),
    .io_out_10(rand_exe_prng_65_io_out_10),
    .io_out_11(rand_exe_prng_65_io_out_11),
    .io_out_12(rand_exe_prng_65_io_out_12),
    .io_out_13(rand_exe_prng_65_io_out_13),
    .io_out_14(rand_exe_prng_65_io_out_14),
    .io_out_15(rand_exe_prng_65_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_66 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_66_clock),
    .reset(rand_exe_prng_66_reset),
    .io_out_0(rand_exe_prng_66_io_out_0),
    .io_out_1(rand_exe_prng_66_io_out_1),
    .io_out_2(rand_exe_prng_66_io_out_2),
    .io_out_3(rand_exe_prng_66_io_out_3),
    .io_out_4(rand_exe_prng_66_io_out_4),
    .io_out_5(rand_exe_prng_66_io_out_5),
    .io_out_6(rand_exe_prng_66_io_out_6),
    .io_out_7(rand_exe_prng_66_io_out_7),
    .io_out_8(rand_exe_prng_66_io_out_8),
    .io_out_9(rand_exe_prng_66_io_out_9),
    .io_out_10(rand_exe_prng_66_io_out_10),
    .io_out_11(rand_exe_prng_66_io_out_11),
    .io_out_12(rand_exe_prng_66_io_out_12),
    .io_out_13(rand_exe_prng_66_io_out_13),
    .io_out_14(rand_exe_prng_66_io_out_14),
    .io_out_15(rand_exe_prng_66_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_67 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_67_clock),
    .reset(rand_exe_prng_67_reset),
    .io_out_0(rand_exe_prng_67_io_out_0),
    .io_out_1(rand_exe_prng_67_io_out_1),
    .io_out_2(rand_exe_prng_67_io_out_2),
    .io_out_3(rand_exe_prng_67_io_out_3),
    .io_out_4(rand_exe_prng_67_io_out_4),
    .io_out_5(rand_exe_prng_67_io_out_5),
    .io_out_6(rand_exe_prng_67_io_out_6),
    .io_out_7(rand_exe_prng_67_io_out_7),
    .io_out_8(rand_exe_prng_67_io_out_8),
    .io_out_9(rand_exe_prng_67_io_out_9),
    .io_out_10(rand_exe_prng_67_io_out_10),
    .io_out_11(rand_exe_prng_67_io_out_11),
    .io_out_12(rand_exe_prng_67_io_out_12),
    .io_out_13(rand_exe_prng_67_io_out_13),
    .io_out_14(rand_exe_prng_67_io_out_14),
    .io_out_15(rand_exe_prng_67_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_68 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_68_clock),
    .reset(rand_exe_prng_68_reset),
    .io_out_0(rand_exe_prng_68_io_out_0),
    .io_out_1(rand_exe_prng_68_io_out_1),
    .io_out_2(rand_exe_prng_68_io_out_2),
    .io_out_3(rand_exe_prng_68_io_out_3),
    .io_out_4(rand_exe_prng_68_io_out_4),
    .io_out_5(rand_exe_prng_68_io_out_5),
    .io_out_6(rand_exe_prng_68_io_out_6),
    .io_out_7(rand_exe_prng_68_io_out_7),
    .io_out_8(rand_exe_prng_68_io_out_8),
    .io_out_9(rand_exe_prng_68_io_out_9),
    .io_out_10(rand_exe_prng_68_io_out_10),
    .io_out_11(rand_exe_prng_68_io_out_11),
    .io_out_12(rand_exe_prng_68_io_out_12),
    .io_out_13(rand_exe_prng_68_io_out_13),
    .io_out_14(rand_exe_prng_68_io_out_14),
    .io_out_15(rand_exe_prng_68_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_69 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_69_clock),
    .reset(rand_exe_prng_69_reset),
    .io_out_0(rand_exe_prng_69_io_out_0),
    .io_out_1(rand_exe_prng_69_io_out_1),
    .io_out_2(rand_exe_prng_69_io_out_2),
    .io_out_3(rand_exe_prng_69_io_out_3),
    .io_out_4(rand_exe_prng_69_io_out_4),
    .io_out_5(rand_exe_prng_69_io_out_5),
    .io_out_6(rand_exe_prng_69_io_out_6),
    .io_out_7(rand_exe_prng_69_io_out_7),
    .io_out_8(rand_exe_prng_69_io_out_8),
    .io_out_9(rand_exe_prng_69_io_out_9),
    .io_out_10(rand_exe_prng_69_io_out_10),
    .io_out_11(rand_exe_prng_69_io_out_11),
    .io_out_12(rand_exe_prng_69_io_out_12),
    .io_out_13(rand_exe_prng_69_io_out_13),
    .io_out_14(rand_exe_prng_69_io_out_14),
    .io_out_15(rand_exe_prng_69_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_70 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_70_clock),
    .reset(rand_exe_prng_70_reset),
    .io_out_0(rand_exe_prng_70_io_out_0),
    .io_out_1(rand_exe_prng_70_io_out_1),
    .io_out_2(rand_exe_prng_70_io_out_2),
    .io_out_3(rand_exe_prng_70_io_out_3),
    .io_out_4(rand_exe_prng_70_io_out_4),
    .io_out_5(rand_exe_prng_70_io_out_5),
    .io_out_6(rand_exe_prng_70_io_out_6),
    .io_out_7(rand_exe_prng_70_io_out_7),
    .io_out_8(rand_exe_prng_70_io_out_8),
    .io_out_9(rand_exe_prng_70_io_out_9),
    .io_out_10(rand_exe_prng_70_io_out_10),
    .io_out_11(rand_exe_prng_70_io_out_11),
    .io_out_12(rand_exe_prng_70_io_out_12),
    .io_out_13(rand_exe_prng_70_io_out_13),
    .io_out_14(rand_exe_prng_70_io_out_14),
    .io_out_15(rand_exe_prng_70_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_71 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_71_clock),
    .reset(rand_exe_prng_71_reset),
    .io_out_0(rand_exe_prng_71_io_out_0),
    .io_out_1(rand_exe_prng_71_io_out_1),
    .io_out_2(rand_exe_prng_71_io_out_2),
    .io_out_3(rand_exe_prng_71_io_out_3),
    .io_out_4(rand_exe_prng_71_io_out_4),
    .io_out_5(rand_exe_prng_71_io_out_5),
    .io_out_6(rand_exe_prng_71_io_out_6),
    .io_out_7(rand_exe_prng_71_io_out_7),
    .io_out_8(rand_exe_prng_71_io_out_8),
    .io_out_9(rand_exe_prng_71_io_out_9),
    .io_out_10(rand_exe_prng_71_io_out_10),
    .io_out_11(rand_exe_prng_71_io_out_11),
    .io_out_12(rand_exe_prng_71_io_out_12),
    .io_out_13(rand_exe_prng_71_io_out_13),
    .io_out_14(rand_exe_prng_71_io_out_14),
    .io_out_15(rand_exe_prng_71_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_72 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_72_clock),
    .reset(rand_exe_prng_72_reset),
    .io_out_0(rand_exe_prng_72_io_out_0),
    .io_out_1(rand_exe_prng_72_io_out_1),
    .io_out_2(rand_exe_prng_72_io_out_2),
    .io_out_3(rand_exe_prng_72_io_out_3),
    .io_out_4(rand_exe_prng_72_io_out_4),
    .io_out_5(rand_exe_prng_72_io_out_5),
    .io_out_6(rand_exe_prng_72_io_out_6),
    .io_out_7(rand_exe_prng_72_io_out_7),
    .io_out_8(rand_exe_prng_72_io_out_8),
    .io_out_9(rand_exe_prng_72_io_out_9),
    .io_out_10(rand_exe_prng_72_io_out_10),
    .io_out_11(rand_exe_prng_72_io_out_11),
    .io_out_12(rand_exe_prng_72_io_out_12),
    .io_out_13(rand_exe_prng_72_io_out_13),
    .io_out_14(rand_exe_prng_72_io_out_14),
    .io_out_15(rand_exe_prng_72_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_73 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_73_clock),
    .reset(rand_exe_prng_73_reset),
    .io_out_0(rand_exe_prng_73_io_out_0),
    .io_out_1(rand_exe_prng_73_io_out_1),
    .io_out_2(rand_exe_prng_73_io_out_2),
    .io_out_3(rand_exe_prng_73_io_out_3),
    .io_out_4(rand_exe_prng_73_io_out_4),
    .io_out_5(rand_exe_prng_73_io_out_5),
    .io_out_6(rand_exe_prng_73_io_out_6),
    .io_out_7(rand_exe_prng_73_io_out_7),
    .io_out_8(rand_exe_prng_73_io_out_8),
    .io_out_9(rand_exe_prng_73_io_out_9),
    .io_out_10(rand_exe_prng_73_io_out_10),
    .io_out_11(rand_exe_prng_73_io_out_11),
    .io_out_12(rand_exe_prng_73_io_out_12),
    .io_out_13(rand_exe_prng_73_io_out_13),
    .io_out_14(rand_exe_prng_73_io_out_14),
    .io_out_15(rand_exe_prng_73_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_74 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_74_clock),
    .reset(rand_exe_prng_74_reset),
    .io_out_0(rand_exe_prng_74_io_out_0),
    .io_out_1(rand_exe_prng_74_io_out_1),
    .io_out_2(rand_exe_prng_74_io_out_2),
    .io_out_3(rand_exe_prng_74_io_out_3),
    .io_out_4(rand_exe_prng_74_io_out_4),
    .io_out_5(rand_exe_prng_74_io_out_5),
    .io_out_6(rand_exe_prng_74_io_out_6),
    .io_out_7(rand_exe_prng_74_io_out_7),
    .io_out_8(rand_exe_prng_74_io_out_8),
    .io_out_9(rand_exe_prng_74_io_out_9),
    .io_out_10(rand_exe_prng_74_io_out_10),
    .io_out_11(rand_exe_prng_74_io_out_11),
    .io_out_12(rand_exe_prng_74_io_out_12),
    .io_out_13(rand_exe_prng_74_io_out_13),
    .io_out_14(rand_exe_prng_74_io_out_14),
    .io_out_15(rand_exe_prng_74_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_75 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_75_clock),
    .reset(rand_exe_prng_75_reset),
    .io_out_0(rand_exe_prng_75_io_out_0),
    .io_out_1(rand_exe_prng_75_io_out_1),
    .io_out_2(rand_exe_prng_75_io_out_2),
    .io_out_3(rand_exe_prng_75_io_out_3),
    .io_out_4(rand_exe_prng_75_io_out_4),
    .io_out_5(rand_exe_prng_75_io_out_5),
    .io_out_6(rand_exe_prng_75_io_out_6),
    .io_out_7(rand_exe_prng_75_io_out_7),
    .io_out_8(rand_exe_prng_75_io_out_8),
    .io_out_9(rand_exe_prng_75_io_out_9),
    .io_out_10(rand_exe_prng_75_io_out_10),
    .io_out_11(rand_exe_prng_75_io_out_11),
    .io_out_12(rand_exe_prng_75_io_out_12),
    .io_out_13(rand_exe_prng_75_io_out_13),
    .io_out_14(rand_exe_prng_75_io_out_14),
    .io_out_15(rand_exe_prng_75_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_76 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_76_clock),
    .reset(rand_exe_prng_76_reset),
    .io_out_0(rand_exe_prng_76_io_out_0),
    .io_out_1(rand_exe_prng_76_io_out_1),
    .io_out_2(rand_exe_prng_76_io_out_2),
    .io_out_3(rand_exe_prng_76_io_out_3),
    .io_out_4(rand_exe_prng_76_io_out_4),
    .io_out_5(rand_exe_prng_76_io_out_5),
    .io_out_6(rand_exe_prng_76_io_out_6),
    .io_out_7(rand_exe_prng_76_io_out_7),
    .io_out_8(rand_exe_prng_76_io_out_8),
    .io_out_9(rand_exe_prng_76_io_out_9),
    .io_out_10(rand_exe_prng_76_io_out_10),
    .io_out_11(rand_exe_prng_76_io_out_11),
    .io_out_12(rand_exe_prng_76_io_out_12),
    .io_out_13(rand_exe_prng_76_io_out_13),
    .io_out_14(rand_exe_prng_76_io_out_14),
    .io_out_15(rand_exe_prng_76_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_77 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_77_clock),
    .reset(rand_exe_prng_77_reset),
    .io_out_0(rand_exe_prng_77_io_out_0),
    .io_out_1(rand_exe_prng_77_io_out_1),
    .io_out_2(rand_exe_prng_77_io_out_2),
    .io_out_3(rand_exe_prng_77_io_out_3),
    .io_out_4(rand_exe_prng_77_io_out_4),
    .io_out_5(rand_exe_prng_77_io_out_5),
    .io_out_6(rand_exe_prng_77_io_out_6),
    .io_out_7(rand_exe_prng_77_io_out_7),
    .io_out_8(rand_exe_prng_77_io_out_8),
    .io_out_9(rand_exe_prng_77_io_out_9),
    .io_out_10(rand_exe_prng_77_io_out_10),
    .io_out_11(rand_exe_prng_77_io_out_11),
    .io_out_12(rand_exe_prng_77_io_out_12),
    .io_out_13(rand_exe_prng_77_io_out_13),
    .io_out_14(rand_exe_prng_77_io_out_14),
    .io_out_15(rand_exe_prng_77_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_78 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_78_clock),
    .reset(rand_exe_prng_78_reset),
    .io_out_0(rand_exe_prng_78_io_out_0),
    .io_out_1(rand_exe_prng_78_io_out_1),
    .io_out_2(rand_exe_prng_78_io_out_2),
    .io_out_3(rand_exe_prng_78_io_out_3),
    .io_out_4(rand_exe_prng_78_io_out_4),
    .io_out_5(rand_exe_prng_78_io_out_5),
    .io_out_6(rand_exe_prng_78_io_out_6),
    .io_out_7(rand_exe_prng_78_io_out_7),
    .io_out_8(rand_exe_prng_78_io_out_8),
    .io_out_9(rand_exe_prng_78_io_out_9),
    .io_out_10(rand_exe_prng_78_io_out_10),
    .io_out_11(rand_exe_prng_78_io_out_11),
    .io_out_12(rand_exe_prng_78_io_out_12),
    .io_out_13(rand_exe_prng_78_io_out_13),
    .io_out_14(rand_exe_prng_78_io_out_14),
    .io_out_15(rand_exe_prng_78_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_79 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_79_clock),
    .reset(rand_exe_prng_79_reset),
    .io_out_0(rand_exe_prng_79_io_out_0),
    .io_out_1(rand_exe_prng_79_io_out_1),
    .io_out_2(rand_exe_prng_79_io_out_2),
    .io_out_3(rand_exe_prng_79_io_out_3),
    .io_out_4(rand_exe_prng_79_io_out_4),
    .io_out_5(rand_exe_prng_79_io_out_5),
    .io_out_6(rand_exe_prng_79_io_out_6),
    .io_out_7(rand_exe_prng_79_io_out_7),
    .io_out_8(rand_exe_prng_79_io_out_8),
    .io_out_9(rand_exe_prng_79_io_out_9),
    .io_out_10(rand_exe_prng_79_io_out_10),
    .io_out_11(rand_exe_prng_79_io_out_11),
    .io_out_12(rand_exe_prng_79_io_out_12),
    .io_out_13(rand_exe_prng_79_io_out_13),
    .io_out_14(rand_exe_prng_79_io_out_14),
    .io_out_15(rand_exe_prng_79_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_80 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_80_clock),
    .reset(rand_exe_prng_80_reset),
    .io_out_0(rand_exe_prng_80_io_out_0),
    .io_out_1(rand_exe_prng_80_io_out_1),
    .io_out_2(rand_exe_prng_80_io_out_2),
    .io_out_3(rand_exe_prng_80_io_out_3),
    .io_out_4(rand_exe_prng_80_io_out_4),
    .io_out_5(rand_exe_prng_80_io_out_5),
    .io_out_6(rand_exe_prng_80_io_out_6),
    .io_out_7(rand_exe_prng_80_io_out_7),
    .io_out_8(rand_exe_prng_80_io_out_8),
    .io_out_9(rand_exe_prng_80_io_out_9),
    .io_out_10(rand_exe_prng_80_io_out_10),
    .io_out_11(rand_exe_prng_80_io_out_11),
    .io_out_12(rand_exe_prng_80_io_out_12),
    .io_out_13(rand_exe_prng_80_io_out_13),
    .io_out_14(rand_exe_prng_80_io_out_14),
    .io_out_15(rand_exe_prng_80_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_81 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_81_clock),
    .reset(rand_exe_prng_81_reset),
    .io_out_0(rand_exe_prng_81_io_out_0),
    .io_out_1(rand_exe_prng_81_io_out_1),
    .io_out_2(rand_exe_prng_81_io_out_2),
    .io_out_3(rand_exe_prng_81_io_out_3),
    .io_out_4(rand_exe_prng_81_io_out_4),
    .io_out_5(rand_exe_prng_81_io_out_5),
    .io_out_6(rand_exe_prng_81_io_out_6),
    .io_out_7(rand_exe_prng_81_io_out_7),
    .io_out_8(rand_exe_prng_81_io_out_8),
    .io_out_9(rand_exe_prng_81_io_out_9),
    .io_out_10(rand_exe_prng_81_io_out_10),
    .io_out_11(rand_exe_prng_81_io_out_11),
    .io_out_12(rand_exe_prng_81_io_out_12),
    .io_out_13(rand_exe_prng_81_io_out_13),
    .io_out_14(rand_exe_prng_81_io_out_14),
    .io_out_15(rand_exe_prng_81_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_82 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_82_clock),
    .reset(rand_exe_prng_82_reset),
    .io_out_0(rand_exe_prng_82_io_out_0),
    .io_out_1(rand_exe_prng_82_io_out_1),
    .io_out_2(rand_exe_prng_82_io_out_2),
    .io_out_3(rand_exe_prng_82_io_out_3),
    .io_out_4(rand_exe_prng_82_io_out_4),
    .io_out_5(rand_exe_prng_82_io_out_5),
    .io_out_6(rand_exe_prng_82_io_out_6),
    .io_out_7(rand_exe_prng_82_io_out_7),
    .io_out_8(rand_exe_prng_82_io_out_8),
    .io_out_9(rand_exe_prng_82_io_out_9),
    .io_out_10(rand_exe_prng_82_io_out_10),
    .io_out_11(rand_exe_prng_82_io_out_11),
    .io_out_12(rand_exe_prng_82_io_out_12),
    .io_out_13(rand_exe_prng_82_io_out_13),
    .io_out_14(rand_exe_prng_82_io_out_14),
    .io_out_15(rand_exe_prng_82_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_83 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_83_clock),
    .reset(rand_exe_prng_83_reset),
    .io_out_0(rand_exe_prng_83_io_out_0),
    .io_out_1(rand_exe_prng_83_io_out_1),
    .io_out_2(rand_exe_prng_83_io_out_2),
    .io_out_3(rand_exe_prng_83_io_out_3),
    .io_out_4(rand_exe_prng_83_io_out_4),
    .io_out_5(rand_exe_prng_83_io_out_5),
    .io_out_6(rand_exe_prng_83_io_out_6),
    .io_out_7(rand_exe_prng_83_io_out_7),
    .io_out_8(rand_exe_prng_83_io_out_8),
    .io_out_9(rand_exe_prng_83_io_out_9),
    .io_out_10(rand_exe_prng_83_io_out_10),
    .io_out_11(rand_exe_prng_83_io_out_11),
    .io_out_12(rand_exe_prng_83_io_out_12),
    .io_out_13(rand_exe_prng_83_io_out_13),
    .io_out_14(rand_exe_prng_83_io_out_14),
    .io_out_15(rand_exe_prng_83_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_84 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_84_clock),
    .reset(rand_exe_prng_84_reset),
    .io_out_0(rand_exe_prng_84_io_out_0),
    .io_out_1(rand_exe_prng_84_io_out_1),
    .io_out_2(rand_exe_prng_84_io_out_2),
    .io_out_3(rand_exe_prng_84_io_out_3),
    .io_out_4(rand_exe_prng_84_io_out_4),
    .io_out_5(rand_exe_prng_84_io_out_5),
    .io_out_6(rand_exe_prng_84_io_out_6),
    .io_out_7(rand_exe_prng_84_io_out_7),
    .io_out_8(rand_exe_prng_84_io_out_8),
    .io_out_9(rand_exe_prng_84_io_out_9),
    .io_out_10(rand_exe_prng_84_io_out_10),
    .io_out_11(rand_exe_prng_84_io_out_11),
    .io_out_12(rand_exe_prng_84_io_out_12),
    .io_out_13(rand_exe_prng_84_io_out_13),
    .io_out_14(rand_exe_prng_84_io_out_14),
    .io_out_15(rand_exe_prng_84_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_85 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_85_clock),
    .reset(rand_exe_prng_85_reset),
    .io_out_0(rand_exe_prng_85_io_out_0),
    .io_out_1(rand_exe_prng_85_io_out_1),
    .io_out_2(rand_exe_prng_85_io_out_2),
    .io_out_3(rand_exe_prng_85_io_out_3),
    .io_out_4(rand_exe_prng_85_io_out_4),
    .io_out_5(rand_exe_prng_85_io_out_5),
    .io_out_6(rand_exe_prng_85_io_out_6),
    .io_out_7(rand_exe_prng_85_io_out_7),
    .io_out_8(rand_exe_prng_85_io_out_8),
    .io_out_9(rand_exe_prng_85_io_out_9),
    .io_out_10(rand_exe_prng_85_io_out_10),
    .io_out_11(rand_exe_prng_85_io_out_11),
    .io_out_12(rand_exe_prng_85_io_out_12),
    .io_out_13(rand_exe_prng_85_io_out_13),
    .io_out_14(rand_exe_prng_85_io_out_14),
    .io_out_15(rand_exe_prng_85_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_86 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_86_clock),
    .reset(rand_exe_prng_86_reset),
    .io_out_0(rand_exe_prng_86_io_out_0),
    .io_out_1(rand_exe_prng_86_io_out_1),
    .io_out_2(rand_exe_prng_86_io_out_2),
    .io_out_3(rand_exe_prng_86_io_out_3),
    .io_out_4(rand_exe_prng_86_io_out_4),
    .io_out_5(rand_exe_prng_86_io_out_5),
    .io_out_6(rand_exe_prng_86_io_out_6),
    .io_out_7(rand_exe_prng_86_io_out_7),
    .io_out_8(rand_exe_prng_86_io_out_8),
    .io_out_9(rand_exe_prng_86_io_out_9),
    .io_out_10(rand_exe_prng_86_io_out_10),
    .io_out_11(rand_exe_prng_86_io_out_11),
    .io_out_12(rand_exe_prng_86_io_out_12),
    .io_out_13(rand_exe_prng_86_io_out_13),
    .io_out_14(rand_exe_prng_86_io_out_14),
    .io_out_15(rand_exe_prng_86_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_87 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_87_clock),
    .reset(rand_exe_prng_87_reset),
    .io_out_0(rand_exe_prng_87_io_out_0),
    .io_out_1(rand_exe_prng_87_io_out_1),
    .io_out_2(rand_exe_prng_87_io_out_2),
    .io_out_3(rand_exe_prng_87_io_out_3),
    .io_out_4(rand_exe_prng_87_io_out_4),
    .io_out_5(rand_exe_prng_87_io_out_5),
    .io_out_6(rand_exe_prng_87_io_out_6),
    .io_out_7(rand_exe_prng_87_io_out_7),
    .io_out_8(rand_exe_prng_87_io_out_8),
    .io_out_9(rand_exe_prng_87_io_out_9),
    .io_out_10(rand_exe_prng_87_io_out_10),
    .io_out_11(rand_exe_prng_87_io_out_11),
    .io_out_12(rand_exe_prng_87_io_out_12),
    .io_out_13(rand_exe_prng_87_io_out_13),
    .io_out_14(rand_exe_prng_87_io_out_14),
    .io_out_15(rand_exe_prng_87_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_88 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_88_clock),
    .reset(rand_exe_prng_88_reset),
    .io_out_0(rand_exe_prng_88_io_out_0),
    .io_out_1(rand_exe_prng_88_io_out_1),
    .io_out_2(rand_exe_prng_88_io_out_2),
    .io_out_3(rand_exe_prng_88_io_out_3),
    .io_out_4(rand_exe_prng_88_io_out_4),
    .io_out_5(rand_exe_prng_88_io_out_5),
    .io_out_6(rand_exe_prng_88_io_out_6),
    .io_out_7(rand_exe_prng_88_io_out_7),
    .io_out_8(rand_exe_prng_88_io_out_8),
    .io_out_9(rand_exe_prng_88_io_out_9),
    .io_out_10(rand_exe_prng_88_io_out_10),
    .io_out_11(rand_exe_prng_88_io_out_11),
    .io_out_12(rand_exe_prng_88_io_out_12),
    .io_out_13(rand_exe_prng_88_io_out_13),
    .io_out_14(rand_exe_prng_88_io_out_14),
    .io_out_15(rand_exe_prng_88_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_89 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_89_clock),
    .reset(rand_exe_prng_89_reset),
    .io_out_0(rand_exe_prng_89_io_out_0),
    .io_out_1(rand_exe_prng_89_io_out_1),
    .io_out_2(rand_exe_prng_89_io_out_2),
    .io_out_3(rand_exe_prng_89_io_out_3),
    .io_out_4(rand_exe_prng_89_io_out_4),
    .io_out_5(rand_exe_prng_89_io_out_5),
    .io_out_6(rand_exe_prng_89_io_out_6),
    .io_out_7(rand_exe_prng_89_io_out_7),
    .io_out_8(rand_exe_prng_89_io_out_8),
    .io_out_9(rand_exe_prng_89_io_out_9),
    .io_out_10(rand_exe_prng_89_io_out_10),
    .io_out_11(rand_exe_prng_89_io_out_11),
    .io_out_12(rand_exe_prng_89_io_out_12),
    .io_out_13(rand_exe_prng_89_io_out_13),
    .io_out_14(rand_exe_prng_89_io_out_14),
    .io_out_15(rand_exe_prng_89_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_90 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_90_clock),
    .reset(rand_exe_prng_90_reset),
    .io_out_0(rand_exe_prng_90_io_out_0),
    .io_out_1(rand_exe_prng_90_io_out_1),
    .io_out_2(rand_exe_prng_90_io_out_2),
    .io_out_3(rand_exe_prng_90_io_out_3),
    .io_out_4(rand_exe_prng_90_io_out_4),
    .io_out_5(rand_exe_prng_90_io_out_5),
    .io_out_6(rand_exe_prng_90_io_out_6),
    .io_out_7(rand_exe_prng_90_io_out_7),
    .io_out_8(rand_exe_prng_90_io_out_8),
    .io_out_9(rand_exe_prng_90_io_out_9),
    .io_out_10(rand_exe_prng_90_io_out_10),
    .io_out_11(rand_exe_prng_90_io_out_11),
    .io_out_12(rand_exe_prng_90_io_out_12),
    .io_out_13(rand_exe_prng_90_io_out_13),
    .io_out_14(rand_exe_prng_90_io_out_14),
    .io_out_15(rand_exe_prng_90_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_91 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_91_clock),
    .reset(rand_exe_prng_91_reset),
    .io_out_0(rand_exe_prng_91_io_out_0),
    .io_out_1(rand_exe_prng_91_io_out_1),
    .io_out_2(rand_exe_prng_91_io_out_2),
    .io_out_3(rand_exe_prng_91_io_out_3),
    .io_out_4(rand_exe_prng_91_io_out_4),
    .io_out_5(rand_exe_prng_91_io_out_5),
    .io_out_6(rand_exe_prng_91_io_out_6),
    .io_out_7(rand_exe_prng_91_io_out_7),
    .io_out_8(rand_exe_prng_91_io_out_8),
    .io_out_9(rand_exe_prng_91_io_out_9),
    .io_out_10(rand_exe_prng_91_io_out_10),
    .io_out_11(rand_exe_prng_91_io_out_11),
    .io_out_12(rand_exe_prng_91_io_out_12),
    .io_out_13(rand_exe_prng_91_io_out_13),
    .io_out_14(rand_exe_prng_91_io_out_14),
    .io_out_15(rand_exe_prng_91_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_92 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_92_clock),
    .reset(rand_exe_prng_92_reset),
    .io_out_0(rand_exe_prng_92_io_out_0),
    .io_out_1(rand_exe_prng_92_io_out_1),
    .io_out_2(rand_exe_prng_92_io_out_2),
    .io_out_3(rand_exe_prng_92_io_out_3),
    .io_out_4(rand_exe_prng_92_io_out_4),
    .io_out_5(rand_exe_prng_92_io_out_5),
    .io_out_6(rand_exe_prng_92_io_out_6),
    .io_out_7(rand_exe_prng_92_io_out_7),
    .io_out_8(rand_exe_prng_92_io_out_8),
    .io_out_9(rand_exe_prng_92_io_out_9),
    .io_out_10(rand_exe_prng_92_io_out_10),
    .io_out_11(rand_exe_prng_92_io_out_11),
    .io_out_12(rand_exe_prng_92_io_out_12),
    .io_out_13(rand_exe_prng_92_io_out_13),
    .io_out_14(rand_exe_prng_92_io_out_14),
    .io_out_15(rand_exe_prng_92_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_93 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_93_clock),
    .reset(rand_exe_prng_93_reset),
    .io_out_0(rand_exe_prng_93_io_out_0),
    .io_out_1(rand_exe_prng_93_io_out_1),
    .io_out_2(rand_exe_prng_93_io_out_2),
    .io_out_3(rand_exe_prng_93_io_out_3),
    .io_out_4(rand_exe_prng_93_io_out_4),
    .io_out_5(rand_exe_prng_93_io_out_5),
    .io_out_6(rand_exe_prng_93_io_out_6),
    .io_out_7(rand_exe_prng_93_io_out_7),
    .io_out_8(rand_exe_prng_93_io_out_8),
    .io_out_9(rand_exe_prng_93_io_out_9),
    .io_out_10(rand_exe_prng_93_io_out_10),
    .io_out_11(rand_exe_prng_93_io_out_11),
    .io_out_12(rand_exe_prng_93_io_out_12),
    .io_out_13(rand_exe_prng_93_io_out_13),
    .io_out_14(rand_exe_prng_93_io_out_14),
    .io_out_15(rand_exe_prng_93_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_94 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_94_clock),
    .reset(rand_exe_prng_94_reset),
    .io_out_0(rand_exe_prng_94_io_out_0),
    .io_out_1(rand_exe_prng_94_io_out_1),
    .io_out_2(rand_exe_prng_94_io_out_2),
    .io_out_3(rand_exe_prng_94_io_out_3),
    .io_out_4(rand_exe_prng_94_io_out_4),
    .io_out_5(rand_exe_prng_94_io_out_5),
    .io_out_6(rand_exe_prng_94_io_out_6),
    .io_out_7(rand_exe_prng_94_io_out_7),
    .io_out_8(rand_exe_prng_94_io_out_8),
    .io_out_9(rand_exe_prng_94_io_out_9),
    .io_out_10(rand_exe_prng_94_io_out_10),
    .io_out_11(rand_exe_prng_94_io_out_11),
    .io_out_12(rand_exe_prng_94_io_out_12),
    .io_out_13(rand_exe_prng_94_io_out_13),
    .io_out_14(rand_exe_prng_94_io_out_14),
    .io_out_15(rand_exe_prng_94_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_95 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_95_clock),
    .reset(rand_exe_prng_95_reset),
    .io_out_0(rand_exe_prng_95_io_out_0),
    .io_out_1(rand_exe_prng_95_io_out_1),
    .io_out_2(rand_exe_prng_95_io_out_2),
    .io_out_3(rand_exe_prng_95_io_out_3),
    .io_out_4(rand_exe_prng_95_io_out_4),
    .io_out_5(rand_exe_prng_95_io_out_5),
    .io_out_6(rand_exe_prng_95_io_out_6),
    .io_out_7(rand_exe_prng_95_io_out_7),
    .io_out_8(rand_exe_prng_95_io_out_8),
    .io_out_9(rand_exe_prng_95_io_out_9),
    .io_out_10(rand_exe_prng_95_io_out_10),
    .io_out_11(rand_exe_prng_95_io_out_11),
    .io_out_12(rand_exe_prng_95_io_out_12),
    .io_out_13(rand_exe_prng_95_io_out_13),
    .io_out_14(rand_exe_prng_95_io_out_14),
    .io_out_15(rand_exe_prng_95_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_96 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_96_clock),
    .reset(rand_exe_prng_96_reset),
    .io_out_0(rand_exe_prng_96_io_out_0),
    .io_out_1(rand_exe_prng_96_io_out_1),
    .io_out_2(rand_exe_prng_96_io_out_2),
    .io_out_3(rand_exe_prng_96_io_out_3),
    .io_out_4(rand_exe_prng_96_io_out_4),
    .io_out_5(rand_exe_prng_96_io_out_5),
    .io_out_6(rand_exe_prng_96_io_out_6),
    .io_out_7(rand_exe_prng_96_io_out_7),
    .io_out_8(rand_exe_prng_96_io_out_8),
    .io_out_9(rand_exe_prng_96_io_out_9),
    .io_out_10(rand_exe_prng_96_io_out_10),
    .io_out_11(rand_exe_prng_96_io_out_11),
    .io_out_12(rand_exe_prng_96_io_out_12),
    .io_out_13(rand_exe_prng_96_io_out_13),
    .io_out_14(rand_exe_prng_96_io_out_14),
    .io_out_15(rand_exe_prng_96_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_97 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_97_clock),
    .reset(rand_exe_prng_97_reset),
    .io_out_0(rand_exe_prng_97_io_out_0),
    .io_out_1(rand_exe_prng_97_io_out_1),
    .io_out_2(rand_exe_prng_97_io_out_2),
    .io_out_3(rand_exe_prng_97_io_out_3),
    .io_out_4(rand_exe_prng_97_io_out_4),
    .io_out_5(rand_exe_prng_97_io_out_5),
    .io_out_6(rand_exe_prng_97_io_out_6),
    .io_out_7(rand_exe_prng_97_io_out_7),
    .io_out_8(rand_exe_prng_97_io_out_8),
    .io_out_9(rand_exe_prng_97_io_out_9),
    .io_out_10(rand_exe_prng_97_io_out_10),
    .io_out_11(rand_exe_prng_97_io_out_11),
    .io_out_12(rand_exe_prng_97_io_out_12),
    .io_out_13(rand_exe_prng_97_io_out_13),
    .io_out_14(rand_exe_prng_97_io_out_14),
    .io_out_15(rand_exe_prng_97_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_98 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_98_clock),
    .reset(rand_exe_prng_98_reset),
    .io_out_0(rand_exe_prng_98_io_out_0),
    .io_out_1(rand_exe_prng_98_io_out_1),
    .io_out_2(rand_exe_prng_98_io_out_2),
    .io_out_3(rand_exe_prng_98_io_out_3),
    .io_out_4(rand_exe_prng_98_io_out_4),
    .io_out_5(rand_exe_prng_98_io_out_5),
    .io_out_6(rand_exe_prng_98_io_out_6),
    .io_out_7(rand_exe_prng_98_io_out_7),
    .io_out_8(rand_exe_prng_98_io_out_8),
    .io_out_9(rand_exe_prng_98_io_out_9),
    .io_out_10(rand_exe_prng_98_io_out_10),
    .io_out_11(rand_exe_prng_98_io_out_11),
    .io_out_12(rand_exe_prng_98_io_out_12),
    .io_out_13(rand_exe_prng_98_io_out_13),
    .io_out_14(rand_exe_prng_98_io_out_14),
    .io_out_15(rand_exe_prng_98_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_99 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_99_clock),
    .reset(rand_exe_prng_99_reset),
    .io_out_0(rand_exe_prng_99_io_out_0),
    .io_out_1(rand_exe_prng_99_io_out_1),
    .io_out_2(rand_exe_prng_99_io_out_2),
    .io_out_3(rand_exe_prng_99_io_out_3),
    .io_out_4(rand_exe_prng_99_io_out_4),
    .io_out_5(rand_exe_prng_99_io_out_5),
    .io_out_6(rand_exe_prng_99_io_out_6),
    .io_out_7(rand_exe_prng_99_io_out_7),
    .io_out_8(rand_exe_prng_99_io_out_8),
    .io_out_9(rand_exe_prng_99_io_out_9),
    .io_out_10(rand_exe_prng_99_io_out_10),
    .io_out_11(rand_exe_prng_99_io_out_11),
    .io_out_12(rand_exe_prng_99_io_out_12),
    .io_out_13(rand_exe_prng_99_io_out_13),
    .io_out_14(rand_exe_prng_99_io_out_14),
    .io_out_15(rand_exe_prng_99_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_100 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_100_clock),
    .reset(rand_exe_prng_100_reset),
    .io_out_0(rand_exe_prng_100_io_out_0),
    .io_out_1(rand_exe_prng_100_io_out_1),
    .io_out_2(rand_exe_prng_100_io_out_2),
    .io_out_3(rand_exe_prng_100_io_out_3),
    .io_out_4(rand_exe_prng_100_io_out_4),
    .io_out_5(rand_exe_prng_100_io_out_5),
    .io_out_6(rand_exe_prng_100_io_out_6),
    .io_out_7(rand_exe_prng_100_io_out_7),
    .io_out_8(rand_exe_prng_100_io_out_8),
    .io_out_9(rand_exe_prng_100_io_out_9),
    .io_out_10(rand_exe_prng_100_io_out_10),
    .io_out_11(rand_exe_prng_100_io_out_11),
    .io_out_12(rand_exe_prng_100_io_out_12),
    .io_out_13(rand_exe_prng_100_io_out_13),
    .io_out_14(rand_exe_prng_100_io_out_14),
    .io_out_15(rand_exe_prng_100_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_101 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_101_clock),
    .reset(rand_exe_prng_101_reset),
    .io_out_0(rand_exe_prng_101_io_out_0),
    .io_out_1(rand_exe_prng_101_io_out_1),
    .io_out_2(rand_exe_prng_101_io_out_2),
    .io_out_3(rand_exe_prng_101_io_out_3),
    .io_out_4(rand_exe_prng_101_io_out_4),
    .io_out_5(rand_exe_prng_101_io_out_5),
    .io_out_6(rand_exe_prng_101_io_out_6),
    .io_out_7(rand_exe_prng_101_io_out_7),
    .io_out_8(rand_exe_prng_101_io_out_8),
    .io_out_9(rand_exe_prng_101_io_out_9),
    .io_out_10(rand_exe_prng_101_io_out_10),
    .io_out_11(rand_exe_prng_101_io_out_11),
    .io_out_12(rand_exe_prng_101_io_out_12),
    .io_out_13(rand_exe_prng_101_io_out_13),
    .io_out_14(rand_exe_prng_101_io_out_14),
    .io_out_15(rand_exe_prng_101_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_102 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_102_clock),
    .reset(rand_exe_prng_102_reset),
    .io_out_0(rand_exe_prng_102_io_out_0),
    .io_out_1(rand_exe_prng_102_io_out_1),
    .io_out_2(rand_exe_prng_102_io_out_2),
    .io_out_3(rand_exe_prng_102_io_out_3),
    .io_out_4(rand_exe_prng_102_io_out_4),
    .io_out_5(rand_exe_prng_102_io_out_5),
    .io_out_6(rand_exe_prng_102_io_out_6),
    .io_out_7(rand_exe_prng_102_io_out_7),
    .io_out_8(rand_exe_prng_102_io_out_8),
    .io_out_9(rand_exe_prng_102_io_out_9),
    .io_out_10(rand_exe_prng_102_io_out_10),
    .io_out_11(rand_exe_prng_102_io_out_11),
    .io_out_12(rand_exe_prng_102_io_out_12),
    .io_out_13(rand_exe_prng_102_io_out_13),
    .io_out_14(rand_exe_prng_102_io_out_14),
    .io_out_15(rand_exe_prng_102_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_103 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_103_clock),
    .reset(rand_exe_prng_103_reset),
    .io_out_0(rand_exe_prng_103_io_out_0),
    .io_out_1(rand_exe_prng_103_io_out_1),
    .io_out_2(rand_exe_prng_103_io_out_2),
    .io_out_3(rand_exe_prng_103_io_out_3),
    .io_out_4(rand_exe_prng_103_io_out_4),
    .io_out_5(rand_exe_prng_103_io_out_5),
    .io_out_6(rand_exe_prng_103_io_out_6),
    .io_out_7(rand_exe_prng_103_io_out_7),
    .io_out_8(rand_exe_prng_103_io_out_8),
    .io_out_9(rand_exe_prng_103_io_out_9),
    .io_out_10(rand_exe_prng_103_io_out_10),
    .io_out_11(rand_exe_prng_103_io_out_11),
    .io_out_12(rand_exe_prng_103_io_out_12),
    .io_out_13(rand_exe_prng_103_io_out_13),
    .io_out_14(rand_exe_prng_103_io_out_14),
    .io_out_15(rand_exe_prng_103_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_104 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_104_clock),
    .reset(rand_exe_prng_104_reset),
    .io_out_0(rand_exe_prng_104_io_out_0),
    .io_out_1(rand_exe_prng_104_io_out_1),
    .io_out_2(rand_exe_prng_104_io_out_2),
    .io_out_3(rand_exe_prng_104_io_out_3),
    .io_out_4(rand_exe_prng_104_io_out_4),
    .io_out_5(rand_exe_prng_104_io_out_5),
    .io_out_6(rand_exe_prng_104_io_out_6),
    .io_out_7(rand_exe_prng_104_io_out_7),
    .io_out_8(rand_exe_prng_104_io_out_8),
    .io_out_9(rand_exe_prng_104_io_out_9),
    .io_out_10(rand_exe_prng_104_io_out_10),
    .io_out_11(rand_exe_prng_104_io_out_11),
    .io_out_12(rand_exe_prng_104_io_out_12),
    .io_out_13(rand_exe_prng_104_io_out_13),
    .io_out_14(rand_exe_prng_104_io_out_14),
    .io_out_15(rand_exe_prng_104_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_105 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_105_clock),
    .reset(rand_exe_prng_105_reset),
    .io_out_0(rand_exe_prng_105_io_out_0),
    .io_out_1(rand_exe_prng_105_io_out_1),
    .io_out_2(rand_exe_prng_105_io_out_2),
    .io_out_3(rand_exe_prng_105_io_out_3),
    .io_out_4(rand_exe_prng_105_io_out_4),
    .io_out_5(rand_exe_prng_105_io_out_5),
    .io_out_6(rand_exe_prng_105_io_out_6),
    .io_out_7(rand_exe_prng_105_io_out_7),
    .io_out_8(rand_exe_prng_105_io_out_8),
    .io_out_9(rand_exe_prng_105_io_out_9),
    .io_out_10(rand_exe_prng_105_io_out_10),
    .io_out_11(rand_exe_prng_105_io_out_11),
    .io_out_12(rand_exe_prng_105_io_out_12),
    .io_out_13(rand_exe_prng_105_io_out_13),
    .io_out_14(rand_exe_prng_105_io_out_14),
    .io_out_15(rand_exe_prng_105_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_106 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_106_clock),
    .reset(rand_exe_prng_106_reset),
    .io_out_0(rand_exe_prng_106_io_out_0),
    .io_out_1(rand_exe_prng_106_io_out_1),
    .io_out_2(rand_exe_prng_106_io_out_2),
    .io_out_3(rand_exe_prng_106_io_out_3),
    .io_out_4(rand_exe_prng_106_io_out_4),
    .io_out_5(rand_exe_prng_106_io_out_5),
    .io_out_6(rand_exe_prng_106_io_out_6),
    .io_out_7(rand_exe_prng_106_io_out_7),
    .io_out_8(rand_exe_prng_106_io_out_8),
    .io_out_9(rand_exe_prng_106_io_out_9),
    .io_out_10(rand_exe_prng_106_io_out_10),
    .io_out_11(rand_exe_prng_106_io_out_11),
    .io_out_12(rand_exe_prng_106_io_out_12),
    .io_out_13(rand_exe_prng_106_io_out_13),
    .io_out_14(rand_exe_prng_106_io_out_14),
    .io_out_15(rand_exe_prng_106_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_107 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_107_clock),
    .reset(rand_exe_prng_107_reset),
    .io_out_0(rand_exe_prng_107_io_out_0),
    .io_out_1(rand_exe_prng_107_io_out_1),
    .io_out_2(rand_exe_prng_107_io_out_2),
    .io_out_3(rand_exe_prng_107_io_out_3),
    .io_out_4(rand_exe_prng_107_io_out_4),
    .io_out_5(rand_exe_prng_107_io_out_5),
    .io_out_6(rand_exe_prng_107_io_out_6),
    .io_out_7(rand_exe_prng_107_io_out_7),
    .io_out_8(rand_exe_prng_107_io_out_8),
    .io_out_9(rand_exe_prng_107_io_out_9),
    .io_out_10(rand_exe_prng_107_io_out_10),
    .io_out_11(rand_exe_prng_107_io_out_11),
    .io_out_12(rand_exe_prng_107_io_out_12),
    .io_out_13(rand_exe_prng_107_io_out_13),
    .io_out_14(rand_exe_prng_107_io_out_14),
    .io_out_15(rand_exe_prng_107_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_108 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_108_clock),
    .reset(rand_exe_prng_108_reset),
    .io_out_0(rand_exe_prng_108_io_out_0),
    .io_out_1(rand_exe_prng_108_io_out_1),
    .io_out_2(rand_exe_prng_108_io_out_2),
    .io_out_3(rand_exe_prng_108_io_out_3),
    .io_out_4(rand_exe_prng_108_io_out_4),
    .io_out_5(rand_exe_prng_108_io_out_5),
    .io_out_6(rand_exe_prng_108_io_out_6),
    .io_out_7(rand_exe_prng_108_io_out_7),
    .io_out_8(rand_exe_prng_108_io_out_8),
    .io_out_9(rand_exe_prng_108_io_out_9),
    .io_out_10(rand_exe_prng_108_io_out_10),
    .io_out_11(rand_exe_prng_108_io_out_11),
    .io_out_12(rand_exe_prng_108_io_out_12),
    .io_out_13(rand_exe_prng_108_io_out_13),
    .io_out_14(rand_exe_prng_108_io_out_14),
    .io_out_15(rand_exe_prng_108_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_109 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_109_clock),
    .reset(rand_exe_prng_109_reset),
    .io_out_0(rand_exe_prng_109_io_out_0),
    .io_out_1(rand_exe_prng_109_io_out_1),
    .io_out_2(rand_exe_prng_109_io_out_2),
    .io_out_3(rand_exe_prng_109_io_out_3),
    .io_out_4(rand_exe_prng_109_io_out_4),
    .io_out_5(rand_exe_prng_109_io_out_5),
    .io_out_6(rand_exe_prng_109_io_out_6),
    .io_out_7(rand_exe_prng_109_io_out_7),
    .io_out_8(rand_exe_prng_109_io_out_8),
    .io_out_9(rand_exe_prng_109_io_out_9),
    .io_out_10(rand_exe_prng_109_io_out_10),
    .io_out_11(rand_exe_prng_109_io_out_11),
    .io_out_12(rand_exe_prng_109_io_out_12),
    .io_out_13(rand_exe_prng_109_io_out_13),
    .io_out_14(rand_exe_prng_109_io_out_14),
    .io_out_15(rand_exe_prng_109_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_110 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_110_clock),
    .reset(rand_exe_prng_110_reset),
    .io_out_0(rand_exe_prng_110_io_out_0),
    .io_out_1(rand_exe_prng_110_io_out_1),
    .io_out_2(rand_exe_prng_110_io_out_2),
    .io_out_3(rand_exe_prng_110_io_out_3),
    .io_out_4(rand_exe_prng_110_io_out_4),
    .io_out_5(rand_exe_prng_110_io_out_5),
    .io_out_6(rand_exe_prng_110_io_out_6),
    .io_out_7(rand_exe_prng_110_io_out_7),
    .io_out_8(rand_exe_prng_110_io_out_8),
    .io_out_9(rand_exe_prng_110_io_out_9),
    .io_out_10(rand_exe_prng_110_io_out_10),
    .io_out_11(rand_exe_prng_110_io_out_11),
    .io_out_12(rand_exe_prng_110_io_out_12),
    .io_out_13(rand_exe_prng_110_io_out_13),
    .io_out_14(rand_exe_prng_110_io_out_14),
    .io_out_15(rand_exe_prng_110_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_111 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_111_clock),
    .reset(rand_exe_prng_111_reset),
    .io_out_0(rand_exe_prng_111_io_out_0),
    .io_out_1(rand_exe_prng_111_io_out_1),
    .io_out_2(rand_exe_prng_111_io_out_2),
    .io_out_3(rand_exe_prng_111_io_out_3),
    .io_out_4(rand_exe_prng_111_io_out_4),
    .io_out_5(rand_exe_prng_111_io_out_5),
    .io_out_6(rand_exe_prng_111_io_out_6),
    .io_out_7(rand_exe_prng_111_io_out_7),
    .io_out_8(rand_exe_prng_111_io_out_8),
    .io_out_9(rand_exe_prng_111_io_out_9),
    .io_out_10(rand_exe_prng_111_io_out_10),
    .io_out_11(rand_exe_prng_111_io_out_11),
    .io_out_12(rand_exe_prng_111_io_out_12),
    .io_out_13(rand_exe_prng_111_io_out_13),
    .io_out_14(rand_exe_prng_111_io_out_14),
    .io_out_15(rand_exe_prng_111_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_112 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_112_clock),
    .reset(rand_exe_prng_112_reset),
    .io_out_0(rand_exe_prng_112_io_out_0),
    .io_out_1(rand_exe_prng_112_io_out_1),
    .io_out_2(rand_exe_prng_112_io_out_2),
    .io_out_3(rand_exe_prng_112_io_out_3),
    .io_out_4(rand_exe_prng_112_io_out_4),
    .io_out_5(rand_exe_prng_112_io_out_5),
    .io_out_6(rand_exe_prng_112_io_out_6),
    .io_out_7(rand_exe_prng_112_io_out_7),
    .io_out_8(rand_exe_prng_112_io_out_8),
    .io_out_9(rand_exe_prng_112_io_out_9),
    .io_out_10(rand_exe_prng_112_io_out_10),
    .io_out_11(rand_exe_prng_112_io_out_11),
    .io_out_12(rand_exe_prng_112_io_out_12),
    .io_out_13(rand_exe_prng_112_io_out_13),
    .io_out_14(rand_exe_prng_112_io_out_14),
    .io_out_15(rand_exe_prng_112_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_113 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_113_clock),
    .reset(rand_exe_prng_113_reset),
    .io_out_0(rand_exe_prng_113_io_out_0),
    .io_out_1(rand_exe_prng_113_io_out_1),
    .io_out_2(rand_exe_prng_113_io_out_2),
    .io_out_3(rand_exe_prng_113_io_out_3),
    .io_out_4(rand_exe_prng_113_io_out_4),
    .io_out_5(rand_exe_prng_113_io_out_5),
    .io_out_6(rand_exe_prng_113_io_out_6),
    .io_out_7(rand_exe_prng_113_io_out_7),
    .io_out_8(rand_exe_prng_113_io_out_8),
    .io_out_9(rand_exe_prng_113_io_out_9),
    .io_out_10(rand_exe_prng_113_io_out_10),
    .io_out_11(rand_exe_prng_113_io_out_11),
    .io_out_12(rand_exe_prng_113_io_out_12),
    .io_out_13(rand_exe_prng_113_io_out_13),
    .io_out_14(rand_exe_prng_113_io_out_14),
    .io_out_15(rand_exe_prng_113_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_114 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_114_clock),
    .reset(rand_exe_prng_114_reset),
    .io_out_0(rand_exe_prng_114_io_out_0),
    .io_out_1(rand_exe_prng_114_io_out_1),
    .io_out_2(rand_exe_prng_114_io_out_2),
    .io_out_3(rand_exe_prng_114_io_out_3),
    .io_out_4(rand_exe_prng_114_io_out_4),
    .io_out_5(rand_exe_prng_114_io_out_5),
    .io_out_6(rand_exe_prng_114_io_out_6),
    .io_out_7(rand_exe_prng_114_io_out_7),
    .io_out_8(rand_exe_prng_114_io_out_8),
    .io_out_9(rand_exe_prng_114_io_out_9),
    .io_out_10(rand_exe_prng_114_io_out_10),
    .io_out_11(rand_exe_prng_114_io_out_11),
    .io_out_12(rand_exe_prng_114_io_out_12),
    .io_out_13(rand_exe_prng_114_io_out_13),
    .io_out_14(rand_exe_prng_114_io_out_14),
    .io_out_15(rand_exe_prng_114_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_115 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_115_clock),
    .reset(rand_exe_prng_115_reset),
    .io_out_0(rand_exe_prng_115_io_out_0),
    .io_out_1(rand_exe_prng_115_io_out_1),
    .io_out_2(rand_exe_prng_115_io_out_2),
    .io_out_3(rand_exe_prng_115_io_out_3),
    .io_out_4(rand_exe_prng_115_io_out_4),
    .io_out_5(rand_exe_prng_115_io_out_5),
    .io_out_6(rand_exe_prng_115_io_out_6),
    .io_out_7(rand_exe_prng_115_io_out_7),
    .io_out_8(rand_exe_prng_115_io_out_8),
    .io_out_9(rand_exe_prng_115_io_out_9),
    .io_out_10(rand_exe_prng_115_io_out_10),
    .io_out_11(rand_exe_prng_115_io_out_11),
    .io_out_12(rand_exe_prng_115_io_out_12),
    .io_out_13(rand_exe_prng_115_io_out_13),
    .io_out_14(rand_exe_prng_115_io_out_14),
    .io_out_15(rand_exe_prng_115_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_116 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_116_clock),
    .reset(rand_exe_prng_116_reset),
    .io_out_0(rand_exe_prng_116_io_out_0),
    .io_out_1(rand_exe_prng_116_io_out_1),
    .io_out_2(rand_exe_prng_116_io_out_2),
    .io_out_3(rand_exe_prng_116_io_out_3),
    .io_out_4(rand_exe_prng_116_io_out_4),
    .io_out_5(rand_exe_prng_116_io_out_5),
    .io_out_6(rand_exe_prng_116_io_out_6),
    .io_out_7(rand_exe_prng_116_io_out_7),
    .io_out_8(rand_exe_prng_116_io_out_8),
    .io_out_9(rand_exe_prng_116_io_out_9),
    .io_out_10(rand_exe_prng_116_io_out_10),
    .io_out_11(rand_exe_prng_116_io_out_11),
    .io_out_12(rand_exe_prng_116_io_out_12),
    .io_out_13(rand_exe_prng_116_io_out_13),
    .io_out_14(rand_exe_prng_116_io_out_14),
    .io_out_15(rand_exe_prng_116_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_117 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_117_clock),
    .reset(rand_exe_prng_117_reset),
    .io_out_0(rand_exe_prng_117_io_out_0),
    .io_out_1(rand_exe_prng_117_io_out_1),
    .io_out_2(rand_exe_prng_117_io_out_2),
    .io_out_3(rand_exe_prng_117_io_out_3),
    .io_out_4(rand_exe_prng_117_io_out_4),
    .io_out_5(rand_exe_prng_117_io_out_5),
    .io_out_6(rand_exe_prng_117_io_out_6),
    .io_out_7(rand_exe_prng_117_io_out_7),
    .io_out_8(rand_exe_prng_117_io_out_8),
    .io_out_9(rand_exe_prng_117_io_out_9),
    .io_out_10(rand_exe_prng_117_io_out_10),
    .io_out_11(rand_exe_prng_117_io_out_11),
    .io_out_12(rand_exe_prng_117_io_out_12),
    .io_out_13(rand_exe_prng_117_io_out_13),
    .io_out_14(rand_exe_prng_117_io_out_14),
    .io_out_15(rand_exe_prng_117_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_118 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_118_clock),
    .reset(rand_exe_prng_118_reset),
    .io_out_0(rand_exe_prng_118_io_out_0),
    .io_out_1(rand_exe_prng_118_io_out_1),
    .io_out_2(rand_exe_prng_118_io_out_2),
    .io_out_3(rand_exe_prng_118_io_out_3),
    .io_out_4(rand_exe_prng_118_io_out_4),
    .io_out_5(rand_exe_prng_118_io_out_5),
    .io_out_6(rand_exe_prng_118_io_out_6),
    .io_out_7(rand_exe_prng_118_io_out_7),
    .io_out_8(rand_exe_prng_118_io_out_8),
    .io_out_9(rand_exe_prng_118_io_out_9),
    .io_out_10(rand_exe_prng_118_io_out_10),
    .io_out_11(rand_exe_prng_118_io_out_11),
    .io_out_12(rand_exe_prng_118_io_out_12),
    .io_out_13(rand_exe_prng_118_io_out_13),
    .io_out_14(rand_exe_prng_118_io_out_14),
    .io_out_15(rand_exe_prng_118_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_119 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_119_clock),
    .reset(rand_exe_prng_119_reset),
    .io_out_0(rand_exe_prng_119_io_out_0),
    .io_out_1(rand_exe_prng_119_io_out_1),
    .io_out_2(rand_exe_prng_119_io_out_2),
    .io_out_3(rand_exe_prng_119_io_out_3),
    .io_out_4(rand_exe_prng_119_io_out_4),
    .io_out_5(rand_exe_prng_119_io_out_5),
    .io_out_6(rand_exe_prng_119_io_out_6),
    .io_out_7(rand_exe_prng_119_io_out_7),
    .io_out_8(rand_exe_prng_119_io_out_8),
    .io_out_9(rand_exe_prng_119_io_out_9),
    .io_out_10(rand_exe_prng_119_io_out_10),
    .io_out_11(rand_exe_prng_119_io_out_11),
    .io_out_12(rand_exe_prng_119_io_out_12),
    .io_out_13(rand_exe_prng_119_io_out_13),
    .io_out_14(rand_exe_prng_119_io_out_14),
    .io_out_15(rand_exe_prng_119_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_120 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_120_clock),
    .reset(rand_exe_prng_120_reset),
    .io_out_0(rand_exe_prng_120_io_out_0),
    .io_out_1(rand_exe_prng_120_io_out_1),
    .io_out_2(rand_exe_prng_120_io_out_2),
    .io_out_3(rand_exe_prng_120_io_out_3),
    .io_out_4(rand_exe_prng_120_io_out_4),
    .io_out_5(rand_exe_prng_120_io_out_5),
    .io_out_6(rand_exe_prng_120_io_out_6),
    .io_out_7(rand_exe_prng_120_io_out_7),
    .io_out_8(rand_exe_prng_120_io_out_8),
    .io_out_9(rand_exe_prng_120_io_out_9),
    .io_out_10(rand_exe_prng_120_io_out_10),
    .io_out_11(rand_exe_prng_120_io_out_11),
    .io_out_12(rand_exe_prng_120_io_out_12),
    .io_out_13(rand_exe_prng_120_io_out_13),
    .io_out_14(rand_exe_prng_120_io_out_14),
    .io_out_15(rand_exe_prng_120_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_121 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_121_clock),
    .reset(rand_exe_prng_121_reset),
    .io_out_0(rand_exe_prng_121_io_out_0),
    .io_out_1(rand_exe_prng_121_io_out_1),
    .io_out_2(rand_exe_prng_121_io_out_2),
    .io_out_3(rand_exe_prng_121_io_out_3),
    .io_out_4(rand_exe_prng_121_io_out_4),
    .io_out_5(rand_exe_prng_121_io_out_5),
    .io_out_6(rand_exe_prng_121_io_out_6),
    .io_out_7(rand_exe_prng_121_io_out_7),
    .io_out_8(rand_exe_prng_121_io_out_8),
    .io_out_9(rand_exe_prng_121_io_out_9),
    .io_out_10(rand_exe_prng_121_io_out_10),
    .io_out_11(rand_exe_prng_121_io_out_11),
    .io_out_12(rand_exe_prng_121_io_out_12),
    .io_out_13(rand_exe_prng_121_io_out_13),
    .io_out_14(rand_exe_prng_121_io_out_14),
    .io_out_15(rand_exe_prng_121_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_122 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_122_clock),
    .reset(rand_exe_prng_122_reset),
    .io_out_0(rand_exe_prng_122_io_out_0),
    .io_out_1(rand_exe_prng_122_io_out_1),
    .io_out_2(rand_exe_prng_122_io_out_2),
    .io_out_3(rand_exe_prng_122_io_out_3),
    .io_out_4(rand_exe_prng_122_io_out_4),
    .io_out_5(rand_exe_prng_122_io_out_5),
    .io_out_6(rand_exe_prng_122_io_out_6),
    .io_out_7(rand_exe_prng_122_io_out_7),
    .io_out_8(rand_exe_prng_122_io_out_8),
    .io_out_9(rand_exe_prng_122_io_out_9),
    .io_out_10(rand_exe_prng_122_io_out_10),
    .io_out_11(rand_exe_prng_122_io_out_11),
    .io_out_12(rand_exe_prng_122_io_out_12),
    .io_out_13(rand_exe_prng_122_io_out_13),
    .io_out_14(rand_exe_prng_122_io_out_14),
    .io_out_15(rand_exe_prng_122_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_123 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_123_clock),
    .reset(rand_exe_prng_123_reset),
    .io_out_0(rand_exe_prng_123_io_out_0),
    .io_out_1(rand_exe_prng_123_io_out_1),
    .io_out_2(rand_exe_prng_123_io_out_2),
    .io_out_3(rand_exe_prng_123_io_out_3),
    .io_out_4(rand_exe_prng_123_io_out_4),
    .io_out_5(rand_exe_prng_123_io_out_5),
    .io_out_6(rand_exe_prng_123_io_out_6),
    .io_out_7(rand_exe_prng_123_io_out_7),
    .io_out_8(rand_exe_prng_123_io_out_8),
    .io_out_9(rand_exe_prng_123_io_out_9),
    .io_out_10(rand_exe_prng_123_io_out_10),
    .io_out_11(rand_exe_prng_123_io_out_11),
    .io_out_12(rand_exe_prng_123_io_out_12),
    .io_out_13(rand_exe_prng_123_io_out_13),
    .io_out_14(rand_exe_prng_123_io_out_14),
    .io_out_15(rand_exe_prng_123_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_124 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_124_clock),
    .reset(rand_exe_prng_124_reset),
    .io_out_0(rand_exe_prng_124_io_out_0),
    .io_out_1(rand_exe_prng_124_io_out_1),
    .io_out_2(rand_exe_prng_124_io_out_2),
    .io_out_3(rand_exe_prng_124_io_out_3),
    .io_out_4(rand_exe_prng_124_io_out_4),
    .io_out_5(rand_exe_prng_124_io_out_5),
    .io_out_6(rand_exe_prng_124_io_out_6),
    .io_out_7(rand_exe_prng_124_io_out_7),
    .io_out_8(rand_exe_prng_124_io_out_8),
    .io_out_9(rand_exe_prng_124_io_out_9),
    .io_out_10(rand_exe_prng_124_io_out_10),
    .io_out_11(rand_exe_prng_124_io_out_11),
    .io_out_12(rand_exe_prng_124_io_out_12),
    .io_out_13(rand_exe_prng_124_io_out_13),
    .io_out_14(rand_exe_prng_124_io_out_14),
    .io_out_15(rand_exe_prng_124_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_125 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_125_clock),
    .reset(rand_exe_prng_125_reset),
    .io_out_0(rand_exe_prng_125_io_out_0),
    .io_out_1(rand_exe_prng_125_io_out_1),
    .io_out_2(rand_exe_prng_125_io_out_2),
    .io_out_3(rand_exe_prng_125_io_out_3),
    .io_out_4(rand_exe_prng_125_io_out_4),
    .io_out_5(rand_exe_prng_125_io_out_5),
    .io_out_6(rand_exe_prng_125_io_out_6),
    .io_out_7(rand_exe_prng_125_io_out_7),
    .io_out_8(rand_exe_prng_125_io_out_8),
    .io_out_9(rand_exe_prng_125_io_out_9),
    .io_out_10(rand_exe_prng_125_io_out_10),
    .io_out_11(rand_exe_prng_125_io_out_11),
    .io_out_12(rand_exe_prng_125_io_out_12),
    .io_out_13(rand_exe_prng_125_io_out_13),
    .io_out_14(rand_exe_prng_125_io_out_14),
    .io_out_15(rand_exe_prng_125_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_126 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_126_clock),
    .reset(rand_exe_prng_126_reset),
    .io_out_0(rand_exe_prng_126_io_out_0),
    .io_out_1(rand_exe_prng_126_io_out_1),
    .io_out_2(rand_exe_prng_126_io_out_2),
    .io_out_3(rand_exe_prng_126_io_out_3),
    .io_out_4(rand_exe_prng_126_io_out_4),
    .io_out_5(rand_exe_prng_126_io_out_5),
    .io_out_6(rand_exe_prng_126_io_out_6),
    .io_out_7(rand_exe_prng_126_io_out_7),
    .io_out_8(rand_exe_prng_126_io_out_8),
    .io_out_9(rand_exe_prng_126_io_out_9),
    .io_out_10(rand_exe_prng_126_io_out_10),
    .io_out_11(rand_exe_prng_126_io_out_11),
    .io_out_12(rand_exe_prng_126_io_out_12),
    .io_out_13(rand_exe_prng_126_io_out_13),
    .io_out_14(rand_exe_prng_126_io_out_14),
    .io_out_15(rand_exe_prng_126_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_127 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_127_clock),
    .reset(rand_exe_prng_127_reset),
    .io_out_0(rand_exe_prng_127_io_out_0),
    .io_out_1(rand_exe_prng_127_io_out_1),
    .io_out_2(rand_exe_prng_127_io_out_2),
    .io_out_3(rand_exe_prng_127_io_out_3),
    .io_out_4(rand_exe_prng_127_io_out_4),
    .io_out_5(rand_exe_prng_127_io_out_5),
    .io_out_6(rand_exe_prng_127_io_out_6),
    .io_out_7(rand_exe_prng_127_io_out_7),
    .io_out_8(rand_exe_prng_127_io_out_8),
    .io_out_9(rand_exe_prng_127_io_out_9),
    .io_out_10(rand_exe_prng_127_io_out_10),
    .io_out_11(rand_exe_prng_127_io_out_11),
    .io_out_12(rand_exe_prng_127_io_out_12),
    .io_out_13(rand_exe_prng_127_io_out_13),
    .io_out_14(rand_exe_prng_127_io_out_14),
    .io_out_15(rand_exe_prng_127_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_128 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_128_clock),
    .reset(rand_exe_prng_128_reset),
    .io_out_0(rand_exe_prng_128_io_out_0),
    .io_out_1(rand_exe_prng_128_io_out_1),
    .io_out_2(rand_exe_prng_128_io_out_2),
    .io_out_3(rand_exe_prng_128_io_out_3),
    .io_out_4(rand_exe_prng_128_io_out_4),
    .io_out_5(rand_exe_prng_128_io_out_5),
    .io_out_6(rand_exe_prng_128_io_out_6),
    .io_out_7(rand_exe_prng_128_io_out_7),
    .io_out_8(rand_exe_prng_128_io_out_8),
    .io_out_9(rand_exe_prng_128_io_out_9),
    .io_out_10(rand_exe_prng_128_io_out_10),
    .io_out_11(rand_exe_prng_128_io_out_11),
    .io_out_12(rand_exe_prng_128_io_out_12),
    .io_out_13(rand_exe_prng_128_io_out_13),
    .io_out_14(rand_exe_prng_128_io_out_14),
    .io_out_15(rand_exe_prng_128_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_129 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_129_clock),
    .reset(rand_exe_prng_129_reset),
    .io_out_0(rand_exe_prng_129_io_out_0),
    .io_out_1(rand_exe_prng_129_io_out_1),
    .io_out_2(rand_exe_prng_129_io_out_2),
    .io_out_3(rand_exe_prng_129_io_out_3),
    .io_out_4(rand_exe_prng_129_io_out_4),
    .io_out_5(rand_exe_prng_129_io_out_5),
    .io_out_6(rand_exe_prng_129_io_out_6),
    .io_out_7(rand_exe_prng_129_io_out_7),
    .io_out_8(rand_exe_prng_129_io_out_8),
    .io_out_9(rand_exe_prng_129_io_out_9),
    .io_out_10(rand_exe_prng_129_io_out_10),
    .io_out_11(rand_exe_prng_129_io_out_11),
    .io_out_12(rand_exe_prng_129_io_out_12),
    .io_out_13(rand_exe_prng_129_io_out_13),
    .io_out_14(rand_exe_prng_129_io_out_14),
    .io_out_15(rand_exe_prng_129_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_130 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_130_clock),
    .reset(rand_exe_prng_130_reset),
    .io_out_0(rand_exe_prng_130_io_out_0),
    .io_out_1(rand_exe_prng_130_io_out_1),
    .io_out_2(rand_exe_prng_130_io_out_2),
    .io_out_3(rand_exe_prng_130_io_out_3),
    .io_out_4(rand_exe_prng_130_io_out_4),
    .io_out_5(rand_exe_prng_130_io_out_5),
    .io_out_6(rand_exe_prng_130_io_out_6),
    .io_out_7(rand_exe_prng_130_io_out_7),
    .io_out_8(rand_exe_prng_130_io_out_8),
    .io_out_9(rand_exe_prng_130_io_out_9),
    .io_out_10(rand_exe_prng_130_io_out_10),
    .io_out_11(rand_exe_prng_130_io_out_11),
    .io_out_12(rand_exe_prng_130_io_out_12),
    .io_out_13(rand_exe_prng_130_io_out_13),
    .io_out_14(rand_exe_prng_130_io_out_14),
    .io_out_15(rand_exe_prng_130_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_131 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_131_clock),
    .reset(rand_exe_prng_131_reset),
    .io_out_0(rand_exe_prng_131_io_out_0),
    .io_out_1(rand_exe_prng_131_io_out_1),
    .io_out_2(rand_exe_prng_131_io_out_2),
    .io_out_3(rand_exe_prng_131_io_out_3),
    .io_out_4(rand_exe_prng_131_io_out_4),
    .io_out_5(rand_exe_prng_131_io_out_5),
    .io_out_6(rand_exe_prng_131_io_out_6),
    .io_out_7(rand_exe_prng_131_io_out_7),
    .io_out_8(rand_exe_prng_131_io_out_8),
    .io_out_9(rand_exe_prng_131_io_out_9),
    .io_out_10(rand_exe_prng_131_io_out_10),
    .io_out_11(rand_exe_prng_131_io_out_11),
    .io_out_12(rand_exe_prng_131_io_out_12),
    .io_out_13(rand_exe_prng_131_io_out_13),
    .io_out_14(rand_exe_prng_131_io_out_14),
    .io_out_15(rand_exe_prng_131_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_132 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_132_clock),
    .reset(rand_exe_prng_132_reset),
    .io_out_0(rand_exe_prng_132_io_out_0),
    .io_out_1(rand_exe_prng_132_io_out_1),
    .io_out_2(rand_exe_prng_132_io_out_2),
    .io_out_3(rand_exe_prng_132_io_out_3),
    .io_out_4(rand_exe_prng_132_io_out_4),
    .io_out_5(rand_exe_prng_132_io_out_5),
    .io_out_6(rand_exe_prng_132_io_out_6),
    .io_out_7(rand_exe_prng_132_io_out_7),
    .io_out_8(rand_exe_prng_132_io_out_8),
    .io_out_9(rand_exe_prng_132_io_out_9),
    .io_out_10(rand_exe_prng_132_io_out_10),
    .io_out_11(rand_exe_prng_132_io_out_11),
    .io_out_12(rand_exe_prng_132_io_out_12),
    .io_out_13(rand_exe_prng_132_io_out_13),
    .io_out_14(rand_exe_prng_132_io_out_14),
    .io_out_15(rand_exe_prng_132_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_133 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_133_clock),
    .reset(rand_exe_prng_133_reset),
    .io_out_0(rand_exe_prng_133_io_out_0),
    .io_out_1(rand_exe_prng_133_io_out_1),
    .io_out_2(rand_exe_prng_133_io_out_2),
    .io_out_3(rand_exe_prng_133_io_out_3),
    .io_out_4(rand_exe_prng_133_io_out_4),
    .io_out_5(rand_exe_prng_133_io_out_5),
    .io_out_6(rand_exe_prng_133_io_out_6),
    .io_out_7(rand_exe_prng_133_io_out_7),
    .io_out_8(rand_exe_prng_133_io_out_8),
    .io_out_9(rand_exe_prng_133_io_out_9),
    .io_out_10(rand_exe_prng_133_io_out_10),
    .io_out_11(rand_exe_prng_133_io_out_11),
    .io_out_12(rand_exe_prng_133_io_out_12),
    .io_out_13(rand_exe_prng_133_io_out_13),
    .io_out_14(rand_exe_prng_133_io_out_14),
    .io_out_15(rand_exe_prng_133_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_134 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_134_clock),
    .reset(rand_exe_prng_134_reset),
    .io_out_0(rand_exe_prng_134_io_out_0),
    .io_out_1(rand_exe_prng_134_io_out_1),
    .io_out_2(rand_exe_prng_134_io_out_2),
    .io_out_3(rand_exe_prng_134_io_out_3),
    .io_out_4(rand_exe_prng_134_io_out_4),
    .io_out_5(rand_exe_prng_134_io_out_5),
    .io_out_6(rand_exe_prng_134_io_out_6),
    .io_out_7(rand_exe_prng_134_io_out_7),
    .io_out_8(rand_exe_prng_134_io_out_8),
    .io_out_9(rand_exe_prng_134_io_out_9),
    .io_out_10(rand_exe_prng_134_io_out_10),
    .io_out_11(rand_exe_prng_134_io_out_11),
    .io_out_12(rand_exe_prng_134_io_out_12),
    .io_out_13(rand_exe_prng_134_io_out_13),
    .io_out_14(rand_exe_prng_134_io_out_14),
    .io_out_15(rand_exe_prng_134_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_135 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_135_clock),
    .reset(rand_exe_prng_135_reset),
    .io_out_0(rand_exe_prng_135_io_out_0),
    .io_out_1(rand_exe_prng_135_io_out_1),
    .io_out_2(rand_exe_prng_135_io_out_2),
    .io_out_3(rand_exe_prng_135_io_out_3),
    .io_out_4(rand_exe_prng_135_io_out_4),
    .io_out_5(rand_exe_prng_135_io_out_5),
    .io_out_6(rand_exe_prng_135_io_out_6),
    .io_out_7(rand_exe_prng_135_io_out_7),
    .io_out_8(rand_exe_prng_135_io_out_8),
    .io_out_9(rand_exe_prng_135_io_out_9),
    .io_out_10(rand_exe_prng_135_io_out_10),
    .io_out_11(rand_exe_prng_135_io_out_11),
    .io_out_12(rand_exe_prng_135_io_out_12),
    .io_out_13(rand_exe_prng_135_io_out_13),
    .io_out_14(rand_exe_prng_135_io_out_14),
    .io_out_15(rand_exe_prng_135_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_136 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_136_clock),
    .reset(rand_exe_prng_136_reset),
    .io_out_0(rand_exe_prng_136_io_out_0),
    .io_out_1(rand_exe_prng_136_io_out_1),
    .io_out_2(rand_exe_prng_136_io_out_2),
    .io_out_3(rand_exe_prng_136_io_out_3),
    .io_out_4(rand_exe_prng_136_io_out_4),
    .io_out_5(rand_exe_prng_136_io_out_5),
    .io_out_6(rand_exe_prng_136_io_out_6),
    .io_out_7(rand_exe_prng_136_io_out_7),
    .io_out_8(rand_exe_prng_136_io_out_8),
    .io_out_9(rand_exe_prng_136_io_out_9),
    .io_out_10(rand_exe_prng_136_io_out_10),
    .io_out_11(rand_exe_prng_136_io_out_11),
    .io_out_12(rand_exe_prng_136_io_out_12),
    .io_out_13(rand_exe_prng_136_io_out_13),
    .io_out_14(rand_exe_prng_136_io_out_14),
    .io_out_15(rand_exe_prng_136_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_137 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_137_clock),
    .reset(rand_exe_prng_137_reset),
    .io_out_0(rand_exe_prng_137_io_out_0),
    .io_out_1(rand_exe_prng_137_io_out_1),
    .io_out_2(rand_exe_prng_137_io_out_2),
    .io_out_3(rand_exe_prng_137_io_out_3),
    .io_out_4(rand_exe_prng_137_io_out_4),
    .io_out_5(rand_exe_prng_137_io_out_5),
    .io_out_6(rand_exe_prng_137_io_out_6),
    .io_out_7(rand_exe_prng_137_io_out_7),
    .io_out_8(rand_exe_prng_137_io_out_8),
    .io_out_9(rand_exe_prng_137_io_out_9),
    .io_out_10(rand_exe_prng_137_io_out_10),
    .io_out_11(rand_exe_prng_137_io_out_11),
    .io_out_12(rand_exe_prng_137_io_out_12),
    .io_out_13(rand_exe_prng_137_io_out_13),
    .io_out_14(rand_exe_prng_137_io_out_14),
    .io_out_15(rand_exe_prng_137_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_138 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_138_clock),
    .reset(rand_exe_prng_138_reset),
    .io_out_0(rand_exe_prng_138_io_out_0),
    .io_out_1(rand_exe_prng_138_io_out_1),
    .io_out_2(rand_exe_prng_138_io_out_2),
    .io_out_3(rand_exe_prng_138_io_out_3),
    .io_out_4(rand_exe_prng_138_io_out_4),
    .io_out_5(rand_exe_prng_138_io_out_5),
    .io_out_6(rand_exe_prng_138_io_out_6),
    .io_out_7(rand_exe_prng_138_io_out_7),
    .io_out_8(rand_exe_prng_138_io_out_8),
    .io_out_9(rand_exe_prng_138_io_out_9),
    .io_out_10(rand_exe_prng_138_io_out_10),
    .io_out_11(rand_exe_prng_138_io_out_11),
    .io_out_12(rand_exe_prng_138_io_out_12),
    .io_out_13(rand_exe_prng_138_io_out_13),
    .io_out_14(rand_exe_prng_138_io_out_14),
    .io_out_15(rand_exe_prng_138_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_139 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_139_clock),
    .reset(rand_exe_prng_139_reset),
    .io_out_0(rand_exe_prng_139_io_out_0),
    .io_out_1(rand_exe_prng_139_io_out_1),
    .io_out_2(rand_exe_prng_139_io_out_2),
    .io_out_3(rand_exe_prng_139_io_out_3),
    .io_out_4(rand_exe_prng_139_io_out_4),
    .io_out_5(rand_exe_prng_139_io_out_5),
    .io_out_6(rand_exe_prng_139_io_out_6),
    .io_out_7(rand_exe_prng_139_io_out_7),
    .io_out_8(rand_exe_prng_139_io_out_8),
    .io_out_9(rand_exe_prng_139_io_out_9),
    .io_out_10(rand_exe_prng_139_io_out_10),
    .io_out_11(rand_exe_prng_139_io_out_11),
    .io_out_12(rand_exe_prng_139_io_out_12),
    .io_out_13(rand_exe_prng_139_io_out_13),
    .io_out_14(rand_exe_prng_139_io_out_14),
    .io_out_15(rand_exe_prng_139_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_140 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_140_clock),
    .reset(rand_exe_prng_140_reset),
    .io_out_0(rand_exe_prng_140_io_out_0),
    .io_out_1(rand_exe_prng_140_io_out_1),
    .io_out_2(rand_exe_prng_140_io_out_2),
    .io_out_3(rand_exe_prng_140_io_out_3),
    .io_out_4(rand_exe_prng_140_io_out_4),
    .io_out_5(rand_exe_prng_140_io_out_5),
    .io_out_6(rand_exe_prng_140_io_out_6),
    .io_out_7(rand_exe_prng_140_io_out_7),
    .io_out_8(rand_exe_prng_140_io_out_8),
    .io_out_9(rand_exe_prng_140_io_out_9),
    .io_out_10(rand_exe_prng_140_io_out_10),
    .io_out_11(rand_exe_prng_140_io_out_11),
    .io_out_12(rand_exe_prng_140_io_out_12),
    .io_out_13(rand_exe_prng_140_io_out_13),
    .io_out_14(rand_exe_prng_140_io_out_14),
    .io_out_15(rand_exe_prng_140_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_141 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_141_clock),
    .reset(rand_exe_prng_141_reset),
    .io_out_0(rand_exe_prng_141_io_out_0),
    .io_out_1(rand_exe_prng_141_io_out_1),
    .io_out_2(rand_exe_prng_141_io_out_2),
    .io_out_3(rand_exe_prng_141_io_out_3),
    .io_out_4(rand_exe_prng_141_io_out_4),
    .io_out_5(rand_exe_prng_141_io_out_5),
    .io_out_6(rand_exe_prng_141_io_out_6),
    .io_out_7(rand_exe_prng_141_io_out_7),
    .io_out_8(rand_exe_prng_141_io_out_8),
    .io_out_9(rand_exe_prng_141_io_out_9),
    .io_out_10(rand_exe_prng_141_io_out_10),
    .io_out_11(rand_exe_prng_141_io_out_11),
    .io_out_12(rand_exe_prng_141_io_out_12),
    .io_out_13(rand_exe_prng_141_io_out_13),
    .io_out_14(rand_exe_prng_141_io_out_14),
    .io_out_15(rand_exe_prng_141_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_142 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_142_clock),
    .reset(rand_exe_prng_142_reset),
    .io_out_0(rand_exe_prng_142_io_out_0),
    .io_out_1(rand_exe_prng_142_io_out_1),
    .io_out_2(rand_exe_prng_142_io_out_2),
    .io_out_3(rand_exe_prng_142_io_out_3),
    .io_out_4(rand_exe_prng_142_io_out_4),
    .io_out_5(rand_exe_prng_142_io_out_5),
    .io_out_6(rand_exe_prng_142_io_out_6),
    .io_out_7(rand_exe_prng_142_io_out_7),
    .io_out_8(rand_exe_prng_142_io_out_8),
    .io_out_9(rand_exe_prng_142_io_out_9),
    .io_out_10(rand_exe_prng_142_io_out_10),
    .io_out_11(rand_exe_prng_142_io_out_11),
    .io_out_12(rand_exe_prng_142_io_out_12),
    .io_out_13(rand_exe_prng_142_io_out_13),
    .io_out_14(rand_exe_prng_142_io_out_14),
    .io_out_15(rand_exe_prng_142_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_143 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_143_clock),
    .reset(rand_exe_prng_143_reset),
    .io_out_0(rand_exe_prng_143_io_out_0),
    .io_out_1(rand_exe_prng_143_io_out_1),
    .io_out_2(rand_exe_prng_143_io_out_2),
    .io_out_3(rand_exe_prng_143_io_out_3),
    .io_out_4(rand_exe_prng_143_io_out_4),
    .io_out_5(rand_exe_prng_143_io_out_5),
    .io_out_6(rand_exe_prng_143_io_out_6),
    .io_out_7(rand_exe_prng_143_io_out_7),
    .io_out_8(rand_exe_prng_143_io_out_8),
    .io_out_9(rand_exe_prng_143_io_out_9),
    .io_out_10(rand_exe_prng_143_io_out_10),
    .io_out_11(rand_exe_prng_143_io_out_11),
    .io_out_12(rand_exe_prng_143_io_out_12),
    .io_out_13(rand_exe_prng_143_io_out_13),
    .io_out_14(rand_exe_prng_143_io_out_14),
    .io_out_15(rand_exe_prng_143_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_144 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_144_clock),
    .reset(rand_exe_prng_144_reset),
    .io_out_0(rand_exe_prng_144_io_out_0),
    .io_out_1(rand_exe_prng_144_io_out_1),
    .io_out_2(rand_exe_prng_144_io_out_2),
    .io_out_3(rand_exe_prng_144_io_out_3),
    .io_out_4(rand_exe_prng_144_io_out_4),
    .io_out_5(rand_exe_prng_144_io_out_5),
    .io_out_6(rand_exe_prng_144_io_out_6),
    .io_out_7(rand_exe_prng_144_io_out_7),
    .io_out_8(rand_exe_prng_144_io_out_8),
    .io_out_9(rand_exe_prng_144_io_out_9),
    .io_out_10(rand_exe_prng_144_io_out_10),
    .io_out_11(rand_exe_prng_144_io_out_11),
    .io_out_12(rand_exe_prng_144_io_out_12),
    .io_out_13(rand_exe_prng_144_io_out_13),
    .io_out_14(rand_exe_prng_144_io_out_14),
    .io_out_15(rand_exe_prng_144_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_145 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_145_clock),
    .reset(rand_exe_prng_145_reset),
    .io_out_0(rand_exe_prng_145_io_out_0),
    .io_out_1(rand_exe_prng_145_io_out_1),
    .io_out_2(rand_exe_prng_145_io_out_2),
    .io_out_3(rand_exe_prng_145_io_out_3),
    .io_out_4(rand_exe_prng_145_io_out_4),
    .io_out_5(rand_exe_prng_145_io_out_5),
    .io_out_6(rand_exe_prng_145_io_out_6),
    .io_out_7(rand_exe_prng_145_io_out_7),
    .io_out_8(rand_exe_prng_145_io_out_8),
    .io_out_9(rand_exe_prng_145_io_out_9),
    .io_out_10(rand_exe_prng_145_io_out_10),
    .io_out_11(rand_exe_prng_145_io_out_11),
    .io_out_12(rand_exe_prng_145_io_out_12),
    .io_out_13(rand_exe_prng_145_io_out_13),
    .io_out_14(rand_exe_prng_145_io_out_14),
    .io_out_15(rand_exe_prng_145_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_146 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_146_clock),
    .reset(rand_exe_prng_146_reset),
    .io_out_0(rand_exe_prng_146_io_out_0),
    .io_out_1(rand_exe_prng_146_io_out_1),
    .io_out_2(rand_exe_prng_146_io_out_2),
    .io_out_3(rand_exe_prng_146_io_out_3),
    .io_out_4(rand_exe_prng_146_io_out_4),
    .io_out_5(rand_exe_prng_146_io_out_5),
    .io_out_6(rand_exe_prng_146_io_out_6),
    .io_out_7(rand_exe_prng_146_io_out_7),
    .io_out_8(rand_exe_prng_146_io_out_8),
    .io_out_9(rand_exe_prng_146_io_out_9),
    .io_out_10(rand_exe_prng_146_io_out_10),
    .io_out_11(rand_exe_prng_146_io_out_11),
    .io_out_12(rand_exe_prng_146_io_out_12),
    .io_out_13(rand_exe_prng_146_io_out_13),
    .io_out_14(rand_exe_prng_146_io_out_14),
    .io_out_15(rand_exe_prng_146_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_147 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_147_clock),
    .reset(rand_exe_prng_147_reset),
    .io_out_0(rand_exe_prng_147_io_out_0),
    .io_out_1(rand_exe_prng_147_io_out_1),
    .io_out_2(rand_exe_prng_147_io_out_2),
    .io_out_3(rand_exe_prng_147_io_out_3),
    .io_out_4(rand_exe_prng_147_io_out_4),
    .io_out_5(rand_exe_prng_147_io_out_5),
    .io_out_6(rand_exe_prng_147_io_out_6),
    .io_out_7(rand_exe_prng_147_io_out_7),
    .io_out_8(rand_exe_prng_147_io_out_8),
    .io_out_9(rand_exe_prng_147_io_out_9),
    .io_out_10(rand_exe_prng_147_io_out_10),
    .io_out_11(rand_exe_prng_147_io_out_11),
    .io_out_12(rand_exe_prng_147_io_out_12),
    .io_out_13(rand_exe_prng_147_io_out_13),
    .io_out_14(rand_exe_prng_147_io_out_14),
    .io_out_15(rand_exe_prng_147_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_148 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_148_clock),
    .reset(rand_exe_prng_148_reset),
    .io_out_0(rand_exe_prng_148_io_out_0),
    .io_out_1(rand_exe_prng_148_io_out_1),
    .io_out_2(rand_exe_prng_148_io_out_2),
    .io_out_3(rand_exe_prng_148_io_out_3),
    .io_out_4(rand_exe_prng_148_io_out_4),
    .io_out_5(rand_exe_prng_148_io_out_5),
    .io_out_6(rand_exe_prng_148_io_out_6),
    .io_out_7(rand_exe_prng_148_io_out_7),
    .io_out_8(rand_exe_prng_148_io_out_8),
    .io_out_9(rand_exe_prng_148_io_out_9),
    .io_out_10(rand_exe_prng_148_io_out_10),
    .io_out_11(rand_exe_prng_148_io_out_11),
    .io_out_12(rand_exe_prng_148_io_out_12),
    .io_out_13(rand_exe_prng_148_io_out_13),
    .io_out_14(rand_exe_prng_148_io_out_14),
    .io_out_15(rand_exe_prng_148_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_149 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_149_clock),
    .reset(rand_exe_prng_149_reset),
    .io_out_0(rand_exe_prng_149_io_out_0),
    .io_out_1(rand_exe_prng_149_io_out_1),
    .io_out_2(rand_exe_prng_149_io_out_2),
    .io_out_3(rand_exe_prng_149_io_out_3),
    .io_out_4(rand_exe_prng_149_io_out_4),
    .io_out_5(rand_exe_prng_149_io_out_5),
    .io_out_6(rand_exe_prng_149_io_out_6),
    .io_out_7(rand_exe_prng_149_io_out_7),
    .io_out_8(rand_exe_prng_149_io_out_8),
    .io_out_9(rand_exe_prng_149_io_out_9),
    .io_out_10(rand_exe_prng_149_io_out_10),
    .io_out_11(rand_exe_prng_149_io_out_11),
    .io_out_12(rand_exe_prng_149_io_out_12),
    .io_out_13(rand_exe_prng_149_io_out_13),
    .io_out_14(rand_exe_prng_149_io_out_14),
    .io_out_15(rand_exe_prng_149_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_150 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_150_clock),
    .reset(rand_exe_prng_150_reset),
    .io_out_0(rand_exe_prng_150_io_out_0),
    .io_out_1(rand_exe_prng_150_io_out_1),
    .io_out_2(rand_exe_prng_150_io_out_2),
    .io_out_3(rand_exe_prng_150_io_out_3),
    .io_out_4(rand_exe_prng_150_io_out_4),
    .io_out_5(rand_exe_prng_150_io_out_5),
    .io_out_6(rand_exe_prng_150_io_out_6),
    .io_out_7(rand_exe_prng_150_io_out_7),
    .io_out_8(rand_exe_prng_150_io_out_8),
    .io_out_9(rand_exe_prng_150_io_out_9),
    .io_out_10(rand_exe_prng_150_io_out_10),
    .io_out_11(rand_exe_prng_150_io_out_11),
    .io_out_12(rand_exe_prng_150_io_out_12),
    .io_out_13(rand_exe_prng_150_io_out_13),
    .io_out_14(rand_exe_prng_150_io_out_14),
    .io_out_15(rand_exe_prng_150_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_151 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_151_clock),
    .reset(rand_exe_prng_151_reset),
    .io_out_0(rand_exe_prng_151_io_out_0),
    .io_out_1(rand_exe_prng_151_io_out_1),
    .io_out_2(rand_exe_prng_151_io_out_2),
    .io_out_3(rand_exe_prng_151_io_out_3),
    .io_out_4(rand_exe_prng_151_io_out_4),
    .io_out_5(rand_exe_prng_151_io_out_5),
    .io_out_6(rand_exe_prng_151_io_out_6),
    .io_out_7(rand_exe_prng_151_io_out_7),
    .io_out_8(rand_exe_prng_151_io_out_8),
    .io_out_9(rand_exe_prng_151_io_out_9),
    .io_out_10(rand_exe_prng_151_io_out_10),
    .io_out_11(rand_exe_prng_151_io_out_11),
    .io_out_12(rand_exe_prng_151_io_out_12),
    .io_out_13(rand_exe_prng_151_io_out_13),
    .io_out_14(rand_exe_prng_151_io_out_14),
    .io_out_15(rand_exe_prng_151_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_152 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_152_clock),
    .reset(rand_exe_prng_152_reset),
    .io_out_0(rand_exe_prng_152_io_out_0),
    .io_out_1(rand_exe_prng_152_io_out_1),
    .io_out_2(rand_exe_prng_152_io_out_2),
    .io_out_3(rand_exe_prng_152_io_out_3),
    .io_out_4(rand_exe_prng_152_io_out_4),
    .io_out_5(rand_exe_prng_152_io_out_5),
    .io_out_6(rand_exe_prng_152_io_out_6),
    .io_out_7(rand_exe_prng_152_io_out_7),
    .io_out_8(rand_exe_prng_152_io_out_8),
    .io_out_9(rand_exe_prng_152_io_out_9),
    .io_out_10(rand_exe_prng_152_io_out_10),
    .io_out_11(rand_exe_prng_152_io_out_11),
    .io_out_12(rand_exe_prng_152_io_out_12),
    .io_out_13(rand_exe_prng_152_io_out_13),
    .io_out_14(rand_exe_prng_152_io_out_14),
    .io_out_15(rand_exe_prng_152_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_153 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_153_clock),
    .reset(rand_exe_prng_153_reset),
    .io_out_0(rand_exe_prng_153_io_out_0),
    .io_out_1(rand_exe_prng_153_io_out_1),
    .io_out_2(rand_exe_prng_153_io_out_2),
    .io_out_3(rand_exe_prng_153_io_out_3),
    .io_out_4(rand_exe_prng_153_io_out_4),
    .io_out_5(rand_exe_prng_153_io_out_5),
    .io_out_6(rand_exe_prng_153_io_out_6),
    .io_out_7(rand_exe_prng_153_io_out_7),
    .io_out_8(rand_exe_prng_153_io_out_8),
    .io_out_9(rand_exe_prng_153_io_out_9),
    .io_out_10(rand_exe_prng_153_io_out_10),
    .io_out_11(rand_exe_prng_153_io_out_11),
    .io_out_12(rand_exe_prng_153_io_out_12),
    .io_out_13(rand_exe_prng_153_io_out_13),
    .io_out_14(rand_exe_prng_153_io_out_14),
    .io_out_15(rand_exe_prng_153_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_154 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_154_clock),
    .reset(rand_exe_prng_154_reset),
    .io_out_0(rand_exe_prng_154_io_out_0),
    .io_out_1(rand_exe_prng_154_io_out_1),
    .io_out_2(rand_exe_prng_154_io_out_2),
    .io_out_3(rand_exe_prng_154_io_out_3),
    .io_out_4(rand_exe_prng_154_io_out_4),
    .io_out_5(rand_exe_prng_154_io_out_5),
    .io_out_6(rand_exe_prng_154_io_out_6),
    .io_out_7(rand_exe_prng_154_io_out_7),
    .io_out_8(rand_exe_prng_154_io_out_8),
    .io_out_9(rand_exe_prng_154_io_out_9),
    .io_out_10(rand_exe_prng_154_io_out_10),
    .io_out_11(rand_exe_prng_154_io_out_11),
    .io_out_12(rand_exe_prng_154_io_out_12),
    .io_out_13(rand_exe_prng_154_io_out_13),
    .io_out_14(rand_exe_prng_154_io_out_14),
    .io_out_15(rand_exe_prng_154_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_155 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_155_clock),
    .reset(rand_exe_prng_155_reset),
    .io_out_0(rand_exe_prng_155_io_out_0),
    .io_out_1(rand_exe_prng_155_io_out_1),
    .io_out_2(rand_exe_prng_155_io_out_2),
    .io_out_3(rand_exe_prng_155_io_out_3),
    .io_out_4(rand_exe_prng_155_io_out_4),
    .io_out_5(rand_exe_prng_155_io_out_5),
    .io_out_6(rand_exe_prng_155_io_out_6),
    .io_out_7(rand_exe_prng_155_io_out_7),
    .io_out_8(rand_exe_prng_155_io_out_8),
    .io_out_9(rand_exe_prng_155_io_out_9),
    .io_out_10(rand_exe_prng_155_io_out_10),
    .io_out_11(rand_exe_prng_155_io_out_11),
    .io_out_12(rand_exe_prng_155_io_out_12),
    .io_out_13(rand_exe_prng_155_io_out_13),
    .io_out_14(rand_exe_prng_155_io_out_14),
    .io_out_15(rand_exe_prng_155_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_156 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_156_clock),
    .reset(rand_exe_prng_156_reset),
    .io_out_0(rand_exe_prng_156_io_out_0),
    .io_out_1(rand_exe_prng_156_io_out_1),
    .io_out_2(rand_exe_prng_156_io_out_2),
    .io_out_3(rand_exe_prng_156_io_out_3),
    .io_out_4(rand_exe_prng_156_io_out_4),
    .io_out_5(rand_exe_prng_156_io_out_5),
    .io_out_6(rand_exe_prng_156_io_out_6),
    .io_out_7(rand_exe_prng_156_io_out_7),
    .io_out_8(rand_exe_prng_156_io_out_8),
    .io_out_9(rand_exe_prng_156_io_out_9),
    .io_out_10(rand_exe_prng_156_io_out_10),
    .io_out_11(rand_exe_prng_156_io_out_11),
    .io_out_12(rand_exe_prng_156_io_out_12),
    .io_out_13(rand_exe_prng_156_io_out_13),
    .io_out_14(rand_exe_prng_156_io_out_14),
    .io_out_15(rand_exe_prng_156_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_157 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_157_clock),
    .reset(rand_exe_prng_157_reset),
    .io_out_0(rand_exe_prng_157_io_out_0),
    .io_out_1(rand_exe_prng_157_io_out_1),
    .io_out_2(rand_exe_prng_157_io_out_2),
    .io_out_3(rand_exe_prng_157_io_out_3),
    .io_out_4(rand_exe_prng_157_io_out_4),
    .io_out_5(rand_exe_prng_157_io_out_5),
    .io_out_6(rand_exe_prng_157_io_out_6),
    .io_out_7(rand_exe_prng_157_io_out_7),
    .io_out_8(rand_exe_prng_157_io_out_8),
    .io_out_9(rand_exe_prng_157_io_out_9),
    .io_out_10(rand_exe_prng_157_io_out_10),
    .io_out_11(rand_exe_prng_157_io_out_11),
    .io_out_12(rand_exe_prng_157_io_out_12),
    .io_out_13(rand_exe_prng_157_io_out_13),
    .io_out_14(rand_exe_prng_157_io_out_14),
    .io_out_15(rand_exe_prng_157_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_158 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_158_clock),
    .reset(rand_exe_prng_158_reset),
    .io_out_0(rand_exe_prng_158_io_out_0),
    .io_out_1(rand_exe_prng_158_io_out_1),
    .io_out_2(rand_exe_prng_158_io_out_2),
    .io_out_3(rand_exe_prng_158_io_out_3),
    .io_out_4(rand_exe_prng_158_io_out_4),
    .io_out_5(rand_exe_prng_158_io_out_5),
    .io_out_6(rand_exe_prng_158_io_out_6),
    .io_out_7(rand_exe_prng_158_io_out_7),
    .io_out_8(rand_exe_prng_158_io_out_8),
    .io_out_9(rand_exe_prng_158_io_out_9),
    .io_out_10(rand_exe_prng_158_io_out_10),
    .io_out_11(rand_exe_prng_158_io_out_11),
    .io_out_12(rand_exe_prng_158_io_out_12),
    .io_out_13(rand_exe_prng_158_io_out_13),
    .io_out_14(rand_exe_prng_158_io_out_14),
    .io_out_15(rand_exe_prng_158_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_159 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_159_clock),
    .reset(rand_exe_prng_159_reset),
    .io_out_0(rand_exe_prng_159_io_out_0),
    .io_out_1(rand_exe_prng_159_io_out_1),
    .io_out_2(rand_exe_prng_159_io_out_2),
    .io_out_3(rand_exe_prng_159_io_out_3),
    .io_out_4(rand_exe_prng_159_io_out_4),
    .io_out_5(rand_exe_prng_159_io_out_5),
    .io_out_6(rand_exe_prng_159_io_out_6),
    .io_out_7(rand_exe_prng_159_io_out_7),
    .io_out_8(rand_exe_prng_159_io_out_8),
    .io_out_9(rand_exe_prng_159_io_out_9),
    .io_out_10(rand_exe_prng_159_io_out_10),
    .io_out_11(rand_exe_prng_159_io_out_11),
    .io_out_12(rand_exe_prng_159_io_out_12),
    .io_out_13(rand_exe_prng_159_io_out_13),
    .io_out_14(rand_exe_prng_159_io_out_14),
    .io_out_15(rand_exe_prng_159_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_160 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_160_clock),
    .reset(rand_exe_prng_160_reset),
    .io_out_0(rand_exe_prng_160_io_out_0),
    .io_out_1(rand_exe_prng_160_io_out_1),
    .io_out_2(rand_exe_prng_160_io_out_2),
    .io_out_3(rand_exe_prng_160_io_out_3),
    .io_out_4(rand_exe_prng_160_io_out_4),
    .io_out_5(rand_exe_prng_160_io_out_5),
    .io_out_6(rand_exe_prng_160_io_out_6),
    .io_out_7(rand_exe_prng_160_io_out_7),
    .io_out_8(rand_exe_prng_160_io_out_8),
    .io_out_9(rand_exe_prng_160_io_out_9),
    .io_out_10(rand_exe_prng_160_io_out_10),
    .io_out_11(rand_exe_prng_160_io_out_11),
    .io_out_12(rand_exe_prng_160_io_out_12),
    .io_out_13(rand_exe_prng_160_io_out_13),
    .io_out_14(rand_exe_prng_160_io_out_14),
    .io_out_15(rand_exe_prng_160_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_161 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_161_clock),
    .reset(rand_exe_prng_161_reset),
    .io_out_0(rand_exe_prng_161_io_out_0),
    .io_out_1(rand_exe_prng_161_io_out_1),
    .io_out_2(rand_exe_prng_161_io_out_2),
    .io_out_3(rand_exe_prng_161_io_out_3),
    .io_out_4(rand_exe_prng_161_io_out_4),
    .io_out_5(rand_exe_prng_161_io_out_5),
    .io_out_6(rand_exe_prng_161_io_out_6),
    .io_out_7(rand_exe_prng_161_io_out_7),
    .io_out_8(rand_exe_prng_161_io_out_8),
    .io_out_9(rand_exe_prng_161_io_out_9),
    .io_out_10(rand_exe_prng_161_io_out_10),
    .io_out_11(rand_exe_prng_161_io_out_11),
    .io_out_12(rand_exe_prng_161_io_out_12),
    .io_out_13(rand_exe_prng_161_io_out_13),
    .io_out_14(rand_exe_prng_161_io_out_14),
    .io_out_15(rand_exe_prng_161_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_162 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_162_clock),
    .reset(rand_exe_prng_162_reset),
    .io_out_0(rand_exe_prng_162_io_out_0),
    .io_out_1(rand_exe_prng_162_io_out_1),
    .io_out_2(rand_exe_prng_162_io_out_2),
    .io_out_3(rand_exe_prng_162_io_out_3),
    .io_out_4(rand_exe_prng_162_io_out_4),
    .io_out_5(rand_exe_prng_162_io_out_5),
    .io_out_6(rand_exe_prng_162_io_out_6),
    .io_out_7(rand_exe_prng_162_io_out_7),
    .io_out_8(rand_exe_prng_162_io_out_8),
    .io_out_9(rand_exe_prng_162_io_out_9),
    .io_out_10(rand_exe_prng_162_io_out_10),
    .io_out_11(rand_exe_prng_162_io_out_11),
    .io_out_12(rand_exe_prng_162_io_out_12),
    .io_out_13(rand_exe_prng_162_io_out_13),
    .io_out_14(rand_exe_prng_162_io_out_14),
    .io_out_15(rand_exe_prng_162_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_163 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_163_clock),
    .reset(rand_exe_prng_163_reset),
    .io_out_0(rand_exe_prng_163_io_out_0),
    .io_out_1(rand_exe_prng_163_io_out_1),
    .io_out_2(rand_exe_prng_163_io_out_2),
    .io_out_3(rand_exe_prng_163_io_out_3),
    .io_out_4(rand_exe_prng_163_io_out_4),
    .io_out_5(rand_exe_prng_163_io_out_5),
    .io_out_6(rand_exe_prng_163_io_out_6),
    .io_out_7(rand_exe_prng_163_io_out_7),
    .io_out_8(rand_exe_prng_163_io_out_8),
    .io_out_9(rand_exe_prng_163_io_out_9),
    .io_out_10(rand_exe_prng_163_io_out_10),
    .io_out_11(rand_exe_prng_163_io_out_11),
    .io_out_12(rand_exe_prng_163_io_out_12),
    .io_out_13(rand_exe_prng_163_io_out_13),
    .io_out_14(rand_exe_prng_163_io_out_14),
    .io_out_15(rand_exe_prng_163_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_164 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_164_clock),
    .reset(rand_exe_prng_164_reset),
    .io_out_0(rand_exe_prng_164_io_out_0),
    .io_out_1(rand_exe_prng_164_io_out_1),
    .io_out_2(rand_exe_prng_164_io_out_2),
    .io_out_3(rand_exe_prng_164_io_out_3),
    .io_out_4(rand_exe_prng_164_io_out_4),
    .io_out_5(rand_exe_prng_164_io_out_5),
    .io_out_6(rand_exe_prng_164_io_out_6),
    .io_out_7(rand_exe_prng_164_io_out_7),
    .io_out_8(rand_exe_prng_164_io_out_8),
    .io_out_9(rand_exe_prng_164_io_out_9),
    .io_out_10(rand_exe_prng_164_io_out_10),
    .io_out_11(rand_exe_prng_164_io_out_11),
    .io_out_12(rand_exe_prng_164_io_out_12),
    .io_out_13(rand_exe_prng_164_io_out_13),
    .io_out_14(rand_exe_prng_164_io_out_14),
    .io_out_15(rand_exe_prng_164_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_165 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_165_clock),
    .reset(rand_exe_prng_165_reset),
    .io_out_0(rand_exe_prng_165_io_out_0),
    .io_out_1(rand_exe_prng_165_io_out_1),
    .io_out_2(rand_exe_prng_165_io_out_2),
    .io_out_3(rand_exe_prng_165_io_out_3),
    .io_out_4(rand_exe_prng_165_io_out_4),
    .io_out_5(rand_exe_prng_165_io_out_5),
    .io_out_6(rand_exe_prng_165_io_out_6),
    .io_out_7(rand_exe_prng_165_io_out_7),
    .io_out_8(rand_exe_prng_165_io_out_8),
    .io_out_9(rand_exe_prng_165_io_out_9),
    .io_out_10(rand_exe_prng_165_io_out_10),
    .io_out_11(rand_exe_prng_165_io_out_11),
    .io_out_12(rand_exe_prng_165_io_out_12),
    .io_out_13(rand_exe_prng_165_io_out_13),
    .io_out_14(rand_exe_prng_165_io_out_14),
    .io_out_15(rand_exe_prng_165_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_166 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_166_clock),
    .reset(rand_exe_prng_166_reset),
    .io_out_0(rand_exe_prng_166_io_out_0),
    .io_out_1(rand_exe_prng_166_io_out_1),
    .io_out_2(rand_exe_prng_166_io_out_2),
    .io_out_3(rand_exe_prng_166_io_out_3),
    .io_out_4(rand_exe_prng_166_io_out_4),
    .io_out_5(rand_exe_prng_166_io_out_5),
    .io_out_6(rand_exe_prng_166_io_out_6),
    .io_out_7(rand_exe_prng_166_io_out_7),
    .io_out_8(rand_exe_prng_166_io_out_8),
    .io_out_9(rand_exe_prng_166_io_out_9),
    .io_out_10(rand_exe_prng_166_io_out_10),
    .io_out_11(rand_exe_prng_166_io_out_11),
    .io_out_12(rand_exe_prng_166_io_out_12),
    .io_out_13(rand_exe_prng_166_io_out_13),
    .io_out_14(rand_exe_prng_166_io_out_14),
    .io_out_15(rand_exe_prng_166_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_167 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_167_clock),
    .reset(rand_exe_prng_167_reset),
    .io_out_0(rand_exe_prng_167_io_out_0),
    .io_out_1(rand_exe_prng_167_io_out_1),
    .io_out_2(rand_exe_prng_167_io_out_2),
    .io_out_3(rand_exe_prng_167_io_out_3),
    .io_out_4(rand_exe_prng_167_io_out_4),
    .io_out_5(rand_exe_prng_167_io_out_5),
    .io_out_6(rand_exe_prng_167_io_out_6),
    .io_out_7(rand_exe_prng_167_io_out_7),
    .io_out_8(rand_exe_prng_167_io_out_8),
    .io_out_9(rand_exe_prng_167_io_out_9),
    .io_out_10(rand_exe_prng_167_io_out_10),
    .io_out_11(rand_exe_prng_167_io_out_11),
    .io_out_12(rand_exe_prng_167_io_out_12),
    .io_out_13(rand_exe_prng_167_io_out_13),
    .io_out_14(rand_exe_prng_167_io_out_14),
    .io_out_15(rand_exe_prng_167_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_168 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_168_clock),
    .reset(rand_exe_prng_168_reset),
    .io_out_0(rand_exe_prng_168_io_out_0),
    .io_out_1(rand_exe_prng_168_io_out_1),
    .io_out_2(rand_exe_prng_168_io_out_2),
    .io_out_3(rand_exe_prng_168_io_out_3),
    .io_out_4(rand_exe_prng_168_io_out_4),
    .io_out_5(rand_exe_prng_168_io_out_5),
    .io_out_6(rand_exe_prng_168_io_out_6),
    .io_out_7(rand_exe_prng_168_io_out_7),
    .io_out_8(rand_exe_prng_168_io_out_8),
    .io_out_9(rand_exe_prng_168_io_out_9),
    .io_out_10(rand_exe_prng_168_io_out_10),
    .io_out_11(rand_exe_prng_168_io_out_11),
    .io_out_12(rand_exe_prng_168_io_out_12),
    .io_out_13(rand_exe_prng_168_io_out_13),
    .io_out_14(rand_exe_prng_168_io_out_14),
    .io_out_15(rand_exe_prng_168_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_169 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_169_clock),
    .reset(rand_exe_prng_169_reset),
    .io_out_0(rand_exe_prng_169_io_out_0),
    .io_out_1(rand_exe_prng_169_io_out_1),
    .io_out_2(rand_exe_prng_169_io_out_2),
    .io_out_3(rand_exe_prng_169_io_out_3),
    .io_out_4(rand_exe_prng_169_io_out_4),
    .io_out_5(rand_exe_prng_169_io_out_5),
    .io_out_6(rand_exe_prng_169_io_out_6),
    .io_out_7(rand_exe_prng_169_io_out_7),
    .io_out_8(rand_exe_prng_169_io_out_8),
    .io_out_9(rand_exe_prng_169_io_out_9),
    .io_out_10(rand_exe_prng_169_io_out_10),
    .io_out_11(rand_exe_prng_169_io_out_11),
    .io_out_12(rand_exe_prng_169_io_out_12),
    .io_out_13(rand_exe_prng_169_io_out_13),
    .io_out_14(rand_exe_prng_169_io_out_14),
    .io_out_15(rand_exe_prng_169_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_170 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_170_clock),
    .reset(rand_exe_prng_170_reset),
    .io_out_0(rand_exe_prng_170_io_out_0),
    .io_out_1(rand_exe_prng_170_io_out_1),
    .io_out_2(rand_exe_prng_170_io_out_2),
    .io_out_3(rand_exe_prng_170_io_out_3),
    .io_out_4(rand_exe_prng_170_io_out_4),
    .io_out_5(rand_exe_prng_170_io_out_5),
    .io_out_6(rand_exe_prng_170_io_out_6),
    .io_out_7(rand_exe_prng_170_io_out_7),
    .io_out_8(rand_exe_prng_170_io_out_8),
    .io_out_9(rand_exe_prng_170_io_out_9),
    .io_out_10(rand_exe_prng_170_io_out_10),
    .io_out_11(rand_exe_prng_170_io_out_11),
    .io_out_12(rand_exe_prng_170_io_out_12),
    .io_out_13(rand_exe_prng_170_io_out_13),
    .io_out_14(rand_exe_prng_170_io_out_14),
    .io_out_15(rand_exe_prng_170_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_171 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_171_clock),
    .reset(rand_exe_prng_171_reset),
    .io_out_0(rand_exe_prng_171_io_out_0),
    .io_out_1(rand_exe_prng_171_io_out_1),
    .io_out_2(rand_exe_prng_171_io_out_2),
    .io_out_3(rand_exe_prng_171_io_out_3),
    .io_out_4(rand_exe_prng_171_io_out_4),
    .io_out_5(rand_exe_prng_171_io_out_5),
    .io_out_6(rand_exe_prng_171_io_out_6),
    .io_out_7(rand_exe_prng_171_io_out_7),
    .io_out_8(rand_exe_prng_171_io_out_8),
    .io_out_9(rand_exe_prng_171_io_out_9),
    .io_out_10(rand_exe_prng_171_io_out_10),
    .io_out_11(rand_exe_prng_171_io_out_11),
    .io_out_12(rand_exe_prng_171_io_out_12),
    .io_out_13(rand_exe_prng_171_io_out_13),
    .io_out_14(rand_exe_prng_171_io_out_14),
    .io_out_15(rand_exe_prng_171_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_172 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_172_clock),
    .reset(rand_exe_prng_172_reset),
    .io_out_0(rand_exe_prng_172_io_out_0),
    .io_out_1(rand_exe_prng_172_io_out_1),
    .io_out_2(rand_exe_prng_172_io_out_2),
    .io_out_3(rand_exe_prng_172_io_out_3),
    .io_out_4(rand_exe_prng_172_io_out_4),
    .io_out_5(rand_exe_prng_172_io_out_5),
    .io_out_6(rand_exe_prng_172_io_out_6),
    .io_out_7(rand_exe_prng_172_io_out_7),
    .io_out_8(rand_exe_prng_172_io_out_8),
    .io_out_9(rand_exe_prng_172_io_out_9),
    .io_out_10(rand_exe_prng_172_io_out_10),
    .io_out_11(rand_exe_prng_172_io_out_11),
    .io_out_12(rand_exe_prng_172_io_out_12),
    .io_out_13(rand_exe_prng_172_io_out_13),
    .io_out_14(rand_exe_prng_172_io_out_14),
    .io_out_15(rand_exe_prng_172_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_173 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_173_clock),
    .reset(rand_exe_prng_173_reset),
    .io_out_0(rand_exe_prng_173_io_out_0),
    .io_out_1(rand_exe_prng_173_io_out_1),
    .io_out_2(rand_exe_prng_173_io_out_2),
    .io_out_3(rand_exe_prng_173_io_out_3),
    .io_out_4(rand_exe_prng_173_io_out_4),
    .io_out_5(rand_exe_prng_173_io_out_5),
    .io_out_6(rand_exe_prng_173_io_out_6),
    .io_out_7(rand_exe_prng_173_io_out_7),
    .io_out_8(rand_exe_prng_173_io_out_8),
    .io_out_9(rand_exe_prng_173_io_out_9),
    .io_out_10(rand_exe_prng_173_io_out_10),
    .io_out_11(rand_exe_prng_173_io_out_11),
    .io_out_12(rand_exe_prng_173_io_out_12),
    .io_out_13(rand_exe_prng_173_io_out_13),
    .io_out_14(rand_exe_prng_173_io_out_14),
    .io_out_15(rand_exe_prng_173_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_174 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_174_clock),
    .reset(rand_exe_prng_174_reset),
    .io_out_0(rand_exe_prng_174_io_out_0),
    .io_out_1(rand_exe_prng_174_io_out_1),
    .io_out_2(rand_exe_prng_174_io_out_2),
    .io_out_3(rand_exe_prng_174_io_out_3),
    .io_out_4(rand_exe_prng_174_io_out_4),
    .io_out_5(rand_exe_prng_174_io_out_5),
    .io_out_6(rand_exe_prng_174_io_out_6),
    .io_out_7(rand_exe_prng_174_io_out_7),
    .io_out_8(rand_exe_prng_174_io_out_8),
    .io_out_9(rand_exe_prng_174_io_out_9),
    .io_out_10(rand_exe_prng_174_io_out_10),
    .io_out_11(rand_exe_prng_174_io_out_11),
    .io_out_12(rand_exe_prng_174_io_out_12),
    .io_out_13(rand_exe_prng_174_io_out_13),
    .io_out_14(rand_exe_prng_174_io_out_14),
    .io_out_15(rand_exe_prng_174_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_175 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_175_clock),
    .reset(rand_exe_prng_175_reset),
    .io_out_0(rand_exe_prng_175_io_out_0),
    .io_out_1(rand_exe_prng_175_io_out_1),
    .io_out_2(rand_exe_prng_175_io_out_2),
    .io_out_3(rand_exe_prng_175_io_out_3),
    .io_out_4(rand_exe_prng_175_io_out_4),
    .io_out_5(rand_exe_prng_175_io_out_5),
    .io_out_6(rand_exe_prng_175_io_out_6),
    .io_out_7(rand_exe_prng_175_io_out_7),
    .io_out_8(rand_exe_prng_175_io_out_8),
    .io_out_9(rand_exe_prng_175_io_out_9),
    .io_out_10(rand_exe_prng_175_io_out_10),
    .io_out_11(rand_exe_prng_175_io_out_11),
    .io_out_12(rand_exe_prng_175_io_out_12),
    .io_out_13(rand_exe_prng_175_io_out_13),
    .io_out_14(rand_exe_prng_175_io_out_14),
    .io_out_15(rand_exe_prng_175_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_176 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_176_clock),
    .reset(rand_exe_prng_176_reset),
    .io_out_0(rand_exe_prng_176_io_out_0),
    .io_out_1(rand_exe_prng_176_io_out_1),
    .io_out_2(rand_exe_prng_176_io_out_2),
    .io_out_3(rand_exe_prng_176_io_out_3),
    .io_out_4(rand_exe_prng_176_io_out_4),
    .io_out_5(rand_exe_prng_176_io_out_5),
    .io_out_6(rand_exe_prng_176_io_out_6),
    .io_out_7(rand_exe_prng_176_io_out_7),
    .io_out_8(rand_exe_prng_176_io_out_8),
    .io_out_9(rand_exe_prng_176_io_out_9),
    .io_out_10(rand_exe_prng_176_io_out_10),
    .io_out_11(rand_exe_prng_176_io_out_11),
    .io_out_12(rand_exe_prng_176_io_out_12),
    .io_out_13(rand_exe_prng_176_io_out_13),
    .io_out_14(rand_exe_prng_176_io_out_14),
    .io_out_15(rand_exe_prng_176_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_177 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_177_clock),
    .reset(rand_exe_prng_177_reset),
    .io_out_0(rand_exe_prng_177_io_out_0),
    .io_out_1(rand_exe_prng_177_io_out_1),
    .io_out_2(rand_exe_prng_177_io_out_2),
    .io_out_3(rand_exe_prng_177_io_out_3),
    .io_out_4(rand_exe_prng_177_io_out_4),
    .io_out_5(rand_exe_prng_177_io_out_5),
    .io_out_6(rand_exe_prng_177_io_out_6),
    .io_out_7(rand_exe_prng_177_io_out_7),
    .io_out_8(rand_exe_prng_177_io_out_8),
    .io_out_9(rand_exe_prng_177_io_out_9),
    .io_out_10(rand_exe_prng_177_io_out_10),
    .io_out_11(rand_exe_prng_177_io_out_11),
    .io_out_12(rand_exe_prng_177_io_out_12),
    .io_out_13(rand_exe_prng_177_io_out_13),
    .io_out_14(rand_exe_prng_177_io_out_14),
    .io_out_15(rand_exe_prng_177_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_178 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_178_clock),
    .reset(rand_exe_prng_178_reset),
    .io_out_0(rand_exe_prng_178_io_out_0),
    .io_out_1(rand_exe_prng_178_io_out_1),
    .io_out_2(rand_exe_prng_178_io_out_2),
    .io_out_3(rand_exe_prng_178_io_out_3),
    .io_out_4(rand_exe_prng_178_io_out_4),
    .io_out_5(rand_exe_prng_178_io_out_5),
    .io_out_6(rand_exe_prng_178_io_out_6),
    .io_out_7(rand_exe_prng_178_io_out_7),
    .io_out_8(rand_exe_prng_178_io_out_8),
    .io_out_9(rand_exe_prng_178_io_out_9),
    .io_out_10(rand_exe_prng_178_io_out_10),
    .io_out_11(rand_exe_prng_178_io_out_11),
    .io_out_12(rand_exe_prng_178_io_out_12),
    .io_out_13(rand_exe_prng_178_io_out_13),
    .io_out_14(rand_exe_prng_178_io_out_14),
    .io_out_15(rand_exe_prng_178_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_179 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_179_clock),
    .reset(rand_exe_prng_179_reset),
    .io_out_0(rand_exe_prng_179_io_out_0),
    .io_out_1(rand_exe_prng_179_io_out_1),
    .io_out_2(rand_exe_prng_179_io_out_2),
    .io_out_3(rand_exe_prng_179_io_out_3),
    .io_out_4(rand_exe_prng_179_io_out_4),
    .io_out_5(rand_exe_prng_179_io_out_5),
    .io_out_6(rand_exe_prng_179_io_out_6),
    .io_out_7(rand_exe_prng_179_io_out_7),
    .io_out_8(rand_exe_prng_179_io_out_8),
    .io_out_9(rand_exe_prng_179_io_out_9),
    .io_out_10(rand_exe_prng_179_io_out_10),
    .io_out_11(rand_exe_prng_179_io_out_11),
    .io_out_12(rand_exe_prng_179_io_out_12),
    .io_out_13(rand_exe_prng_179_io_out_13),
    .io_out_14(rand_exe_prng_179_io_out_14),
    .io_out_15(rand_exe_prng_179_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_180 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_180_clock),
    .reset(rand_exe_prng_180_reset),
    .io_out_0(rand_exe_prng_180_io_out_0),
    .io_out_1(rand_exe_prng_180_io_out_1),
    .io_out_2(rand_exe_prng_180_io_out_2),
    .io_out_3(rand_exe_prng_180_io_out_3),
    .io_out_4(rand_exe_prng_180_io_out_4),
    .io_out_5(rand_exe_prng_180_io_out_5),
    .io_out_6(rand_exe_prng_180_io_out_6),
    .io_out_7(rand_exe_prng_180_io_out_7),
    .io_out_8(rand_exe_prng_180_io_out_8),
    .io_out_9(rand_exe_prng_180_io_out_9),
    .io_out_10(rand_exe_prng_180_io_out_10),
    .io_out_11(rand_exe_prng_180_io_out_11),
    .io_out_12(rand_exe_prng_180_io_out_12),
    .io_out_13(rand_exe_prng_180_io_out_13),
    .io_out_14(rand_exe_prng_180_io_out_14),
    .io_out_15(rand_exe_prng_180_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_181 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_181_clock),
    .reset(rand_exe_prng_181_reset),
    .io_out_0(rand_exe_prng_181_io_out_0),
    .io_out_1(rand_exe_prng_181_io_out_1),
    .io_out_2(rand_exe_prng_181_io_out_2),
    .io_out_3(rand_exe_prng_181_io_out_3),
    .io_out_4(rand_exe_prng_181_io_out_4),
    .io_out_5(rand_exe_prng_181_io_out_5),
    .io_out_6(rand_exe_prng_181_io_out_6),
    .io_out_7(rand_exe_prng_181_io_out_7),
    .io_out_8(rand_exe_prng_181_io_out_8),
    .io_out_9(rand_exe_prng_181_io_out_9),
    .io_out_10(rand_exe_prng_181_io_out_10),
    .io_out_11(rand_exe_prng_181_io_out_11),
    .io_out_12(rand_exe_prng_181_io_out_12),
    .io_out_13(rand_exe_prng_181_io_out_13),
    .io_out_14(rand_exe_prng_181_io_out_14),
    .io_out_15(rand_exe_prng_181_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_182 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_182_clock),
    .reset(rand_exe_prng_182_reset),
    .io_out_0(rand_exe_prng_182_io_out_0),
    .io_out_1(rand_exe_prng_182_io_out_1),
    .io_out_2(rand_exe_prng_182_io_out_2),
    .io_out_3(rand_exe_prng_182_io_out_3),
    .io_out_4(rand_exe_prng_182_io_out_4),
    .io_out_5(rand_exe_prng_182_io_out_5),
    .io_out_6(rand_exe_prng_182_io_out_6),
    .io_out_7(rand_exe_prng_182_io_out_7),
    .io_out_8(rand_exe_prng_182_io_out_8),
    .io_out_9(rand_exe_prng_182_io_out_9),
    .io_out_10(rand_exe_prng_182_io_out_10),
    .io_out_11(rand_exe_prng_182_io_out_11),
    .io_out_12(rand_exe_prng_182_io_out_12),
    .io_out_13(rand_exe_prng_182_io_out_13),
    .io_out_14(rand_exe_prng_182_io_out_14),
    .io_out_15(rand_exe_prng_182_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_183 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_183_clock),
    .reset(rand_exe_prng_183_reset),
    .io_out_0(rand_exe_prng_183_io_out_0),
    .io_out_1(rand_exe_prng_183_io_out_1),
    .io_out_2(rand_exe_prng_183_io_out_2),
    .io_out_3(rand_exe_prng_183_io_out_3),
    .io_out_4(rand_exe_prng_183_io_out_4),
    .io_out_5(rand_exe_prng_183_io_out_5),
    .io_out_6(rand_exe_prng_183_io_out_6),
    .io_out_7(rand_exe_prng_183_io_out_7),
    .io_out_8(rand_exe_prng_183_io_out_8),
    .io_out_9(rand_exe_prng_183_io_out_9),
    .io_out_10(rand_exe_prng_183_io_out_10),
    .io_out_11(rand_exe_prng_183_io_out_11),
    .io_out_12(rand_exe_prng_183_io_out_12),
    .io_out_13(rand_exe_prng_183_io_out_13),
    .io_out_14(rand_exe_prng_183_io_out_14),
    .io_out_15(rand_exe_prng_183_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_184 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_184_clock),
    .reset(rand_exe_prng_184_reset),
    .io_out_0(rand_exe_prng_184_io_out_0),
    .io_out_1(rand_exe_prng_184_io_out_1),
    .io_out_2(rand_exe_prng_184_io_out_2),
    .io_out_3(rand_exe_prng_184_io_out_3),
    .io_out_4(rand_exe_prng_184_io_out_4),
    .io_out_5(rand_exe_prng_184_io_out_5),
    .io_out_6(rand_exe_prng_184_io_out_6),
    .io_out_7(rand_exe_prng_184_io_out_7),
    .io_out_8(rand_exe_prng_184_io_out_8),
    .io_out_9(rand_exe_prng_184_io_out_9),
    .io_out_10(rand_exe_prng_184_io_out_10),
    .io_out_11(rand_exe_prng_184_io_out_11),
    .io_out_12(rand_exe_prng_184_io_out_12),
    .io_out_13(rand_exe_prng_184_io_out_13),
    .io_out_14(rand_exe_prng_184_io_out_14),
    .io_out_15(rand_exe_prng_184_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_185 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_185_clock),
    .reset(rand_exe_prng_185_reset),
    .io_out_0(rand_exe_prng_185_io_out_0),
    .io_out_1(rand_exe_prng_185_io_out_1),
    .io_out_2(rand_exe_prng_185_io_out_2),
    .io_out_3(rand_exe_prng_185_io_out_3),
    .io_out_4(rand_exe_prng_185_io_out_4),
    .io_out_5(rand_exe_prng_185_io_out_5),
    .io_out_6(rand_exe_prng_185_io_out_6),
    .io_out_7(rand_exe_prng_185_io_out_7),
    .io_out_8(rand_exe_prng_185_io_out_8),
    .io_out_9(rand_exe_prng_185_io_out_9),
    .io_out_10(rand_exe_prng_185_io_out_10),
    .io_out_11(rand_exe_prng_185_io_out_11),
    .io_out_12(rand_exe_prng_185_io_out_12),
    .io_out_13(rand_exe_prng_185_io_out_13),
    .io_out_14(rand_exe_prng_185_io_out_14),
    .io_out_15(rand_exe_prng_185_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_186 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_186_clock),
    .reset(rand_exe_prng_186_reset),
    .io_out_0(rand_exe_prng_186_io_out_0),
    .io_out_1(rand_exe_prng_186_io_out_1),
    .io_out_2(rand_exe_prng_186_io_out_2),
    .io_out_3(rand_exe_prng_186_io_out_3),
    .io_out_4(rand_exe_prng_186_io_out_4),
    .io_out_5(rand_exe_prng_186_io_out_5),
    .io_out_6(rand_exe_prng_186_io_out_6),
    .io_out_7(rand_exe_prng_186_io_out_7),
    .io_out_8(rand_exe_prng_186_io_out_8),
    .io_out_9(rand_exe_prng_186_io_out_9),
    .io_out_10(rand_exe_prng_186_io_out_10),
    .io_out_11(rand_exe_prng_186_io_out_11),
    .io_out_12(rand_exe_prng_186_io_out_12),
    .io_out_13(rand_exe_prng_186_io_out_13),
    .io_out_14(rand_exe_prng_186_io_out_14),
    .io_out_15(rand_exe_prng_186_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_187 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_187_clock),
    .reset(rand_exe_prng_187_reset),
    .io_out_0(rand_exe_prng_187_io_out_0),
    .io_out_1(rand_exe_prng_187_io_out_1),
    .io_out_2(rand_exe_prng_187_io_out_2),
    .io_out_3(rand_exe_prng_187_io_out_3),
    .io_out_4(rand_exe_prng_187_io_out_4),
    .io_out_5(rand_exe_prng_187_io_out_5),
    .io_out_6(rand_exe_prng_187_io_out_6),
    .io_out_7(rand_exe_prng_187_io_out_7),
    .io_out_8(rand_exe_prng_187_io_out_8),
    .io_out_9(rand_exe_prng_187_io_out_9),
    .io_out_10(rand_exe_prng_187_io_out_10),
    .io_out_11(rand_exe_prng_187_io_out_11),
    .io_out_12(rand_exe_prng_187_io_out_12),
    .io_out_13(rand_exe_prng_187_io_out_13),
    .io_out_14(rand_exe_prng_187_io_out_14),
    .io_out_15(rand_exe_prng_187_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_188 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_188_clock),
    .reset(rand_exe_prng_188_reset),
    .io_out_0(rand_exe_prng_188_io_out_0),
    .io_out_1(rand_exe_prng_188_io_out_1),
    .io_out_2(rand_exe_prng_188_io_out_2),
    .io_out_3(rand_exe_prng_188_io_out_3),
    .io_out_4(rand_exe_prng_188_io_out_4),
    .io_out_5(rand_exe_prng_188_io_out_5),
    .io_out_6(rand_exe_prng_188_io_out_6),
    .io_out_7(rand_exe_prng_188_io_out_7),
    .io_out_8(rand_exe_prng_188_io_out_8),
    .io_out_9(rand_exe_prng_188_io_out_9),
    .io_out_10(rand_exe_prng_188_io_out_10),
    .io_out_11(rand_exe_prng_188_io_out_11),
    .io_out_12(rand_exe_prng_188_io_out_12),
    .io_out_13(rand_exe_prng_188_io_out_13),
    .io_out_14(rand_exe_prng_188_io_out_14),
    .io_out_15(rand_exe_prng_188_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_189 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_189_clock),
    .reset(rand_exe_prng_189_reset),
    .io_out_0(rand_exe_prng_189_io_out_0),
    .io_out_1(rand_exe_prng_189_io_out_1),
    .io_out_2(rand_exe_prng_189_io_out_2),
    .io_out_3(rand_exe_prng_189_io_out_3),
    .io_out_4(rand_exe_prng_189_io_out_4),
    .io_out_5(rand_exe_prng_189_io_out_5),
    .io_out_6(rand_exe_prng_189_io_out_6),
    .io_out_7(rand_exe_prng_189_io_out_7),
    .io_out_8(rand_exe_prng_189_io_out_8),
    .io_out_9(rand_exe_prng_189_io_out_9),
    .io_out_10(rand_exe_prng_189_io_out_10),
    .io_out_11(rand_exe_prng_189_io_out_11),
    .io_out_12(rand_exe_prng_189_io_out_12),
    .io_out_13(rand_exe_prng_189_io_out_13),
    .io_out_14(rand_exe_prng_189_io_out_14),
    .io_out_15(rand_exe_prng_189_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_190 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_190_clock),
    .reset(rand_exe_prng_190_reset),
    .io_out_0(rand_exe_prng_190_io_out_0),
    .io_out_1(rand_exe_prng_190_io_out_1),
    .io_out_2(rand_exe_prng_190_io_out_2),
    .io_out_3(rand_exe_prng_190_io_out_3),
    .io_out_4(rand_exe_prng_190_io_out_4),
    .io_out_5(rand_exe_prng_190_io_out_5),
    .io_out_6(rand_exe_prng_190_io_out_6),
    .io_out_7(rand_exe_prng_190_io_out_7),
    .io_out_8(rand_exe_prng_190_io_out_8),
    .io_out_9(rand_exe_prng_190_io_out_9),
    .io_out_10(rand_exe_prng_190_io_out_10),
    .io_out_11(rand_exe_prng_190_io_out_11),
    .io_out_12(rand_exe_prng_190_io_out_12),
    .io_out_13(rand_exe_prng_190_io_out_13),
    .io_out_14(rand_exe_prng_190_io_out_14),
    .io_out_15(rand_exe_prng_190_io_out_15)
  );
  MaxPeriodFibonacciLFSR rand_exe_prng_191 ( // @[PRNG.scala 82:22]
    .clock(rand_exe_prng_191_clock),
    .reset(rand_exe_prng_191_reset),
    .io_out_0(rand_exe_prng_191_io_out_0),
    .io_out_1(rand_exe_prng_191_io_out_1),
    .io_out_2(rand_exe_prng_191_io_out_2),
    .io_out_3(rand_exe_prng_191_io_out_3),
    .io_out_4(rand_exe_prng_191_io_out_4),
    .io_out_5(rand_exe_prng_191_io_out_5),
    .io_out_6(rand_exe_prng_191_io_out_6),
    .io_out_7(rand_exe_prng_191_io_out_7),
    .io_out_8(rand_exe_prng_191_io_out_8),
    .io_out_9(rand_exe_prng_191_io_out_9),
    .io_out_10(rand_exe_prng_191_io_out_10),
    .io_out_11(rand_exe_prng_191_io_out_11),
    .io_out_12(rand_exe_prng_191_io_out_12),
    .io_out_13(rand_exe_prng_191_io_out_13),
    .io_out_14(rand_exe_prng_191_io_out_14),
    .io_out_15(rand_exe_prng_191_io_out_15)
  );
  assign io_phv_out_data_0 = rand_0[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_1 = rand_0[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_2 = rand_1[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_3 = rand_1[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_4 = rand_2[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_5 = rand_2[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_6 = rand_3[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_7 = rand_3[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_8 = rand_4[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_9 = rand_4[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_10 = rand_5[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_11 = rand_5[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_12 = rand_6[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_13 = rand_6[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_14 = rand_7[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_15 = rand_7[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_16 = rand_8[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_17 = rand_8[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_18 = rand_9[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_19 = rand_9[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_20 = rand_10[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_21 = rand_10[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_22 = rand_11[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_23 = rand_11[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_24 = rand_12[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_25 = rand_12[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_26 = rand_13[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_27 = rand_13[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_28 = rand_14[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_29 = rand_14[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_30 = rand_15[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_31 = rand_15[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_32 = rand_16[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_33 = rand_16[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_34 = rand_17[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_35 = rand_17[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_36 = rand_18[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_37 = rand_18[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_38 = rand_19[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_39 = rand_19[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_40 = rand_20[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_41 = rand_20[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_42 = rand_21[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_43 = rand_21[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_44 = rand_22[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_45 = rand_22[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_46 = rand_23[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_47 = rand_23[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_48 = rand_24[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_49 = rand_24[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_50 = rand_25[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_51 = rand_25[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_52 = rand_26[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_53 = rand_26[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_54 = rand_27[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_55 = rand_27[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_56 = rand_28[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_57 = rand_28[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_58 = rand_29[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_59 = rand_29[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_60 = rand_30[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_61 = rand_30[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_62 = rand_31[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_63 = rand_31[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_64 = rand_32[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_65 = rand_32[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_66 = rand_33[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_67 = rand_33[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_68 = rand_34[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_69 = rand_34[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_70 = rand_35[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_71 = rand_35[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_72 = rand_36[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_73 = rand_36[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_74 = rand_37[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_75 = rand_37[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_76 = rand_38[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_77 = rand_38[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_78 = rand_39[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_79 = rand_39[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_80 = rand_40[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_81 = rand_40[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_82 = rand_41[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_83 = rand_41[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_84 = rand_42[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_85 = rand_42[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_86 = rand_43[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_87 = rand_43[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_88 = rand_44[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_89 = rand_44[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_90 = rand_45[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_91 = rand_45[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_92 = rand_46[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_93 = rand_46[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_94 = rand_47[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_95 = rand_47[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_96 = rand_48[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_97 = rand_48[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_98 = rand_49[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_99 = rand_49[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_100 = rand_50[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_101 = rand_50[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_102 = rand_51[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_103 = rand_51[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_104 = rand_52[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_105 = rand_52[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_106 = rand_53[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_107 = rand_53[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_108 = rand_54[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_109 = rand_54[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_110 = rand_55[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_111 = rand_55[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_112 = rand_56[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_113 = rand_56[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_114 = rand_57[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_115 = rand_57[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_116 = rand_58[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_117 = rand_58[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_118 = rand_59[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_119 = rand_59[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_120 = rand_60[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_121 = rand_60[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_122 = rand_61[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_123 = rand_61[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_124 = rand_62[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_125 = rand_62[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_126 = rand_63[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_127 = rand_63[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_128 = rand_64[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_129 = rand_64[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_130 = rand_65[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_131 = rand_65[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_132 = rand_66[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_133 = rand_66[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_134 = rand_67[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_135 = rand_67[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_136 = rand_68[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_137 = rand_68[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_138 = rand_69[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_139 = rand_69[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_140 = rand_70[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_141 = rand_70[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_142 = rand_71[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_143 = rand_71[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_144 = rand_72[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_145 = rand_72[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_146 = rand_73[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_147 = rand_73[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_148 = rand_74[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_149 = rand_74[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_150 = rand_75[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_151 = rand_75[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_152 = rand_76[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_153 = rand_76[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_154 = rand_77[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_155 = rand_77[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_156 = rand_78[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_157 = rand_78[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_158 = rand_79[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_159 = rand_79[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_160 = rand_80[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_161 = rand_80[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_162 = rand_81[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_163 = rand_81[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_164 = rand_82[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_165 = rand_82[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_166 = rand_83[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_167 = rand_83[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_168 = rand_84[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_169 = rand_84[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_170 = rand_85[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_171 = rand_85[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_172 = rand_86[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_173 = rand_86[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_174 = rand_87[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_175 = rand_87[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_176 = rand_88[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_177 = rand_88[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_178 = rand_89[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_179 = rand_89[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_180 = rand_90[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_181 = rand_90[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_182 = rand_91[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_183 = rand_91[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_184 = rand_92[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_185 = rand_92[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_186 = rand_93[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_187 = rand_93[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_188 = rand_94[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_189 = rand_94[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_190 = rand_95[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_191 = rand_95[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_192 = rand_96[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_193 = rand_96[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_194 = rand_97[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_195 = rand_97[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_196 = rand_98[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_197 = rand_98[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_198 = rand_99[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_199 = rand_99[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_200 = rand_100[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_201 = rand_100[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_202 = rand_101[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_203 = rand_101[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_204 = rand_102[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_205 = rand_102[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_206 = rand_103[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_207 = rand_103[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_208 = rand_104[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_209 = rand_104[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_210 = rand_105[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_211 = rand_105[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_212 = rand_106[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_213 = rand_106[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_214 = rand_107[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_215 = rand_107[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_216 = rand_108[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_217 = rand_108[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_218 = rand_109[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_219 = rand_109[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_220 = rand_110[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_221 = rand_110[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_222 = rand_111[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_223 = rand_111[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_224 = rand_112[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_225 = rand_112[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_226 = rand_113[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_227 = rand_113[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_228 = rand_114[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_229 = rand_114[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_230 = rand_115[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_231 = rand_115[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_232 = rand_116[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_233 = rand_116[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_234 = rand_117[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_235 = rand_117[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_236 = rand_118[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_237 = rand_118[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_238 = rand_119[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_239 = rand_119[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_240 = rand_120[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_241 = rand_120[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_242 = rand_121[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_243 = rand_121[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_244 = rand_122[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_245 = rand_122[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_246 = rand_123[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_247 = rand_123[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_248 = rand_124[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_249 = rand_124[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_250 = rand_125[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_251 = rand_125[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_252 = rand_126[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_253 = rand_126[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_254 = rand_127[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_255 = rand_127[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_256 = rand_128[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_257 = rand_128[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_258 = rand_129[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_259 = rand_129[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_260 = rand_130[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_261 = rand_130[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_262 = rand_131[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_263 = rand_131[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_264 = rand_132[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_265 = rand_132[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_266 = rand_133[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_267 = rand_133[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_268 = rand_134[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_269 = rand_134[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_270 = rand_135[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_271 = rand_135[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_272 = rand_136[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_273 = rand_136[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_274 = rand_137[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_275 = rand_137[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_276 = rand_138[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_277 = rand_138[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_278 = rand_139[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_279 = rand_139[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_280 = rand_140[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_281 = rand_140[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_282 = rand_141[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_283 = rand_141[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_284 = rand_142[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_285 = rand_142[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_286 = rand_143[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_287 = rand_143[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_288 = rand_144[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_289 = rand_144[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_290 = rand_145[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_291 = rand_145[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_292 = rand_146[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_293 = rand_146[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_294 = rand_147[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_295 = rand_147[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_296 = rand_148[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_297 = rand_148[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_298 = rand_149[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_299 = rand_149[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_300 = rand_150[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_301 = rand_150[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_302 = rand_151[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_303 = rand_151[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_304 = rand_152[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_305 = rand_152[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_306 = rand_153[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_307 = rand_153[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_308 = rand_154[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_309 = rand_154[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_310 = rand_155[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_311 = rand_155[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_312 = rand_156[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_313 = rand_156[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_314 = rand_157[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_315 = rand_157[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_316 = rand_158[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_317 = rand_158[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_318 = rand_159[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_319 = rand_159[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_320 = rand_160[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_321 = rand_160[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_322 = rand_161[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_323 = rand_161[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_324 = rand_162[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_325 = rand_162[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_326 = rand_163[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_327 = rand_163[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_328 = rand_164[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_329 = rand_164[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_330 = rand_165[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_331 = rand_165[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_332 = rand_166[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_333 = rand_166[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_334 = rand_167[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_335 = rand_167[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_336 = rand_168[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_337 = rand_168[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_338 = rand_169[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_339 = rand_169[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_340 = rand_170[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_341 = rand_170[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_342 = rand_171[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_343 = rand_171[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_344 = rand_172[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_345 = rand_172[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_346 = rand_173[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_347 = rand_173[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_348 = rand_174[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_349 = rand_174[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_350 = rand_175[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_351 = rand_175[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_352 = rand_176[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_353 = rand_176[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_354 = rand_177[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_355 = rand_177[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_356 = rand_178[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_357 = rand_178[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_358 = rand_179[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_359 = rand_179[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_360 = rand_180[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_361 = rand_180[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_362 = rand_181[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_363 = rand_181[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_364 = rand_182[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_365 = rand_182[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_366 = rand_183[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_367 = rand_183[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_368 = rand_184[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_369 = rand_184[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_370 = rand_185[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_371 = rand_185[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_372 = rand_186[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_373 = rand_186[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_374 = rand_187[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_375 = rand_187[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_376 = rand_188[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_377 = rand_188[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_378 = rand_189[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_379 = rand_189[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_380 = rand_190[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_381 = rand_190[7:0]; // @[inport.scala 19:42]
  assign io_phv_out_data_382 = rand_191[15:8]; // @[inport.scala 18:42]
  assign io_phv_out_data_383 = rand_191[7:0]; // @[inport.scala 19:42]
  assign rand_exe_prng_clock = clock;
  assign rand_exe_prng_reset = reset;
  assign rand_exe_prng_1_clock = clock;
  assign rand_exe_prng_1_reset = reset;
  assign rand_exe_prng_2_clock = clock;
  assign rand_exe_prng_2_reset = reset;
  assign rand_exe_prng_3_clock = clock;
  assign rand_exe_prng_3_reset = reset;
  assign rand_exe_prng_4_clock = clock;
  assign rand_exe_prng_4_reset = reset;
  assign rand_exe_prng_5_clock = clock;
  assign rand_exe_prng_5_reset = reset;
  assign rand_exe_prng_6_clock = clock;
  assign rand_exe_prng_6_reset = reset;
  assign rand_exe_prng_7_clock = clock;
  assign rand_exe_prng_7_reset = reset;
  assign rand_exe_prng_8_clock = clock;
  assign rand_exe_prng_8_reset = reset;
  assign rand_exe_prng_9_clock = clock;
  assign rand_exe_prng_9_reset = reset;
  assign rand_exe_prng_10_clock = clock;
  assign rand_exe_prng_10_reset = reset;
  assign rand_exe_prng_11_clock = clock;
  assign rand_exe_prng_11_reset = reset;
  assign rand_exe_prng_12_clock = clock;
  assign rand_exe_prng_12_reset = reset;
  assign rand_exe_prng_13_clock = clock;
  assign rand_exe_prng_13_reset = reset;
  assign rand_exe_prng_14_clock = clock;
  assign rand_exe_prng_14_reset = reset;
  assign rand_exe_prng_15_clock = clock;
  assign rand_exe_prng_15_reset = reset;
  assign rand_exe_prng_16_clock = clock;
  assign rand_exe_prng_16_reset = reset;
  assign rand_exe_prng_17_clock = clock;
  assign rand_exe_prng_17_reset = reset;
  assign rand_exe_prng_18_clock = clock;
  assign rand_exe_prng_18_reset = reset;
  assign rand_exe_prng_19_clock = clock;
  assign rand_exe_prng_19_reset = reset;
  assign rand_exe_prng_20_clock = clock;
  assign rand_exe_prng_20_reset = reset;
  assign rand_exe_prng_21_clock = clock;
  assign rand_exe_prng_21_reset = reset;
  assign rand_exe_prng_22_clock = clock;
  assign rand_exe_prng_22_reset = reset;
  assign rand_exe_prng_23_clock = clock;
  assign rand_exe_prng_23_reset = reset;
  assign rand_exe_prng_24_clock = clock;
  assign rand_exe_prng_24_reset = reset;
  assign rand_exe_prng_25_clock = clock;
  assign rand_exe_prng_25_reset = reset;
  assign rand_exe_prng_26_clock = clock;
  assign rand_exe_prng_26_reset = reset;
  assign rand_exe_prng_27_clock = clock;
  assign rand_exe_prng_27_reset = reset;
  assign rand_exe_prng_28_clock = clock;
  assign rand_exe_prng_28_reset = reset;
  assign rand_exe_prng_29_clock = clock;
  assign rand_exe_prng_29_reset = reset;
  assign rand_exe_prng_30_clock = clock;
  assign rand_exe_prng_30_reset = reset;
  assign rand_exe_prng_31_clock = clock;
  assign rand_exe_prng_31_reset = reset;
  assign rand_exe_prng_32_clock = clock;
  assign rand_exe_prng_32_reset = reset;
  assign rand_exe_prng_33_clock = clock;
  assign rand_exe_prng_33_reset = reset;
  assign rand_exe_prng_34_clock = clock;
  assign rand_exe_prng_34_reset = reset;
  assign rand_exe_prng_35_clock = clock;
  assign rand_exe_prng_35_reset = reset;
  assign rand_exe_prng_36_clock = clock;
  assign rand_exe_prng_36_reset = reset;
  assign rand_exe_prng_37_clock = clock;
  assign rand_exe_prng_37_reset = reset;
  assign rand_exe_prng_38_clock = clock;
  assign rand_exe_prng_38_reset = reset;
  assign rand_exe_prng_39_clock = clock;
  assign rand_exe_prng_39_reset = reset;
  assign rand_exe_prng_40_clock = clock;
  assign rand_exe_prng_40_reset = reset;
  assign rand_exe_prng_41_clock = clock;
  assign rand_exe_prng_41_reset = reset;
  assign rand_exe_prng_42_clock = clock;
  assign rand_exe_prng_42_reset = reset;
  assign rand_exe_prng_43_clock = clock;
  assign rand_exe_prng_43_reset = reset;
  assign rand_exe_prng_44_clock = clock;
  assign rand_exe_prng_44_reset = reset;
  assign rand_exe_prng_45_clock = clock;
  assign rand_exe_prng_45_reset = reset;
  assign rand_exe_prng_46_clock = clock;
  assign rand_exe_prng_46_reset = reset;
  assign rand_exe_prng_47_clock = clock;
  assign rand_exe_prng_47_reset = reset;
  assign rand_exe_prng_48_clock = clock;
  assign rand_exe_prng_48_reset = reset;
  assign rand_exe_prng_49_clock = clock;
  assign rand_exe_prng_49_reset = reset;
  assign rand_exe_prng_50_clock = clock;
  assign rand_exe_prng_50_reset = reset;
  assign rand_exe_prng_51_clock = clock;
  assign rand_exe_prng_51_reset = reset;
  assign rand_exe_prng_52_clock = clock;
  assign rand_exe_prng_52_reset = reset;
  assign rand_exe_prng_53_clock = clock;
  assign rand_exe_prng_53_reset = reset;
  assign rand_exe_prng_54_clock = clock;
  assign rand_exe_prng_54_reset = reset;
  assign rand_exe_prng_55_clock = clock;
  assign rand_exe_prng_55_reset = reset;
  assign rand_exe_prng_56_clock = clock;
  assign rand_exe_prng_56_reset = reset;
  assign rand_exe_prng_57_clock = clock;
  assign rand_exe_prng_57_reset = reset;
  assign rand_exe_prng_58_clock = clock;
  assign rand_exe_prng_58_reset = reset;
  assign rand_exe_prng_59_clock = clock;
  assign rand_exe_prng_59_reset = reset;
  assign rand_exe_prng_60_clock = clock;
  assign rand_exe_prng_60_reset = reset;
  assign rand_exe_prng_61_clock = clock;
  assign rand_exe_prng_61_reset = reset;
  assign rand_exe_prng_62_clock = clock;
  assign rand_exe_prng_62_reset = reset;
  assign rand_exe_prng_63_clock = clock;
  assign rand_exe_prng_63_reset = reset;
  assign rand_exe_prng_64_clock = clock;
  assign rand_exe_prng_64_reset = reset;
  assign rand_exe_prng_65_clock = clock;
  assign rand_exe_prng_65_reset = reset;
  assign rand_exe_prng_66_clock = clock;
  assign rand_exe_prng_66_reset = reset;
  assign rand_exe_prng_67_clock = clock;
  assign rand_exe_prng_67_reset = reset;
  assign rand_exe_prng_68_clock = clock;
  assign rand_exe_prng_68_reset = reset;
  assign rand_exe_prng_69_clock = clock;
  assign rand_exe_prng_69_reset = reset;
  assign rand_exe_prng_70_clock = clock;
  assign rand_exe_prng_70_reset = reset;
  assign rand_exe_prng_71_clock = clock;
  assign rand_exe_prng_71_reset = reset;
  assign rand_exe_prng_72_clock = clock;
  assign rand_exe_prng_72_reset = reset;
  assign rand_exe_prng_73_clock = clock;
  assign rand_exe_prng_73_reset = reset;
  assign rand_exe_prng_74_clock = clock;
  assign rand_exe_prng_74_reset = reset;
  assign rand_exe_prng_75_clock = clock;
  assign rand_exe_prng_75_reset = reset;
  assign rand_exe_prng_76_clock = clock;
  assign rand_exe_prng_76_reset = reset;
  assign rand_exe_prng_77_clock = clock;
  assign rand_exe_prng_77_reset = reset;
  assign rand_exe_prng_78_clock = clock;
  assign rand_exe_prng_78_reset = reset;
  assign rand_exe_prng_79_clock = clock;
  assign rand_exe_prng_79_reset = reset;
  assign rand_exe_prng_80_clock = clock;
  assign rand_exe_prng_80_reset = reset;
  assign rand_exe_prng_81_clock = clock;
  assign rand_exe_prng_81_reset = reset;
  assign rand_exe_prng_82_clock = clock;
  assign rand_exe_prng_82_reset = reset;
  assign rand_exe_prng_83_clock = clock;
  assign rand_exe_prng_83_reset = reset;
  assign rand_exe_prng_84_clock = clock;
  assign rand_exe_prng_84_reset = reset;
  assign rand_exe_prng_85_clock = clock;
  assign rand_exe_prng_85_reset = reset;
  assign rand_exe_prng_86_clock = clock;
  assign rand_exe_prng_86_reset = reset;
  assign rand_exe_prng_87_clock = clock;
  assign rand_exe_prng_87_reset = reset;
  assign rand_exe_prng_88_clock = clock;
  assign rand_exe_prng_88_reset = reset;
  assign rand_exe_prng_89_clock = clock;
  assign rand_exe_prng_89_reset = reset;
  assign rand_exe_prng_90_clock = clock;
  assign rand_exe_prng_90_reset = reset;
  assign rand_exe_prng_91_clock = clock;
  assign rand_exe_prng_91_reset = reset;
  assign rand_exe_prng_92_clock = clock;
  assign rand_exe_prng_92_reset = reset;
  assign rand_exe_prng_93_clock = clock;
  assign rand_exe_prng_93_reset = reset;
  assign rand_exe_prng_94_clock = clock;
  assign rand_exe_prng_94_reset = reset;
  assign rand_exe_prng_95_clock = clock;
  assign rand_exe_prng_95_reset = reset;
  assign rand_exe_prng_96_clock = clock;
  assign rand_exe_prng_96_reset = reset;
  assign rand_exe_prng_97_clock = clock;
  assign rand_exe_prng_97_reset = reset;
  assign rand_exe_prng_98_clock = clock;
  assign rand_exe_prng_98_reset = reset;
  assign rand_exe_prng_99_clock = clock;
  assign rand_exe_prng_99_reset = reset;
  assign rand_exe_prng_100_clock = clock;
  assign rand_exe_prng_100_reset = reset;
  assign rand_exe_prng_101_clock = clock;
  assign rand_exe_prng_101_reset = reset;
  assign rand_exe_prng_102_clock = clock;
  assign rand_exe_prng_102_reset = reset;
  assign rand_exe_prng_103_clock = clock;
  assign rand_exe_prng_103_reset = reset;
  assign rand_exe_prng_104_clock = clock;
  assign rand_exe_prng_104_reset = reset;
  assign rand_exe_prng_105_clock = clock;
  assign rand_exe_prng_105_reset = reset;
  assign rand_exe_prng_106_clock = clock;
  assign rand_exe_prng_106_reset = reset;
  assign rand_exe_prng_107_clock = clock;
  assign rand_exe_prng_107_reset = reset;
  assign rand_exe_prng_108_clock = clock;
  assign rand_exe_prng_108_reset = reset;
  assign rand_exe_prng_109_clock = clock;
  assign rand_exe_prng_109_reset = reset;
  assign rand_exe_prng_110_clock = clock;
  assign rand_exe_prng_110_reset = reset;
  assign rand_exe_prng_111_clock = clock;
  assign rand_exe_prng_111_reset = reset;
  assign rand_exe_prng_112_clock = clock;
  assign rand_exe_prng_112_reset = reset;
  assign rand_exe_prng_113_clock = clock;
  assign rand_exe_prng_113_reset = reset;
  assign rand_exe_prng_114_clock = clock;
  assign rand_exe_prng_114_reset = reset;
  assign rand_exe_prng_115_clock = clock;
  assign rand_exe_prng_115_reset = reset;
  assign rand_exe_prng_116_clock = clock;
  assign rand_exe_prng_116_reset = reset;
  assign rand_exe_prng_117_clock = clock;
  assign rand_exe_prng_117_reset = reset;
  assign rand_exe_prng_118_clock = clock;
  assign rand_exe_prng_118_reset = reset;
  assign rand_exe_prng_119_clock = clock;
  assign rand_exe_prng_119_reset = reset;
  assign rand_exe_prng_120_clock = clock;
  assign rand_exe_prng_120_reset = reset;
  assign rand_exe_prng_121_clock = clock;
  assign rand_exe_prng_121_reset = reset;
  assign rand_exe_prng_122_clock = clock;
  assign rand_exe_prng_122_reset = reset;
  assign rand_exe_prng_123_clock = clock;
  assign rand_exe_prng_123_reset = reset;
  assign rand_exe_prng_124_clock = clock;
  assign rand_exe_prng_124_reset = reset;
  assign rand_exe_prng_125_clock = clock;
  assign rand_exe_prng_125_reset = reset;
  assign rand_exe_prng_126_clock = clock;
  assign rand_exe_prng_126_reset = reset;
  assign rand_exe_prng_127_clock = clock;
  assign rand_exe_prng_127_reset = reset;
  assign rand_exe_prng_128_clock = clock;
  assign rand_exe_prng_128_reset = reset;
  assign rand_exe_prng_129_clock = clock;
  assign rand_exe_prng_129_reset = reset;
  assign rand_exe_prng_130_clock = clock;
  assign rand_exe_prng_130_reset = reset;
  assign rand_exe_prng_131_clock = clock;
  assign rand_exe_prng_131_reset = reset;
  assign rand_exe_prng_132_clock = clock;
  assign rand_exe_prng_132_reset = reset;
  assign rand_exe_prng_133_clock = clock;
  assign rand_exe_prng_133_reset = reset;
  assign rand_exe_prng_134_clock = clock;
  assign rand_exe_prng_134_reset = reset;
  assign rand_exe_prng_135_clock = clock;
  assign rand_exe_prng_135_reset = reset;
  assign rand_exe_prng_136_clock = clock;
  assign rand_exe_prng_136_reset = reset;
  assign rand_exe_prng_137_clock = clock;
  assign rand_exe_prng_137_reset = reset;
  assign rand_exe_prng_138_clock = clock;
  assign rand_exe_prng_138_reset = reset;
  assign rand_exe_prng_139_clock = clock;
  assign rand_exe_prng_139_reset = reset;
  assign rand_exe_prng_140_clock = clock;
  assign rand_exe_prng_140_reset = reset;
  assign rand_exe_prng_141_clock = clock;
  assign rand_exe_prng_141_reset = reset;
  assign rand_exe_prng_142_clock = clock;
  assign rand_exe_prng_142_reset = reset;
  assign rand_exe_prng_143_clock = clock;
  assign rand_exe_prng_143_reset = reset;
  assign rand_exe_prng_144_clock = clock;
  assign rand_exe_prng_144_reset = reset;
  assign rand_exe_prng_145_clock = clock;
  assign rand_exe_prng_145_reset = reset;
  assign rand_exe_prng_146_clock = clock;
  assign rand_exe_prng_146_reset = reset;
  assign rand_exe_prng_147_clock = clock;
  assign rand_exe_prng_147_reset = reset;
  assign rand_exe_prng_148_clock = clock;
  assign rand_exe_prng_148_reset = reset;
  assign rand_exe_prng_149_clock = clock;
  assign rand_exe_prng_149_reset = reset;
  assign rand_exe_prng_150_clock = clock;
  assign rand_exe_prng_150_reset = reset;
  assign rand_exe_prng_151_clock = clock;
  assign rand_exe_prng_151_reset = reset;
  assign rand_exe_prng_152_clock = clock;
  assign rand_exe_prng_152_reset = reset;
  assign rand_exe_prng_153_clock = clock;
  assign rand_exe_prng_153_reset = reset;
  assign rand_exe_prng_154_clock = clock;
  assign rand_exe_prng_154_reset = reset;
  assign rand_exe_prng_155_clock = clock;
  assign rand_exe_prng_155_reset = reset;
  assign rand_exe_prng_156_clock = clock;
  assign rand_exe_prng_156_reset = reset;
  assign rand_exe_prng_157_clock = clock;
  assign rand_exe_prng_157_reset = reset;
  assign rand_exe_prng_158_clock = clock;
  assign rand_exe_prng_158_reset = reset;
  assign rand_exe_prng_159_clock = clock;
  assign rand_exe_prng_159_reset = reset;
  assign rand_exe_prng_160_clock = clock;
  assign rand_exe_prng_160_reset = reset;
  assign rand_exe_prng_161_clock = clock;
  assign rand_exe_prng_161_reset = reset;
  assign rand_exe_prng_162_clock = clock;
  assign rand_exe_prng_162_reset = reset;
  assign rand_exe_prng_163_clock = clock;
  assign rand_exe_prng_163_reset = reset;
  assign rand_exe_prng_164_clock = clock;
  assign rand_exe_prng_164_reset = reset;
  assign rand_exe_prng_165_clock = clock;
  assign rand_exe_prng_165_reset = reset;
  assign rand_exe_prng_166_clock = clock;
  assign rand_exe_prng_166_reset = reset;
  assign rand_exe_prng_167_clock = clock;
  assign rand_exe_prng_167_reset = reset;
  assign rand_exe_prng_168_clock = clock;
  assign rand_exe_prng_168_reset = reset;
  assign rand_exe_prng_169_clock = clock;
  assign rand_exe_prng_169_reset = reset;
  assign rand_exe_prng_170_clock = clock;
  assign rand_exe_prng_170_reset = reset;
  assign rand_exe_prng_171_clock = clock;
  assign rand_exe_prng_171_reset = reset;
  assign rand_exe_prng_172_clock = clock;
  assign rand_exe_prng_172_reset = reset;
  assign rand_exe_prng_173_clock = clock;
  assign rand_exe_prng_173_reset = reset;
  assign rand_exe_prng_174_clock = clock;
  assign rand_exe_prng_174_reset = reset;
  assign rand_exe_prng_175_clock = clock;
  assign rand_exe_prng_175_reset = reset;
  assign rand_exe_prng_176_clock = clock;
  assign rand_exe_prng_176_reset = reset;
  assign rand_exe_prng_177_clock = clock;
  assign rand_exe_prng_177_reset = reset;
  assign rand_exe_prng_178_clock = clock;
  assign rand_exe_prng_178_reset = reset;
  assign rand_exe_prng_179_clock = clock;
  assign rand_exe_prng_179_reset = reset;
  assign rand_exe_prng_180_clock = clock;
  assign rand_exe_prng_180_reset = reset;
  assign rand_exe_prng_181_clock = clock;
  assign rand_exe_prng_181_reset = reset;
  assign rand_exe_prng_182_clock = clock;
  assign rand_exe_prng_182_reset = reset;
  assign rand_exe_prng_183_clock = clock;
  assign rand_exe_prng_183_reset = reset;
  assign rand_exe_prng_184_clock = clock;
  assign rand_exe_prng_184_reset = reset;
  assign rand_exe_prng_185_clock = clock;
  assign rand_exe_prng_185_reset = reset;
  assign rand_exe_prng_186_clock = clock;
  assign rand_exe_prng_186_reset = reset;
  assign rand_exe_prng_187_clock = clock;
  assign rand_exe_prng_187_reset = reset;
  assign rand_exe_prng_188_clock = clock;
  assign rand_exe_prng_188_reset = reset;
  assign rand_exe_prng_189_clock = clock;
  assign rand_exe_prng_189_reset = reset;
  assign rand_exe_prng_190_clock = clock;
  assign rand_exe_prng_190_reset = reset;
  assign rand_exe_prng_191_clock = clock;
  assign rand_exe_prng_191_reset = reset;
endmodule
