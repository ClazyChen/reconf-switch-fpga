module Parser(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_en,
  input         io_mod_last_mau_id_mod,
  input  [1:0]  io_mod_last_mau_id,
  input  [1:0]  io_mod_cs,
  input         io_mod_module_mod_state_id_mod,
  input  [7:0]  io_mod_module_mod_state_id,
  input         io_mod_module_mod_sram_w_cs,
  input         io_mod_module_mod_sram_w_en,
  input  [7:0]  io_mod_module_mod_sram_w_addr,
  input  [63:0] io_mod_module_mod_sram_w_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mau_0_clock; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_0_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_0_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_0_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_0_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_0_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_0_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_0_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_0_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_0_io_mod_sram_w_data; // @[parser.scala 21:25]
  wire  mau_1_clock; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_1_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_1_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_1_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_1_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_1_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_1_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_1_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_1_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_1_io_mod_sram_w_data; // @[parser.scala 21:25]
  wire  mau_2_clock; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_2_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_2_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_2_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_2_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_2_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_2_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_2_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_2_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_2_io_mod_sram_w_data; // @[parser.scala 21:25]
  wire  mau_3_clock; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_in_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_in_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_3_io_pipe_phv_in_next_processor_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_in_next_config_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_in_is_valid_processor; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_0; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_1; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_2; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_3; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_4; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_5; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_6; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_7; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_8; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_9; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_10; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_11; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_12; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_13; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_14; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_16; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_17; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_18; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_19; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_20; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_21; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_22; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_23; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_24; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_25; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_26; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_27; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_28; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_29; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_30; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_31; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_32; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_33; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_34; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_35; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_36; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_37; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_38; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_39; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_40; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_41; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_42; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_43; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_44; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_45; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_46; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_47; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_48; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_49; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_50; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_51; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_52; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_53; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_54; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_55; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_56; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_57; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_58; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_59; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_60; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_61; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_62; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_63; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_64; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_65; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_66; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_67; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_68; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_69; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_70; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_71; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_72; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_73; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_74; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_75; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_76; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_77; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_78; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_79; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_80; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_81; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_82; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_83; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_84; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_85; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_86; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_87; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_88; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_89; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_90; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_91; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_92; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_93; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_94; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_95; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_96; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_97; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_98; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_99; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_100; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_101; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_102; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_103; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_104; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_105; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_106; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_107; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_108; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_109; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_110; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_111; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_112; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_113; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_114; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_115; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_116; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_117; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_118; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_119; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_120; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_121; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_122; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_123; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_124; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_125; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_126; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_127; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_128; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_129; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_130; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_131; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_132; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_133; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_134; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_135; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_136; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_137; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_138; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_139; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_140; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_141; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_142; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_143; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_144; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_145; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_146; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_147; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_148; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_149; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_150; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_151; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_152; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_153; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_154; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_155; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_156; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_157; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_158; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_159; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_160; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_161; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_162; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_163; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_164; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_165; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_166; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_167; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_168; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_169; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_170; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_171; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_172; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_173; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_174; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_175; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_176; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_177; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_178; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_179; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_180; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_181; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_182; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_183; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_184; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_185; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_186; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_187; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_188; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_189; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_190; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_191; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_192; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_193; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_194; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_195; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_196; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_197; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_198; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_199; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_200; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_201; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_202; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_203; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_204; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_205; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_206; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_207; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_208; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_209; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_210; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_211; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_212; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_213; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_214; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_215; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_216; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_217; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_218; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_219; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_220; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_221; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_222; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_223; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_224; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_225; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_226; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_227; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_228; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_229; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_230; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_231; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_232; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_233; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_234; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_235; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_236; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_237; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_238; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_239; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_240; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_241; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_242; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_243; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_244; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_245; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_246; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_247; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_248; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_249; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_250; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_251; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_252; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_253; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_254; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_255; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_256; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_257; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_258; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_259; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_260; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_261; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_262; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_263; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_264; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_265; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_266; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_267; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_268; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_269; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_270; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_271; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_272; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_273; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_274; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_275; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_276; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_277; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_278; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_279; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_280; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_281; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_282; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_283; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_284; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_285; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_286; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_287; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_288; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_289; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_290; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_291; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_292; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_293; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_294; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_295; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_296; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_297; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_298; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_299; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_300; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_301; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_302; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_303; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_304; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_305; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_306; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_307; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_308; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_309; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_310; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_311; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_312; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_313; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_314; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_315; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_316; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_317; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_318; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_319; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_320; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_321; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_322; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_323; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_324; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_325; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_326; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_327; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_328; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_329; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_330; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_331; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_332; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_333; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_334; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_335; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_336; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_337; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_338; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_339; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_340; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_341; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_342; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_343; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_344; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_345; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_346; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_347; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_348; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_349; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_350; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_351; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_352; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_353; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_354; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_355; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_356; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_357; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_358; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_359; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_360; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_361; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_362; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_363; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_364; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_365; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_366; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_367; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_368; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_369; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_370; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_371; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_372; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_373; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_374; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_375; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_376; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_377; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_378; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_379; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_380; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_381; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_382; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_383; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_384; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_385; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_386; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_387; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_388; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_389; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_390; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_391; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_392; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_393; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_394; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_395; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_396; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_397; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_398; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_399; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_400; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_401; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_402; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_403; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_404; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_405; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_406; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_407; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_408; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_409; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_410; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_411; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_412; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_413; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_414; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_415; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_416; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_417; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_418; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_419; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_420; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_421; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_422; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_423; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_424; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_425; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_426; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_427; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_428; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_429; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_430; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_431; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_432; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_433; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_434; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_435; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_436; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_437; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_438; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_439; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_440; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_441; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_442; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_443; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_444; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_445; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_446; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_447; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_448; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_449; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_450; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_451; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_452; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_453; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_454; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_455; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_456; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_457; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_458; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_459; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_460; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_461; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_462; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_463; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_464; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_465; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_466; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_467; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_468; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_469; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_470; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_471; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_472; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_473; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_474; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_475; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_476; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_477; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_478; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_479; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_480; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_481; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_482; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_483; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_484; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_485; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_486; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_487; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_488; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_489; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_490; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_491; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_492; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_493; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_494; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_495; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_496; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_497; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_498; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_499; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_500; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_501; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_502; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_503; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_504; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_505; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_506; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_507; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_508; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_509; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_510; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_data_511; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_0; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_1; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_2; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_3; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_4; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_5; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_6; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_7; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_8; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_9; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_10; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_11; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_12; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_13; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_14; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_header_15; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_state; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_pipe_phv_out_parse_current_offset; // @[parser.scala 21:25]
  wire [15:0] mau_3_io_pipe_phv_out_parse_transition_field; // @[parser.scala 21:25]
  wire [3:0] mau_3_io_pipe_phv_out_next_processor_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_out_next_config_id; // @[parser.scala 21:25]
  wire  mau_3_io_pipe_phv_out_is_valid_processor; // @[parser.scala 21:25]
  wire  mau_3_io_mod_state_id_mod; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_mod_state_id; // @[parser.scala 21:25]
  wire  mau_3_io_mod_sram_w_cs; // @[parser.scala 21:25]
  wire  mau_3_io_mod_sram_w_en; // @[parser.scala 21:25]
  wire [7:0] mau_3_io_mod_sram_w_addr; // @[parser.scala 21:25]
  wire [63:0] mau_3_io_mod_sram_w_data; // @[parser.scala 21:25]
  reg [2:0] last_mau_id; // @[parser.scala 14:26]
  wire  _GEN_0 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_is_valid_processor : io_pipe_phv_in_is_valid_processor; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire  _GEN_1 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_next_config_id : io_pipe_phv_in_next_config_id; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [3:0] _GEN_2 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_next_processor_id : io_pipe_phv_in_next_processor_id; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_3 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_parse_transition_field :
    io_pipe_phv_in_parse_transition_field; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_4 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_parse_current_offset :
    io_pipe_phv_in_parse_current_offset; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_5 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_parse_current_state :
    io_pipe_phv_in_parse_current_state; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_6 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_0 : io_pipe_phv_in_header_0; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_7 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_1 : io_pipe_phv_in_header_1; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_8 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_2 : io_pipe_phv_in_header_2; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_9 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_3 : io_pipe_phv_in_header_3; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_10 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_4 : io_pipe_phv_in_header_4; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_11 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_5 : io_pipe_phv_in_header_5; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_12 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_6 : io_pipe_phv_in_header_6; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_13 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_7 : io_pipe_phv_in_header_7; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_14 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_8 : io_pipe_phv_in_header_8; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_15 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_9 : io_pipe_phv_in_header_9; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_16 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_10 : io_pipe_phv_in_header_10; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_17 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_11 : io_pipe_phv_in_header_11; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_18 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_12 : io_pipe_phv_in_header_12; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_19 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_13 : io_pipe_phv_in_header_13; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_20 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_14 : io_pipe_phv_in_header_14; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [15:0] _GEN_21 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_header_15 : io_pipe_phv_in_header_15; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_22 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_0 : io_pipe_phv_in_data_0; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_23 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_1 : io_pipe_phv_in_data_1; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_24 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_2 : io_pipe_phv_in_data_2; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_25 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_3 : io_pipe_phv_in_data_3; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_26 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_4 : io_pipe_phv_in_data_4; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_27 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_5 : io_pipe_phv_in_data_5; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_28 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_6 : io_pipe_phv_in_data_6; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_29 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_7 : io_pipe_phv_in_data_7; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_30 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_8 : io_pipe_phv_in_data_8; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_31 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_9 : io_pipe_phv_in_data_9; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_32 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_10 : io_pipe_phv_in_data_10; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_33 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_11 : io_pipe_phv_in_data_11; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_34 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_12 : io_pipe_phv_in_data_12; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_35 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_13 : io_pipe_phv_in_data_13; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_36 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_14 : io_pipe_phv_in_data_14; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_37 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_15 : io_pipe_phv_in_data_15; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_38 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_16 : io_pipe_phv_in_data_16; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_39 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_17 : io_pipe_phv_in_data_17; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_40 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_18 : io_pipe_phv_in_data_18; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_41 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_19 : io_pipe_phv_in_data_19; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_42 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_20 : io_pipe_phv_in_data_20; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_43 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_21 : io_pipe_phv_in_data_21; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_44 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_22 : io_pipe_phv_in_data_22; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_45 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_23 : io_pipe_phv_in_data_23; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_46 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_24 : io_pipe_phv_in_data_24; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_47 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_25 : io_pipe_phv_in_data_25; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_48 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_26 : io_pipe_phv_in_data_26; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_49 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_27 : io_pipe_phv_in_data_27; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_50 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_28 : io_pipe_phv_in_data_28; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_51 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_29 : io_pipe_phv_in_data_29; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_52 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_30 : io_pipe_phv_in_data_30; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_53 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_31 : io_pipe_phv_in_data_31; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_54 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_32 : io_pipe_phv_in_data_32; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_55 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_33 : io_pipe_phv_in_data_33; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_56 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_34 : io_pipe_phv_in_data_34; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_57 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_35 : io_pipe_phv_in_data_35; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_58 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_36 : io_pipe_phv_in_data_36; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_59 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_37 : io_pipe_phv_in_data_37; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_60 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_38 : io_pipe_phv_in_data_38; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_61 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_39 : io_pipe_phv_in_data_39; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_62 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_40 : io_pipe_phv_in_data_40; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_63 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_41 : io_pipe_phv_in_data_41; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_64 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_42 : io_pipe_phv_in_data_42; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_65 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_43 : io_pipe_phv_in_data_43; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_66 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_44 : io_pipe_phv_in_data_44; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_67 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_45 : io_pipe_phv_in_data_45; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_68 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_46 : io_pipe_phv_in_data_46; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_69 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_47 : io_pipe_phv_in_data_47; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_70 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_48 : io_pipe_phv_in_data_48; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_71 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_49 : io_pipe_phv_in_data_49; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_72 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_50 : io_pipe_phv_in_data_50; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_73 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_51 : io_pipe_phv_in_data_51; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_74 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_52 : io_pipe_phv_in_data_52; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_75 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_53 : io_pipe_phv_in_data_53; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_76 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_54 : io_pipe_phv_in_data_54; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_77 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_55 : io_pipe_phv_in_data_55; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_78 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_56 : io_pipe_phv_in_data_56; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_79 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_57 : io_pipe_phv_in_data_57; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_80 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_58 : io_pipe_phv_in_data_58; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_81 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_59 : io_pipe_phv_in_data_59; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_82 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_60 : io_pipe_phv_in_data_60; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_83 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_61 : io_pipe_phv_in_data_61; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_84 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_62 : io_pipe_phv_in_data_62; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_85 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_63 : io_pipe_phv_in_data_63; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_86 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_64 : io_pipe_phv_in_data_64; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_87 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_65 : io_pipe_phv_in_data_65; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_88 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_66 : io_pipe_phv_in_data_66; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_89 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_67 : io_pipe_phv_in_data_67; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_90 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_68 : io_pipe_phv_in_data_68; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_91 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_69 : io_pipe_phv_in_data_69; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_92 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_70 : io_pipe_phv_in_data_70; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_93 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_71 : io_pipe_phv_in_data_71; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_94 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_72 : io_pipe_phv_in_data_72; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_95 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_73 : io_pipe_phv_in_data_73; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_96 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_74 : io_pipe_phv_in_data_74; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_97 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_75 : io_pipe_phv_in_data_75; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_98 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_76 : io_pipe_phv_in_data_76; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_99 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_77 : io_pipe_phv_in_data_77; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_100 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_78 : io_pipe_phv_in_data_78; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_101 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_79 : io_pipe_phv_in_data_79; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_102 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_80 : io_pipe_phv_in_data_80; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_103 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_81 : io_pipe_phv_in_data_81; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_104 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_82 : io_pipe_phv_in_data_82; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_105 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_83 : io_pipe_phv_in_data_83; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_106 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_84 : io_pipe_phv_in_data_84; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_107 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_85 : io_pipe_phv_in_data_85; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_108 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_86 : io_pipe_phv_in_data_86; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_109 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_87 : io_pipe_phv_in_data_87; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_110 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_88 : io_pipe_phv_in_data_88; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_111 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_89 : io_pipe_phv_in_data_89; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_112 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_90 : io_pipe_phv_in_data_90; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_113 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_91 : io_pipe_phv_in_data_91; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_114 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_92 : io_pipe_phv_in_data_92; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_115 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_93 : io_pipe_phv_in_data_93; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_116 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_94 : io_pipe_phv_in_data_94; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_117 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_95 : io_pipe_phv_in_data_95; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_118 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_96 : io_pipe_phv_in_data_96; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_119 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_97 : io_pipe_phv_in_data_97; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_120 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_98 : io_pipe_phv_in_data_98; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_121 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_99 : io_pipe_phv_in_data_99; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_122 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_100 : io_pipe_phv_in_data_100; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_123 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_101 : io_pipe_phv_in_data_101; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_124 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_102 : io_pipe_phv_in_data_102; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_125 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_103 : io_pipe_phv_in_data_103; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_126 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_104 : io_pipe_phv_in_data_104; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_127 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_105 : io_pipe_phv_in_data_105; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_128 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_106 : io_pipe_phv_in_data_106; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_129 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_107 : io_pipe_phv_in_data_107; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_130 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_108 : io_pipe_phv_in_data_108; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_131 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_109 : io_pipe_phv_in_data_109; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_132 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_110 : io_pipe_phv_in_data_110; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_133 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_111 : io_pipe_phv_in_data_111; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_134 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_112 : io_pipe_phv_in_data_112; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_135 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_113 : io_pipe_phv_in_data_113; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_136 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_114 : io_pipe_phv_in_data_114; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_137 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_115 : io_pipe_phv_in_data_115; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_138 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_116 : io_pipe_phv_in_data_116; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_139 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_117 : io_pipe_phv_in_data_117; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_140 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_118 : io_pipe_phv_in_data_118; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_141 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_119 : io_pipe_phv_in_data_119; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_142 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_120 : io_pipe_phv_in_data_120; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_143 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_121 : io_pipe_phv_in_data_121; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_144 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_122 : io_pipe_phv_in_data_122; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_145 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_123 : io_pipe_phv_in_data_123; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_146 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_124 : io_pipe_phv_in_data_124; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_147 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_125 : io_pipe_phv_in_data_125; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_148 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_126 : io_pipe_phv_in_data_126; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_149 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_127 : io_pipe_phv_in_data_127; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_150 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_128 : io_pipe_phv_in_data_128; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_151 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_129 : io_pipe_phv_in_data_129; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_152 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_130 : io_pipe_phv_in_data_130; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_153 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_131 : io_pipe_phv_in_data_131; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_154 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_132 : io_pipe_phv_in_data_132; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_155 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_133 : io_pipe_phv_in_data_133; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_156 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_134 : io_pipe_phv_in_data_134; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_157 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_135 : io_pipe_phv_in_data_135; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_158 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_136 : io_pipe_phv_in_data_136; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_159 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_137 : io_pipe_phv_in_data_137; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_160 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_138 : io_pipe_phv_in_data_138; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_161 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_139 : io_pipe_phv_in_data_139; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_162 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_140 : io_pipe_phv_in_data_140; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_163 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_141 : io_pipe_phv_in_data_141; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_164 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_142 : io_pipe_phv_in_data_142; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_165 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_143 : io_pipe_phv_in_data_143; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_166 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_144 : io_pipe_phv_in_data_144; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_167 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_145 : io_pipe_phv_in_data_145; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_168 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_146 : io_pipe_phv_in_data_146; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_169 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_147 : io_pipe_phv_in_data_147; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_170 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_148 : io_pipe_phv_in_data_148; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_171 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_149 : io_pipe_phv_in_data_149; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_172 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_150 : io_pipe_phv_in_data_150; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_173 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_151 : io_pipe_phv_in_data_151; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_174 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_152 : io_pipe_phv_in_data_152; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_175 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_153 : io_pipe_phv_in_data_153; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_176 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_154 : io_pipe_phv_in_data_154; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_177 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_155 : io_pipe_phv_in_data_155; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_178 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_156 : io_pipe_phv_in_data_156; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_179 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_157 : io_pipe_phv_in_data_157; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_180 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_158 : io_pipe_phv_in_data_158; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_181 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_159 : io_pipe_phv_in_data_159; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_182 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_160 : io_pipe_phv_in_data_160; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_183 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_161 : io_pipe_phv_in_data_161; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_184 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_162 : io_pipe_phv_in_data_162; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_185 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_163 : io_pipe_phv_in_data_163; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_186 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_164 : io_pipe_phv_in_data_164; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_187 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_165 : io_pipe_phv_in_data_165; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_188 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_166 : io_pipe_phv_in_data_166; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_189 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_167 : io_pipe_phv_in_data_167; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_190 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_168 : io_pipe_phv_in_data_168; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_191 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_169 : io_pipe_phv_in_data_169; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_192 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_170 : io_pipe_phv_in_data_170; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_193 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_171 : io_pipe_phv_in_data_171; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_194 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_172 : io_pipe_phv_in_data_172; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_195 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_173 : io_pipe_phv_in_data_173; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_196 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_174 : io_pipe_phv_in_data_174; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_197 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_175 : io_pipe_phv_in_data_175; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_198 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_176 : io_pipe_phv_in_data_176; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_199 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_177 : io_pipe_phv_in_data_177; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_200 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_178 : io_pipe_phv_in_data_178; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_201 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_179 : io_pipe_phv_in_data_179; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_202 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_180 : io_pipe_phv_in_data_180; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_203 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_181 : io_pipe_phv_in_data_181; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_204 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_182 : io_pipe_phv_in_data_182; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_205 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_183 : io_pipe_phv_in_data_183; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_206 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_184 : io_pipe_phv_in_data_184; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_207 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_185 : io_pipe_phv_in_data_185; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_208 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_186 : io_pipe_phv_in_data_186; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_209 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_187 : io_pipe_phv_in_data_187; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_210 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_188 : io_pipe_phv_in_data_188; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_211 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_189 : io_pipe_phv_in_data_189; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_212 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_190 : io_pipe_phv_in_data_190; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_213 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_191 : io_pipe_phv_in_data_191; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_214 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_192 : io_pipe_phv_in_data_192; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_215 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_193 : io_pipe_phv_in_data_193; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_216 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_194 : io_pipe_phv_in_data_194; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_217 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_195 : io_pipe_phv_in_data_195; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_218 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_196 : io_pipe_phv_in_data_196; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_219 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_197 : io_pipe_phv_in_data_197; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_220 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_198 : io_pipe_phv_in_data_198; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_221 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_199 : io_pipe_phv_in_data_199; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_222 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_200 : io_pipe_phv_in_data_200; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_223 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_201 : io_pipe_phv_in_data_201; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_224 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_202 : io_pipe_phv_in_data_202; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_225 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_203 : io_pipe_phv_in_data_203; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_226 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_204 : io_pipe_phv_in_data_204; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_227 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_205 : io_pipe_phv_in_data_205; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_228 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_206 : io_pipe_phv_in_data_206; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_229 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_207 : io_pipe_phv_in_data_207; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_230 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_208 : io_pipe_phv_in_data_208; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_231 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_209 : io_pipe_phv_in_data_209; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_232 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_210 : io_pipe_phv_in_data_210; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_233 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_211 : io_pipe_phv_in_data_211; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_234 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_212 : io_pipe_phv_in_data_212; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_235 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_213 : io_pipe_phv_in_data_213; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_236 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_214 : io_pipe_phv_in_data_214; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_237 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_215 : io_pipe_phv_in_data_215; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_238 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_216 : io_pipe_phv_in_data_216; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_239 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_217 : io_pipe_phv_in_data_217; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_240 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_218 : io_pipe_phv_in_data_218; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_241 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_219 : io_pipe_phv_in_data_219; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_242 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_220 : io_pipe_phv_in_data_220; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_243 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_221 : io_pipe_phv_in_data_221; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_244 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_222 : io_pipe_phv_in_data_222; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_245 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_223 : io_pipe_phv_in_data_223; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_246 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_224 : io_pipe_phv_in_data_224; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_247 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_225 : io_pipe_phv_in_data_225; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_248 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_226 : io_pipe_phv_in_data_226; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_249 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_227 : io_pipe_phv_in_data_227; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_250 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_228 : io_pipe_phv_in_data_228; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_251 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_229 : io_pipe_phv_in_data_229; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_252 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_230 : io_pipe_phv_in_data_230; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_253 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_231 : io_pipe_phv_in_data_231; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_254 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_232 : io_pipe_phv_in_data_232; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_255 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_233 : io_pipe_phv_in_data_233; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_256 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_234 : io_pipe_phv_in_data_234; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_257 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_235 : io_pipe_phv_in_data_235; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_258 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_236 : io_pipe_phv_in_data_236; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_259 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_237 : io_pipe_phv_in_data_237; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_260 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_238 : io_pipe_phv_in_data_238; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_261 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_239 : io_pipe_phv_in_data_239; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_262 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_240 : io_pipe_phv_in_data_240; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_263 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_241 : io_pipe_phv_in_data_241; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_264 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_242 : io_pipe_phv_in_data_242; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_265 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_243 : io_pipe_phv_in_data_243; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_266 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_244 : io_pipe_phv_in_data_244; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_267 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_245 : io_pipe_phv_in_data_245; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_268 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_246 : io_pipe_phv_in_data_246; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_269 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_247 : io_pipe_phv_in_data_247; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_270 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_248 : io_pipe_phv_in_data_248; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_271 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_249 : io_pipe_phv_in_data_249; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_272 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_250 : io_pipe_phv_in_data_250; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_273 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_251 : io_pipe_phv_in_data_251; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_274 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_252 : io_pipe_phv_in_data_252; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_275 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_253 : io_pipe_phv_in_data_253; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_276 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_254 : io_pipe_phv_in_data_254; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_277 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_255 : io_pipe_phv_in_data_255; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_278 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_256 : io_pipe_phv_in_data_256; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_279 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_257 : io_pipe_phv_in_data_257; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_280 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_258 : io_pipe_phv_in_data_258; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_281 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_259 : io_pipe_phv_in_data_259; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_282 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_260 : io_pipe_phv_in_data_260; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_283 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_261 : io_pipe_phv_in_data_261; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_284 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_262 : io_pipe_phv_in_data_262; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_285 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_263 : io_pipe_phv_in_data_263; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_286 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_264 : io_pipe_phv_in_data_264; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_287 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_265 : io_pipe_phv_in_data_265; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_288 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_266 : io_pipe_phv_in_data_266; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_289 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_267 : io_pipe_phv_in_data_267; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_290 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_268 : io_pipe_phv_in_data_268; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_291 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_269 : io_pipe_phv_in_data_269; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_292 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_270 : io_pipe_phv_in_data_270; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_293 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_271 : io_pipe_phv_in_data_271; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_294 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_272 : io_pipe_phv_in_data_272; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_295 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_273 : io_pipe_phv_in_data_273; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_296 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_274 : io_pipe_phv_in_data_274; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_297 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_275 : io_pipe_phv_in_data_275; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_298 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_276 : io_pipe_phv_in_data_276; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_299 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_277 : io_pipe_phv_in_data_277; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_300 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_278 : io_pipe_phv_in_data_278; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_301 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_279 : io_pipe_phv_in_data_279; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_302 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_280 : io_pipe_phv_in_data_280; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_303 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_281 : io_pipe_phv_in_data_281; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_304 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_282 : io_pipe_phv_in_data_282; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_305 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_283 : io_pipe_phv_in_data_283; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_306 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_284 : io_pipe_phv_in_data_284; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_307 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_285 : io_pipe_phv_in_data_285; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_308 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_286 : io_pipe_phv_in_data_286; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_309 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_287 : io_pipe_phv_in_data_287; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_310 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_288 : io_pipe_phv_in_data_288; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_311 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_289 : io_pipe_phv_in_data_289; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_312 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_290 : io_pipe_phv_in_data_290; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_313 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_291 : io_pipe_phv_in_data_291; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_314 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_292 : io_pipe_phv_in_data_292; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_315 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_293 : io_pipe_phv_in_data_293; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_316 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_294 : io_pipe_phv_in_data_294; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_317 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_295 : io_pipe_phv_in_data_295; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_318 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_296 : io_pipe_phv_in_data_296; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_319 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_297 : io_pipe_phv_in_data_297; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_320 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_298 : io_pipe_phv_in_data_298; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_321 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_299 : io_pipe_phv_in_data_299; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_322 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_300 : io_pipe_phv_in_data_300; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_323 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_301 : io_pipe_phv_in_data_301; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_324 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_302 : io_pipe_phv_in_data_302; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_325 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_303 : io_pipe_phv_in_data_303; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_326 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_304 : io_pipe_phv_in_data_304; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_327 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_305 : io_pipe_phv_in_data_305; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_328 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_306 : io_pipe_phv_in_data_306; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_329 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_307 : io_pipe_phv_in_data_307; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_330 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_308 : io_pipe_phv_in_data_308; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_331 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_309 : io_pipe_phv_in_data_309; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_332 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_310 : io_pipe_phv_in_data_310; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_333 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_311 : io_pipe_phv_in_data_311; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_334 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_312 : io_pipe_phv_in_data_312; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_335 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_313 : io_pipe_phv_in_data_313; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_336 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_314 : io_pipe_phv_in_data_314; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_337 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_315 : io_pipe_phv_in_data_315; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_338 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_316 : io_pipe_phv_in_data_316; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_339 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_317 : io_pipe_phv_in_data_317; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_340 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_318 : io_pipe_phv_in_data_318; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_341 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_319 : io_pipe_phv_in_data_319; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_342 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_320 : io_pipe_phv_in_data_320; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_343 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_321 : io_pipe_phv_in_data_321; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_344 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_322 : io_pipe_phv_in_data_322; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_345 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_323 : io_pipe_phv_in_data_323; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_346 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_324 : io_pipe_phv_in_data_324; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_347 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_325 : io_pipe_phv_in_data_325; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_348 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_326 : io_pipe_phv_in_data_326; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_349 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_327 : io_pipe_phv_in_data_327; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_350 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_328 : io_pipe_phv_in_data_328; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_351 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_329 : io_pipe_phv_in_data_329; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_352 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_330 : io_pipe_phv_in_data_330; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_353 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_331 : io_pipe_phv_in_data_331; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_354 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_332 : io_pipe_phv_in_data_332; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_355 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_333 : io_pipe_phv_in_data_333; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_356 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_334 : io_pipe_phv_in_data_334; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_357 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_335 : io_pipe_phv_in_data_335; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_358 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_336 : io_pipe_phv_in_data_336; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_359 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_337 : io_pipe_phv_in_data_337; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_360 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_338 : io_pipe_phv_in_data_338; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_361 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_339 : io_pipe_phv_in_data_339; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_362 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_340 : io_pipe_phv_in_data_340; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_363 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_341 : io_pipe_phv_in_data_341; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_364 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_342 : io_pipe_phv_in_data_342; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_365 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_343 : io_pipe_phv_in_data_343; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_366 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_344 : io_pipe_phv_in_data_344; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_367 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_345 : io_pipe_phv_in_data_345; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_368 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_346 : io_pipe_phv_in_data_346; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_369 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_347 : io_pipe_phv_in_data_347; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_370 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_348 : io_pipe_phv_in_data_348; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_371 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_349 : io_pipe_phv_in_data_349; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_372 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_350 : io_pipe_phv_in_data_350; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_373 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_351 : io_pipe_phv_in_data_351; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_374 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_352 : io_pipe_phv_in_data_352; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_375 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_353 : io_pipe_phv_in_data_353; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_376 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_354 : io_pipe_phv_in_data_354; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_377 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_355 : io_pipe_phv_in_data_355; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_378 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_356 : io_pipe_phv_in_data_356; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_379 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_357 : io_pipe_phv_in_data_357; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_380 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_358 : io_pipe_phv_in_data_358; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_381 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_359 : io_pipe_phv_in_data_359; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_382 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_360 : io_pipe_phv_in_data_360; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_383 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_361 : io_pipe_phv_in_data_361; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_384 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_362 : io_pipe_phv_in_data_362; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_385 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_363 : io_pipe_phv_in_data_363; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_386 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_364 : io_pipe_phv_in_data_364; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_387 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_365 : io_pipe_phv_in_data_365; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_388 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_366 : io_pipe_phv_in_data_366; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_389 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_367 : io_pipe_phv_in_data_367; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_390 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_368 : io_pipe_phv_in_data_368; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_391 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_369 : io_pipe_phv_in_data_369; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_392 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_370 : io_pipe_phv_in_data_370; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_393 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_371 : io_pipe_phv_in_data_371; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_394 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_372 : io_pipe_phv_in_data_372; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_395 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_373 : io_pipe_phv_in_data_373; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_396 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_374 : io_pipe_phv_in_data_374; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_397 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_375 : io_pipe_phv_in_data_375; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_398 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_376 : io_pipe_phv_in_data_376; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_399 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_377 : io_pipe_phv_in_data_377; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_400 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_378 : io_pipe_phv_in_data_378; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_401 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_379 : io_pipe_phv_in_data_379; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_402 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_380 : io_pipe_phv_in_data_380; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_403 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_381 : io_pipe_phv_in_data_381; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_404 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_382 : io_pipe_phv_in_data_382; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_405 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_383 : io_pipe_phv_in_data_383; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_406 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_384 : io_pipe_phv_in_data_384; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_407 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_385 : io_pipe_phv_in_data_385; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_408 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_386 : io_pipe_phv_in_data_386; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_409 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_387 : io_pipe_phv_in_data_387; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_410 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_388 : io_pipe_phv_in_data_388; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_411 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_389 : io_pipe_phv_in_data_389; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_412 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_390 : io_pipe_phv_in_data_390; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_413 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_391 : io_pipe_phv_in_data_391; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_414 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_392 : io_pipe_phv_in_data_392; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_415 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_393 : io_pipe_phv_in_data_393; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_416 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_394 : io_pipe_phv_in_data_394; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_417 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_395 : io_pipe_phv_in_data_395; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_418 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_396 : io_pipe_phv_in_data_396; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_419 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_397 : io_pipe_phv_in_data_397; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_420 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_398 : io_pipe_phv_in_data_398; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_421 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_399 : io_pipe_phv_in_data_399; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_422 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_400 : io_pipe_phv_in_data_400; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_423 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_401 : io_pipe_phv_in_data_401; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_424 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_402 : io_pipe_phv_in_data_402; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_425 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_403 : io_pipe_phv_in_data_403; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_426 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_404 : io_pipe_phv_in_data_404; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_427 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_405 : io_pipe_phv_in_data_405; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_428 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_406 : io_pipe_phv_in_data_406; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_429 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_407 : io_pipe_phv_in_data_407; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_430 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_408 : io_pipe_phv_in_data_408; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_431 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_409 : io_pipe_phv_in_data_409; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_432 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_410 : io_pipe_phv_in_data_410; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_433 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_411 : io_pipe_phv_in_data_411; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_434 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_412 : io_pipe_phv_in_data_412; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_435 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_413 : io_pipe_phv_in_data_413; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_436 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_414 : io_pipe_phv_in_data_414; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_437 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_415 : io_pipe_phv_in_data_415; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_438 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_416 : io_pipe_phv_in_data_416; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_439 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_417 : io_pipe_phv_in_data_417; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_440 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_418 : io_pipe_phv_in_data_418; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_441 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_419 : io_pipe_phv_in_data_419; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_442 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_420 : io_pipe_phv_in_data_420; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_443 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_421 : io_pipe_phv_in_data_421; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_444 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_422 : io_pipe_phv_in_data_422; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_445 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_423 : io_pipe_phv_in_data_423; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_446 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_424 : io_pipe_phv_in_data_424; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_447 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_425 : io_pipe_phv_in_data_425; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_448 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_426 : io_pipe_phv_in_data_426; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_449 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_427 : io_pipe_phv_in_data_427; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_450 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_428 : io_pipe_phv_in_data_428; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_451 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_429 : io_pipe_phv_in_data_429; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_452 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_430 : io_pipe_phv_in_data_430; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_453 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_431 : io_pipe_phv_in_data_431; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_454 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_432 : io_pipe_phv_in_data_432; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_455 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_433 : io_pipe_phv_in_data_433; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_456 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_434 : io_pipe_phv_in_data_434; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_457 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_435 : io_pipe_phv_in_data_435; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_458 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_436 : io_pipe_phv_in_data_436; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_459 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_437 : io_pipe_phv_in_data_437; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_460 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_438 : io_pipe_phv_in_data_438; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_461 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_439 : io_pipe_phv_in_data_439; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_462 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_440 : io_pipe_phv_in_data_440; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_463 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_441 : io_pipe_phv_in_data_441; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_464 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_442 : io_pipe_phv_in_data_442; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_465 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_443 : io_pipe_phv_in_data_443; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_466 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_444 : io_pipe_phv_in_data_444; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_467 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_445 : io_pipe_phv_in_data_445; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_468 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_446 : io_pipe_phv_in_data_446; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_469 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_447 : io_pipe_phv_in_data_447; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_470 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_448 : io_pipe_phv_in_data_448; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_471 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_449 : io_pipe_phv_in_data_449; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_472 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_450 : io_pipe_phv_in_data_450; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_473 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_451 : io_pipe_phv_in_data_451; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_474 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_452 : io_pipe_phv_in_data_452; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_475 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_453 : io_pipe_phv_in_data_453; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_476 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_454 : io_pipe_phv_in_data_454; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_477 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_455 : io_pipe_phv_in_data_455; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_478 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_456 : io_pipe_phv_in_data_456; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_479 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_457 : io_pipe_phv_in_data_457; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_480 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_458 : io_pipe_phv_in_data_458; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_481 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_459 : io_pipe_phv_in_data_459; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_482 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_460 : io_pipe_phv_in_data_460; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_483 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_461 : io_pipe_phv_in_data_461; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_484 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_462 : io_pipe_phv_in_data_462; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_485 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_463 : io_pipe_phv_in_data_463; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_486 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_464 : io_pipe_phv_in_data_464; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_487 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_465 : io_pipe_phv_in_data_465; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_488 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_466 : io_pipe_phv_in_data_466; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_489 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_467 : io_pipe_phv_in_data_467; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_490 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_468 : io_pipe_phv_in_data_468; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_491 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_469 : io_pipe_phv_in_data_469; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_492 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_470 : io_pipe_phv_in_data_470; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_493 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_471 : io_pipe_phv_in_data_471; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_494 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_472 : io_pipe_phv_in_data_472; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_495 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_473 : io_pipe_phv_in_data_473; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_496 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_474 : io_pipe_phv_in_data_474; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_497 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_475 : io_pipe_phv_in_data_475; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_498 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_476 : io_pipe_phv_in_data_476; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_499 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_477 : io_pipe_phv_in_data_477; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_500 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_478 : io_pipe_phv_in_data_478; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_501 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_479 : io_pipe_phv_in_data_479; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_502 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_480 : io_pipe_phv_in_data_480; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_503 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_481 : io_pipe_phv_in_data_481; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_504 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_482 : io_pipe_phv_in_data_482; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_505 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_483 : io_pipe_phv_in_data_483; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_506 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_484 : io_pipe_phv_in_data_484; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_507 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_485 : io_pipe_phv_in_data_485; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_508 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_486 : io_pipe_phv_in_data_486; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_509 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_487 : io_pipe_phv_in_data_487; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_510 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_488 : io_pipe_phv_in_data_488; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_511 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_489 : io_pipe_phv_in_data_489; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_512 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_490 : io_pipe_phv_in_data_490; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_513 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_491 : io_pipe_phv_in_data_491; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_514 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_492 : io_pipe_phv_in_data_492; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_515 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_493 : io_pipe_phv_in_data_493; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_516 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_494 : io_pipe_phv_in_data_494; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_517 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_495 : io_pipe_phv_in_data_495; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_518 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_496 : io_pipe_phv_in_data_496; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_519 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_497 : io_pipe_phv_in_data_497; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_520 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_498 : io_pipe_phv_in_data_498; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_521 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_499 : io_pipe_phv_in_data_499; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_522 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_500 : io_pipe_phv_in_data_500; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_523 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_501 : io_pipe_phv_in_data_501; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_524 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_502 : io_pipe_phv_in_data_502; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_525 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_503 : io_pipe_phv_in_data_503; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_526 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_504 : io_pipe_phv_in_data_504; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_527 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_505 : io_pipe_phv_in_data_505; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_528 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_506 : io_pipe_phv_in_data_506; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_529 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_507 : io_pipe_phv_in_data_507; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_530 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_508 : io_pipe_phv_in_data_508; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_531 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_509 : io_pipe_phv_in_data_509; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_532 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_510 : io_pipe_phv_in_data_510; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire [7:0] _GEN_533 = 3'h1 == last_mau_id ? mau_1_io_pipe_phv_out_data_511 : io_pipe_phv_in_data_511; // @[parser.scala 33:62 parser.scala 34:35 parser.scala 26:21]
  wire  _GEN_534 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_is_valid_processor : _GEN_0; // @[parser.scala 33:62 parser.scala 34:35]
  wire  _GEN_535 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_config_id : _GEN_1; // @[parser.scala 33:62 parser.scala 34:35]
  wire [3:0] _GEN_536 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_next_processor_id : _GEN_2; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_537 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_parse_transition_field : _GEN_3; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_538 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_parse_current_offset : _GEN_4; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_539 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_parse_current_state : _GEN_5; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_540 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_0 : _GEN_6; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_541 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_1 : _GEN_7; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_542 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_2 : _GEN_8; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_543 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_3 : _GEN_9; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_544 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_4 : _GEN_10; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_545 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_5 : _GEN_11; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_546 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_6 : _GEN_12; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_547 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_7 : _GEN_13; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_548 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_8 : _GEN_14; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_549 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_9 : _GEN_15; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_550 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_10 : _GEN_16; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_551 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_11 : _GEN_17; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_552 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_12 : _GEN_18; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_553 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_13 : _GEN_19; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_554 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_14 : _GEN_20; // @[parser.scala 33:62 parser.scala 34:35]
  wire [15:0] _GEN_555 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_header_15 : _GEN_21; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_556 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_0 : _GEN_22; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_557 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_1 : _GEN_23; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_558 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_2 : _GEN_24; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_559 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_3 : _GEN_25; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_560 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_4 : _GEN_26; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_561 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_5 : _GEN_27; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_562 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_6 : _GEN_28; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_563 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_7 : _GEN_29; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_564 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_8 : _GEN_30; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_565 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_9 : _GEN_31; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_566 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_10 : _GEN_32; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_567 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_11 : _GEN_33; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_568 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_12 : _GEN_34; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_569 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_13 : _GEN_35; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_570 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_14 : _GEN_36; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_571 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_15 : _GEN_37; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_572 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_16 : _GEN_38; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_573 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_17 : _GEN_39; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_574 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_18 : _GEN_40; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_575 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_19 : _GEN_41; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_576 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_20 : _GEN_42; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_577 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_21 : _GEN_43; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_578 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_22 : _GEN_44; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_579 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_23 : _GEN_45; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_580 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_24 : _GEN_46; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_581 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_25 : _GEN_47; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_582 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_26 : _GEN_48; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_583 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_27 : _GEN_49; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_584 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_28 : _GEN_50; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_585 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_29 : _GEN_51; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_586 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_30 : _GEN_52; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_587 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_31 : _GEN_53; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_588 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_32 : _GEN_54; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_589 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_33 : _GEN_55; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_590 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_34 : _GEN_56; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_591 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_35 : _GEN_57; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_592 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_36 : _GEN_58; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_593 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_37 : _GEN_59; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_594 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_38 : _GEN_60; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_595 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_39 : _GEN_61; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_596 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_40 : _GEN_62; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_597 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_41 : _GEN_63; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_598 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_42 : _GEN_64; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_599 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_43 : _GEN_65; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_600 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_44 : _GEN_66; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_601 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_45 : _GEN_67; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_602 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_46 : _GEN_68; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_603 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_47 : _GEN_69; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_604 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_48 : _GEN_70; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_605 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_49 : _GEN_71; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_606 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_50 : _GEN_72; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_607 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_51 : _GEN_73; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_608 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_52 : _GEN_74; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_609 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_53 : _GEN_75; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_610 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_54 : _GEN_76; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_611 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_55 : _GEN_77; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_612 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_56 : _GEN_78; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_613 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_57 : _GEN_79; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_614 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_58 : _GEN_80; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_615 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_59 : _GEN_81; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_616 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_60 : _GEN_82; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_617 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_61 : _GEN_83; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_618 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_62 : _GEN_84; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_619 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_63 : _GEN_85; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_620 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_64 : _GEN_86; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_621 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_65 : _GEN_87; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_622 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_66 : _GEN_88; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_623 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_67 : _GEN_89; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_624 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_68 : _GEN_90; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_625 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_69 : _GEN_91; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_626 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_70 : _GEN_92; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_627 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_71 : _GEN_93; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_628 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_72 : _GEN_94; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_629 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_73 : _GEN_95; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_630 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_74 : _GEN_96; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_631 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_75 : _GEN_97; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_632 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_76 : _GEN_98; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_633 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_77 : _GEN_99; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_634 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_78 : _GEN_100; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_635 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_79 : _GEN_101; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_636 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_80 : _GEN_102; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_637 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_81 : _GEN_103; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_638 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_82 : _GEN_104; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_639 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_83 : _GEN_105; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_640 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_84 : _GEN_106; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_641 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_85 : _GEN_107; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_642 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_86 : _GEN_108; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_643 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_87 : _GEN_109; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_644 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_88 : _GEN_110; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_645 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_89 : _GEN_111; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_646 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_90 : _GEN_112; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_647 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_91 : _GEN_113; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_648 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_92 : _GEN_114; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_649 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_93 : _GEN_115; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_650 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_94 : _GEN_116; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_651 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_95 : _GEN_117; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_652 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_96 : _GEN_118; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_653 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_97 : _GEN_119; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_654 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_98 : _GEN_120; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_655 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_99 : _GEN_121; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_656 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_100 : _GEN_122; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_657 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_101 : _GEN_123; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_658 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_102 : _GEN_124; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_659 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_103 : _GEN_125; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_660 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_104 : _GEN_126; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_661 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_105 : _GEN_127; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_662 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_106 : _GEN_128; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_663 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_107 : _GEN_129; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_664 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_108 : _GEN_130; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_665 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_109 : _GEN_131; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_666 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_110 : _GEN_132; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_667 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_111 : _GEN_133; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_668 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_112 : _GEN_134; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_669 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_113 : _GEN_135; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_670 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_114 : _GEN_136; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_671 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_115 : _GEN_137; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_672 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_116 : _GEN_138; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_673 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_117 : _GEN_139; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_674 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_118 : _GEN_140; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_675 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_119 : _GEN_141; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_676 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_120 : _GEN_142; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_677 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_121 : _GEN_143; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_678 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_122 : _GEN_144; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_679 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_123 : _GEN_145; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_680 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_124 : _GEN_146; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_681 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_125 : _GEN_147; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_682 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_126 : _GEN_148; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_683 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_127 : _GEN_149; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_684 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_128 : _GEN_150; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_685 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_129 : _GEN_151; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_686 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_130 : _GEN_152; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_687 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_131 : _GEN_153; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_688 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_132 : _GEN_154; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_689 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_133 : _GEN_155; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_690 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_134 : _GEN_156; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_691 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_135 : _GEN_157; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_692 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_136 : _GEN_158; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_693 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_137 : _GEN_159; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_694 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_138 : _GEN_160; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_695 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_139 : _GEN_161; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_696 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_140 : _GEN_162; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_697 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_141 : _GEN_163; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_698 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_142 : _GEN_164; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_699 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_143 : _GEN_165; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_700 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_144 : _GEN_166; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_701 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_145 : _GEN_167; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_702 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_146 : _GEN_168; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_703 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_147 : _GEN_169; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_704 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_148 : _GEN_170; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_705 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_149 : _GEN_171; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_706 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_150 : _GEN_172; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_707 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_151 : _GEN_173; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_708 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_152 : _GEN_174; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_709 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_153 : _GEN_175; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_710 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_154 : _GEN_176; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_711 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_155 : _GEN_177; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_712 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_156 : _GEN_178; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_713 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_157 : _GEN_179; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_714 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_158 : _GEN_180; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_715 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_159 : _GEN_181; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_716 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_160 : _GEN_182; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_717 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_161 : _GEN_183; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_718 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_162 : _GEN_184; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_719 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_163 : _GEN_185; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_720 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_164 : _GEN_186; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_721 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_165 : _GEN_187; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_722 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_166 : _GEN_188; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_723 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_167 : _GEN_189; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_724 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_168 : _GEN_190; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_725 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_169 : _GEN_191; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_726 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_170 : _GEN_192; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_727 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_171 : _GEN_193; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_728 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_172 : _GEN_194; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_729 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_173 : _GEN_195; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_730 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_174 : _GEN_196; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_731 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_175 : _GEN_197; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_732 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_176 : _GEN_198; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_733 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_177 : _GEN_199; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_734 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_178 : _GEN_200; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_735 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_179 : _GEN_201; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_736 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_180 : _GEN_202; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_737 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_181 : _GEN_203; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_738 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_182 : _GEN_204; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_739 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_183 : _GEN_205; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_740 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_184 : _GEN_206; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_741 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_185 : _GEN_207; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_742 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_186 : _GEN_208; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_743 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_187 : _GEN_209; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_744 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_188 : _GEN_210; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_745 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_189 : _GEN_211; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_746 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_190 : _GEN_212; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_747 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_191 : _GEN_213; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_748 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_192 : _GEN_214; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_749 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_193 : _GEN_215; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_750 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_194 : _GEN_216; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_751 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_195 : _GEN_217; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_752 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_196 : _GEN_218; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_753 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_197 : _GEN_219; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_754 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_198 : _GEN_220; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_755 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_199 : _GEN_221; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_756 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_200 : _GEN_222; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_757 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_201 : _GEN_223; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_758 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_202 : _GEN_224; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_759 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_203 : _GEN_225; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_760 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_204 : _GEN_226; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_761 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_205 : _GEN_227; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_762 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_206 : _GEN_228; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_763 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_207 : _GEN_229; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_764 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_208 : _GEN_230; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_765 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_209 : _GEN_231; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_766 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_210 : _GEN_232; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_767 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_211 : _GEN_233; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_768 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_212 : _GEN_234; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_769 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_213 : _GEN_235; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_770 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_214 : _GEN_236; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_771 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_215 : _GEN_237; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_772 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_216 : _GEN_238; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_773 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_217 : _GEN_239; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_774 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_218 : _GEN_240; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_775 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_219 : _GEN_241; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_776 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_220 : _GEN_242; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_777 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_221 : _GEN_243; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_778 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_222 : _GEN_244; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_779 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_223 : _GEN_245; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_780 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_224 : _GEN_246; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_781 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_225 : _GEN_247; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_782 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_226 : _GEN_248; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_783 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_227 : _GEN_249; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_784 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_228 : _GEN_250; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_785 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_229 : _GEN_251; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_786 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_230 : _GEN_252; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_787 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_231 : _GEN_253; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_788 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_232 : _GEN_254; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_789 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_233 : _GEN_255; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_790 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_234 : _GEN_256; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_791 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_235 : _GEN_257; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_792 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_236 : _GEN_258; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_793 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_237 : _GEN_259; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_794 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_238 : _GEN_260; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_795 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_239 : _GEN_261; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_796 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_240 : _GEN_262; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_797 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_241 : _GEN_263; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_798 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_242 : _GEN_264; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_799 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_243 : _GEN_265; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_800 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_244 : _GEN_266; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_801 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_245 : _GEN_267; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_802 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_246 : _GEN_268; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_803 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_247 : _GEN_269; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_804 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_248 : _GEN_270; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_805 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_249 : _GEN_271; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_806 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_250 : _GEN_272; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_807 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_251 : _GEN_273; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_808 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_252 : _GEN_274; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_809 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_253 : _GEN_275; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_810 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_254 : _GEN_276; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_811 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_255 : _GEN_277; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_812 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_256 : _GEN_278; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_813 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_257 : _GEN_279; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_814 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_258 : _GEN_280; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_815 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_259 : _GEN_281; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_816 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_260 : _GEN_282; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_817 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_261 : _GEN_283; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_818 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_262 : _GEN_284; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_819 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_263 : _GEN_285; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_820 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_264 : _GEN_286; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_821 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_265 : _GEN_287; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_822 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_266 : _GEN_288; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_823 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_267 : _GEN_289; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_824 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_268 : _GEN_290; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_825 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_269 : _GEN_291; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_826 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_270 : _GEN_292; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_827 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_271 : _GEN_293; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_828 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_272 : _GEN_294; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_829 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_273 : _GEN_295; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_830 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_274 : _GEN_296; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_831 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_275 : _GEN_297; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_832 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_276 : _GEN_298; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_833 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_277 : _GEN_299; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_834 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_278 : _GEN_300; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_835 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_279 : _GEN_301; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_836 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_280 : _GEN_302; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_837 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_281 : _GEN_303; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_838 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_282 : _GEN_304; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_839 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_283 : _GEN_305; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_840 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_284 : _GEN_306; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_841 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_285 : _GEN_307; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_842 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_286 : _GEN_308; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_843 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_287 : _GEN_309; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_844 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_288 : _GEN_310; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_845 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_289 : _GEN_311; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_846 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_290 : _GEN_312; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_847 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_291 : _GEN_313; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_848 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_292 : _GEN_314; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_849 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_293 : _GEN_315; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_850 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_294 : _GEN_316; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_851 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_295 : _GEN_317; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_852 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_296 : _GEN_318; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_853 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_297 : _GEN_319; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_854 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_298 : _GEN_320; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_855 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_299 : _GEN_321; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_856 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_300 : _GEN_322; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_857 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_301 : _GEN_323; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_858 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_302 : _GEN_324; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_859 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_303 : _GEN_325; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_860 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_304 : _GEN_326; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_861 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_305 : _GEN_327; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_862 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_306 : _GEN_328; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_863 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_307 : _GEN_329; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_864 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_308 : _GEN_330; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_865 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_309 : _GEN_331; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_866 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_310 : _GEN_332; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_867 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_311 : _GEN_333; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_868 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_312 : _GEN_334; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_869 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_313 : _GEN_335; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_870 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_314 : _GEN_336; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_871 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_315 : _GEN_337; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_872 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_316 : _GEN_338; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_873 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_317 : _GEN_339; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_874 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_318 : _GEN_340; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_875 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_319 : _GEN_341; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_876 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_320 : _GEN_342; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_877 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_321 : _GEN_343; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_878 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_322 : _GEN_344; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_879 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_323 : _GEN_345; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_880 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_324 : _GEN_346; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_881 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_325 : _GEN_347; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_882 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_326 : _GEN_348; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_883 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_327 : _GEN_349; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_884 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_328 : _GEN_350; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_885 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_329 : _GEN_351; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_886 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_330 : _GEN_352; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_887 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_331 : _GEN_353; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_888 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_332 : _GEN_354; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_889 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_333 : _GEN_355; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_890 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_334 : _GEN_356; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_891 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_335 : _GEN_357; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_892 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_336 : _GEN_358; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_893 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_337 : _GEN_359; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_894 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_338 : _GEN_360; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_895 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_339 : _GEN_361; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_896 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_340 : _GEN_362; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_897 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_341 : _GEN_363; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_898 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_342 : _GEN_364; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_899 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_343 : _GEN_365; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_900 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_344 : _GEN_366; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_901 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_345 : _GEN_367; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_902 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_346 : _GEN_368; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_903 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_347 : _GEN_369; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_904 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_348 : _GEN_370; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_905 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_349 : _GEN_371; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_906 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_350 : _GEN_372; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_907 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_351 : _GEN_373; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_908 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_352 : _GEN_374; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_909 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_353 : _GEN_375; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_910 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_354 : _GEN_376; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_911 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_355 : _GEN_377; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_912 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_356 : _GEN_378; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_913 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_357 : _GEN_379; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_914 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_358 : _GEN_380; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_915 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_359 : _GEN_381; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_916 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_360 : _GEN_382; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_917 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_361 : _GEN_383; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_918 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_362 : _GEN_384; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_919 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_363 : _GEN_385; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_920 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_364 : _GEN_386; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_921 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_365 : _GEN_387; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_922 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_366 : _GEN_388; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_923 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_367 : _GEN_389; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_924 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_368 : _GEN_390; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_925 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_369 : _GEN_391; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_926 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_370 : _GEN_392; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_927 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_371 : _GEN_393; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_928 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_372 : _GEN_394; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_929 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_373 : _GEN_395; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_930 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_374 : _GEN_396; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_931 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_375 : _GEN_397; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_932 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_376 : _GEN_398; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_933 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_377 : _GEN_399; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_934 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_378 : _GEN_400; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_935 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_379 : _GEN_401; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_936 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_380 : _GEN_402; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_937 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_381 : _GEN_403; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_938 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_382 : _GEN_404; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_939 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_383 : _GEN_405; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_940 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_384 : _GEN_406; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_941 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_385 : _GEN_407; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_942 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_386 : _GEN_408; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_943 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_387 : _GEN_409; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_944 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_388 : _GEN_410; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_945 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_389 : _GEN_411; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_946 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_390 : _GEN_412; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_947 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_391 : _GEN_413; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_948 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_392 : _GEN_414; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_949 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_393 : _GEN_415; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_950 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_394 : _GEN_416; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_951 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_395 : _GEN_417; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_952 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_396 : _GEN_418; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_953 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_397 : _GEN_419; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_954 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_398 : _GEN_420; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_955 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_399 : _GEN_421; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_956 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_400 : _GEN_422; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_957 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_401 : _GEN_423; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_958 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_402 : _GEN_424; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_959 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_403 : _GEN_425; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_960 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_404 : _GEN_426; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_961 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_405 : _GEN_427; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_962 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_406 : _GEN_428; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_963 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_407 : _GEN_429; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_964 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_408 : _GEN_430; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_965 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_409 : _GEN_431; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_966 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_410 : _GEN_432; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_967 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_411 : _GEN_433; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_968 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_412 : _GEN_434; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_969 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_413 : _GEN_435; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_970 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_414 : _GEN_436; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_971 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_415 : _GEN_437; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_972 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_416 : _GEN_438; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_973 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_417 : _GEN_439; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_974 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_418 : _GEN_440; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_975 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_419 : _GEN_441; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_976 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_420 : _GEN_442; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_977 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_421 : _GEN_443; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_978 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_422 : _GEN_444; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_979 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_423 : _GEN_445; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_980 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_424 : _GEN_446; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_981 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_425 : _GEN_447; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_982 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_426 : _GEN_448; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_983 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_427 : _GEN_449; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_984 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_428 : _GEN_450; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_985 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_429 : _GEN_451; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_986 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_430 : _GEN_452; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_987 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_431 : _GEN_453; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_988 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_432 : _GEN_454; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_989 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_433 : _GEN_455; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_990 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_434 : _GEN_456; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_991 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_435 : _GEN_457; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_992 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_436 : _GEN_458; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_993 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_437 : _GEN_459; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_994 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_438 : _GEN_460; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_995 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_439 : _GEN_461; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_996 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_440 : _GEN_462; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_997 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_441 : _GEN_463; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_998 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_442 : _GEN_464; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_999 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_443 : _GEN_465; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1000 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_444 : _GEN_466; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1001 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_445 : _GEN_467; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1002 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_446 : _GEN_468; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1003 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_447 : _GEN_469; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1004 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_448 : _GEN_470; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1005 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_449 : _GEN_471; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1006 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_450 : _GEN_472; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1007 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_451 : _GEN_473; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1008 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_452 : _GEN_474; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1009 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_453 : _GEN_475; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1010 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_454 : _GEN_476; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1011 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_455 : _GEN_477; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1012 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_456 : _GEN_478; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1013 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_457 : _GEN_479; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1014 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_458 : _GEN_480; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1015 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_459 : _GEN_481; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1016 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_460 : _GEN_482; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1017 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_461 : _GEN_483; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1018 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_462 : _GEN_484; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1019 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_463 : _GEN_485; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1020 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_464 : _GEN_486; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1021 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_465 : _GEN_487; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1022 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_466 : _GEN_488; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1023 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_467 : _GEN_489; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1024 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_468 : _GEN_490; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1025 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_469 : _GEN_491; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1026 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_470 : _GEN_492; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1027 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_471 : _GEN_493; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1028 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_472 : _GEN_494; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1029 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_473 : _GEN_495; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1030 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_474 : _GEN_496; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1031 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_475 : _GEN_497; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1032 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_476 : _GEN_498; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1033 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_477 : _GEN_499; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1034 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_478 : _GEN_500; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1035 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_479 : _GEN_501; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1036 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_480 : _GEN_502; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1037 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_481 : _GEN_503; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1038 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_482 : _GEN_504; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1039 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_483 : _GEN_505; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1040 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_484 : _GEN_506; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1041 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_485 : _GEN_507; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1042 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_486 : _GEN_508; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1043 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_487 : _GEN_509; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1044 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_488 : _GEN_510; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1045 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_489 : _GEN_511; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1046 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_490 : _GEN_512; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1047 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_491 : _GEN_513; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1048 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_492 : _GEN_514; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1049 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_493 : _GEN_515; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1050 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_494 : _GEN_516; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1051 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_495 : _GEN_517; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1052 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_496 : _GEN_518; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1053 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_497 : _GEN_519; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1054 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_498 : _GEN_520; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1055 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_499 : _GEN_521; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1056 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_500 : _GEN_522; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1057 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_501 : _GEN_523; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1058 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_502 : _GEN_524; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1059 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_503 : _GEN_525; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1060 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_504 : _GEN_526; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1061 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_505 : _GEN_527; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1062 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_506 : _GEN_528; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1063 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_507 : _GEN_529; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1064 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_508 : _GEN_530; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1065 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_509 : _GEN_531; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1066 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_510 : _GEN_532; // @[parser.scala 33:62 parser.scala 34:35]
  wire [7:0] _GEN_1067 = 3'h2 == last_mau_id ? mau_2_io_pipe_phv_out_data_511 : _GEN_533; // @[parser.scala 33:62 parser.scala 34:35]
  wire  mod_j = io_mod_cs == 2'h0; // @[parser.scala 46:35]
  wire  mod_j_1 = io_mod_cs == 2'h1; // @[parser.scala 46:35]
  wire  mod_j_2 = io_mod_cs == 2'h2; // @[parser.scala 46:35]
  wire  mod_j_3 = io_mod_cs == 2'h3; // @[parser.scala 46:35]
  ParseModule mau_0 ( // @[parser.scala 21:25]
    .clock(mau_0_clock),
    .io_pipe_phv_in_data_0(mau_0_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_0_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_0_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_0_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_0_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_0_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_0_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_0_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_0_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_0_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_0_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_0_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_0_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_0_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_0_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_0_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_0_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_0_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_0_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_0_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_0_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_0_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_0_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_0_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_0_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_0_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_0_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_0_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_0_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_0_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_0_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_0_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_0_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_0_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_0_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_0_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_0_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_0_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_0_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_0_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_0_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_0_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_0_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_0_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_0_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_0_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_0_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_0_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_0_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_0_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_0_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_0_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_0_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_0_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_0_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_0_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_0_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_0_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_0_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_0_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_0_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_0_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_0_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_0_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_0_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_0_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_0_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_0_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_0_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_0_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_0_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_0_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_0_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_0_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_0_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_0_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_0_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_0_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_0_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_0_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_0_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_0_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_0_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_0_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_0_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_0_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_0_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_0_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_0_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_0_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_0_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_0_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_0_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_0_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_0_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_0_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_0_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_0_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_0_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_0_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_0_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_0_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_0_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_0_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_0_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_0_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_0_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_0_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_0_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_0_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_0_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_0_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_0_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_0_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_0_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_0_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_0_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_0_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_0_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_0_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_0_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_0_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_0_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_0_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_0_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_0_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_0_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_0_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_0_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_0_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_0_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_0_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_0_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_0_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_0_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_0_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_0_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_0_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_0_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_0_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_0_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_0_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_0_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_0_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_0_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_0_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_0_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_0_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_0_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_0_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_0_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_0_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_0_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_0_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_0_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_0_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_0_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_0_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_0_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_0_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_0_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_0_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_0_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_0_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_0_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_0_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_0_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_0_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_0_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_0_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_0_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_0_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_0_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_0_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_0_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_0_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_0_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_0_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_0_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_0_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_0_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_0_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_0_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_0_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_0_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_0_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_0_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_0_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_0_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_0_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_0_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_0_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_0_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_0_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_0_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_0_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_0_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_0_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_0_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_0_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_0_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_0_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_0_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_0_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_0_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_0_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_0_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_0_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_0_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_0_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_0_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_0_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_0_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_0_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_0_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_0_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_0_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_0_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_0_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_0_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_0_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_0_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_0_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_0_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_0_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_0_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_0_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_0_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_0_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_0_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_0_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_0_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_0_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_0_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_0_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_0_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_0_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_0_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_0_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_0_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_0_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_0_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_0_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_0_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_0_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_0_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_0_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_0_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_0_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_0_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_0_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_0_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_0_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_0_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_0_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_0_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_0_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_0_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_0_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_0_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_0_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_0_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_0_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_0_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_0_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_0_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_0_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_0_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_0_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_0_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_0_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_0_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_0_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_0_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_0_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_0_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_0_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_0_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_0_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_0_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_0_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_0_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_0_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_0_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_0_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_0_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_0_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_0_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_0_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_0_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_0_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_0_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_0_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_0_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_0_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_0_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_0_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_0_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_0_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_0_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_0_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_0_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_0_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_0_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_0_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_0_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_0_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_0_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_0_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_0_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_0_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_0_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_0_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_0_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_0_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_0_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_0_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_0_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_0_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_0_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_0_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_0_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_0_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_0_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_0_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_0_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_0_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_0_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_0_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_0_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_0_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_0_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_0_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_0_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_0_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_0_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_0_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_0_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_0_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_0_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_0_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_0_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_0_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_0_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_0_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_0_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_0_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_0_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_0_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_0_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_0_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_0_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_0_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_0_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_0_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_0_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_0_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_0_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_0_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_0_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_0_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_0_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_0_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_0_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_0_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_0_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_0_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_0_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_0_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_0_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_0_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_0_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_0_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_0_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_0_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_0_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_0_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_0_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_0_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_0_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_0_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_0_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_0_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_0_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_0_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_0_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_0_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_0_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_0_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_0_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_0_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_0_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_0_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_0_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_0_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_0_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_0_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_0_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_0_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_0_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_0_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_0_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_0_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_0_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_0_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_0_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_0_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_0_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_0_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_0_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_0_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_0_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_0_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_0_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_0_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_0_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_0_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_0_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_0_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_0_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_0_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_0_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_0_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_0_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_0_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_0_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_0_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_0_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_0_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_0_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_0_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_0_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_0_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_0_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_0_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_0_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_0_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_0_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_0_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_0_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_0_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_0_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_0_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_0_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_0_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_0_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_0_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_0_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_0_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_0_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_0_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_0_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_0_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_0_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_0_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_0_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_0_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_0_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_0_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_0_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_0_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_0_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_0_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_0_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_0_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_0_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_0_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_0_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_0_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_0_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_0_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_0_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_0_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_0_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_0_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_0_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_0_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_0_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_0_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_0_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_0_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_0_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_0_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_0_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_0_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_0_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_0_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_0_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_0_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_0_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_0_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_0_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_0_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_0_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_0_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_0_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_0_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_0_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_0_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_0_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_0_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_0_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_0_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_0_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_0_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_0_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_0_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_0_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_0_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_0_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_0_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_0_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_0_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_0_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_0_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_0_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_0_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_0_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_0_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_0_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_0_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_0_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_0_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_0_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_0_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_0_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_0_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_0_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_0_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_0_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_0_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_0_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_0_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_0_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_0_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_0_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_0_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_0_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_0_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_0_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_0_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_0_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_0_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_0_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_0_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_0_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_0_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_0_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_0_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_0_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_0_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_0_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_0_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_0_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_0_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_0_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_0_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_0_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_0_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_0_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_0_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_0_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_0_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_0_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_0_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_0_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_0_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_0_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_0_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_0_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_0_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_0_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_0_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_0_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_0_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_0_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_0_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_0_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_0_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_0_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_0_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_0_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_0_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_0_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_0_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_0_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_0_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_0_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_0_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_0_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_0_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_0_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_0_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_0_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_0_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_0_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_0_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_0_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_0_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_0_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_0_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_0_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_0_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_0_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_0_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_0_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_0_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_0_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_0_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_0_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_0_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_0_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_0_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_0_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_0_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_0_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_0_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_0_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_0_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_0_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_0_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_0_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_0_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_0_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_0_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_0_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_0_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_0_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_0_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_0_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_0_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_0_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_0_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_0_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_0_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_0_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_0_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_0_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_0_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_0_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_0_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_0_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_0_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_0_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_0_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_0_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_0_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_0_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_0_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_0_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_0_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_0_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_0_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_0_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_0_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_0_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_0_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_0_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_0_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_0_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_0_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_0_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_0_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_0_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_0_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_0_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_0_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_0_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_0_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_0_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_0_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_0_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_0_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_0_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_0_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_0_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_0_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_0_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_0_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_0_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_0_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_0_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_0_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_0_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_0_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_0_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_0_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_0_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_0_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_0_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_0_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_0_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_0_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_0_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_0_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_0_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_0_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_0_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_0_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_0_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_0_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_0_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_0_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_0_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_0_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_0_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_0_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_0_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_0_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_0_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_0_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_0_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_0_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_0_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_0_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_0_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_0_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_0_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_0_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_0_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_0_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_0_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_0_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_0_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_0_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_0_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_0_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_0_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_0_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_0_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_0_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_0_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_0_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_0_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_0_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_0_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_0_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_0_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_0_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_0_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_0_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_0_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_0_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_0_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_0_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_0_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_0_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_0_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_0_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_0_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_0_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_0_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_0_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_0_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_0_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_0_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_0_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_0_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_0_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_0_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_0_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_0_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_0_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_0_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_0_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_0_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_0_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_0_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_0_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_0_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_0_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_0_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_0_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_0_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_0_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_0_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_0_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_0_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_0_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_0_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_0_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_0_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_0_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_0_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_0_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_0_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_0_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_0_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_0_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_0_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_0_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_0_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_0_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_0_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_0_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_0_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_0_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_0_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_0_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_0_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_0_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_0_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_0_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_0_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_0_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_0_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_0_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_0_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_0_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_0_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_0_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_0_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_0_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_0_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_0_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_0_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_0_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_0_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_0_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_0_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_0_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_0_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_0_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_0_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_0_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_0_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_0_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_0_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_0_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_0_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_0_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_0_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_0_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_0_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_0_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_0_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_0_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_0_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_0_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_0_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_0_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_0_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_0_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_0_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_0_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_0_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_0_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_0_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_0_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_0_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_0_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_0_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_0_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_0_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_0_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_0_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_0_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_0_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_0_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_0_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_0_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_0_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_0_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_0_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_0_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_0_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_0_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_0_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_0_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_0_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_0_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_0_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_0_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_0_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_0_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_0_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_0_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_0_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_0_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_0_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_0_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_0_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_0_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_0_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_0_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_0_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_0_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_0_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_0_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_0_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_0_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_0_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_0_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_0_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_0_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_0_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_0_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_0_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_0_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_0_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_0_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_0_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_0_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_0_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_0_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_0_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_0_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_0_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_0_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_0_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_0_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_0_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_0_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_0_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_0_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_0_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_0_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_0_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_0_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_0_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_0_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_0_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_0_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_0_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_0_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_0_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_0_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_0_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_0_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_0_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_0_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_0_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_0_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_0_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_0_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_0_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_0_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_0_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_0_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_0_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_0_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_0_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_0_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_0_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_0_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_0_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_0_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_0_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_0_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_0_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_0_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_0_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_0_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_0_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_0_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_0_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_0_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_0_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_0_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_0_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_0_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_0_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_0_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_0_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_0_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_0_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_0_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_0_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_0_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_0_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_0_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_0_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_0_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_0_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_0_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_0_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_0_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_0_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_0_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_0_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_0_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_0_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_0_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_0_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_0_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_0_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_0_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_0_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_0_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_0_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_0_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_0_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_0_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_0_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_0_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_0_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_0_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_0_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_0_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_0_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_0_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_0_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_0_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_0_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_0_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_0_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_0_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_0_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_0_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_0_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_0_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_0_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_0_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_0_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_0_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_0_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_0_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_0_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_0_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_0_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_0_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_0_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_0_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_0_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_0_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_0_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_0_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_0_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_0_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_0_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_0_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_0_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_0_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_0_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_0_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_0_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_0_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_0_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_0_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_0_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_0_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_0_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_0_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_0_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_0_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_0_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_0_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_0_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_0_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_0_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_0_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_0_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_0_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_0_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_0_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_0_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_0_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_0_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_0_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_0_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_0_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_0_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_0_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_0_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_0_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_0_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_0_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_0_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_0_io_mod_state_id_mod),
    .io_mod_state_id(mau_0_io_mod_state_id),
    .io_mod_sram_w_cs(mau_0_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_0_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_0_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_0_io_mod_sram_w_data)
  );
  ParseModule mau_1 ( // @[parser.scala 21:25]
    .clock(mau_1_clock),
    .io_pipe_phv_in_data_0(mau_1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_1_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_1_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_1_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_1_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_1_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_1_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_1_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_1_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_1_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_1_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_1_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_1_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_1_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_1_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_1_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_1_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_1_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_1_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_1_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_1_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_1_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_1_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_1_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_1_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_1_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_1_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_1_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_1_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_1_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_1_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_1_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_1_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_1_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_1_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_1_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_1_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_1_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_1_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_1_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_1_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_1_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_1_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_1_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_1_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_1_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_1_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_1_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_1_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_1_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_1_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_1_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_1_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_1_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_1_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_1_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_1_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_1_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_1_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_1_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_1_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_1_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_1_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_1_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_1_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_1_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_1_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_1_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_1_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_1_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_1_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_1_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_1_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_1_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_1_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_1_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_1_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_1_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_1_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_1_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_1_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_1_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_1_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_1_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_1_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_1_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_1_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_1_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_1_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_1_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_1_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_1_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_1_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_1_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_1_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_1_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_1_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_1_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_1_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_1_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_1_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_1_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_1_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_1_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_1_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_1_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_1_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_1_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_1_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_1_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_1_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_1_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_1_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_1_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_1_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_1_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_1_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_1_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_1_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_1_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_1_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_1_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_1_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_1_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_1_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_1_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_1_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_1_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_1_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_1_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_1_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_1_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_1_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_1_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_1_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_1_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_1_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_1_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_1_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_1_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_1_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_1_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_1_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_1_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_1_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_1_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_1_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_1_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_1_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_1_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_1_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_1_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_1_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_1_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_1_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_1_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_1_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_1_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_1_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_1_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_1_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_1_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_1_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_1_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_1_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_1_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_1_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_1_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_1_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_1_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_1_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_1_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_1_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_1_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_1_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_1_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_1_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_1_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_1_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_1_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_1_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_1_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_1_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_1_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_1_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_1_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_1_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_1_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_1_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_1_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_1_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_1_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_1_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_1_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_1_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_1_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_1_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_1_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_1_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_1_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_1_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_1_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_1_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_1_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_1_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_1_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_1_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_1_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_1_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_1_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_1_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_1_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_1_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_1_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_1_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_1_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_1_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_1_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_1_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_1_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_1_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_1_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_1_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_1_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_1_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_1_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_1_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_1_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_1_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_1_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_1_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_1_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_1_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_1_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_1_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_1_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_1_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_1_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_1_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_1_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_1_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_1_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_1_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_1_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_1_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_1_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_1_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_1_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_1_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_1_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_1_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_1_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_1_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_1_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_1_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_1_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_1_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_1_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_1_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_1_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_1_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_1_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_1_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_1_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_1_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_1_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_1_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_1_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_1_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_1_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_1_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_1_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_1_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_1_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_1_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_1_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_1_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_1_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_1_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_1_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_1_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_1_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_1_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_1_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_1_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_1_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_1_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_1_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_1_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_1_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_1_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_1_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_1_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_1_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_1_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_1_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_1_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_1_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_1_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_1_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_1_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_1_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_1_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_1_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_1_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_1_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_1_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_1_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_1_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_1_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_1_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_1_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_1_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_1_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_1_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_1_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_1_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_1_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_1_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_1_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_1_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_1_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_1_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_1_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_1_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_1_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_1_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_1_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_1_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_1_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_1_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_1_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_1_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_1_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_1_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_1_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_1_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_1_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_1_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_1_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_1_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_1_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_1_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_1_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_1_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_1_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_1_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_1_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_1_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_1_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_1_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_1_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_1_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_1_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_1_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_1_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_1_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_1_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_1_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_1_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_1_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_1_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_1_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_1_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_1_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_1_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_1_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_1_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_1_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_1_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_1_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_1_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_1_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_1_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_1_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_1_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_1_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_1_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_1_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_1_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_1_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_1_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_1_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_1_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_1_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_1_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_1_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_1_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_1_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_1_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_1_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_1_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_1_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_1_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_1_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_1_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_1_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_1_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_1_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_1_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_1_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_1_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_1_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_1_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_1_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_1_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_1_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_1_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_1_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_1_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_1_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_1_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_1_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_1_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_1_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_1_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_1_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_1_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_1_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_1_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_1_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_1_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_1_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_1_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_1_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_1_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_1_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_1_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_1_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_1_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_1_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_1_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_1_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_1_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_1_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_1_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_1_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_1_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_1_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_1_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_1_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_1_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_1_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_1_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_1_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_1_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_1_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_1_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_1_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_1_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_1_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_1_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_1_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_1_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_1_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_1_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_1_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_1_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_1_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_1_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_1_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_1_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_1_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_1_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_1_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_1_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_1_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_1_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_1_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_1_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_1_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_1_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_1_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_1_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_1_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_1_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_1_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_1_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_1_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_1_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_1_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_1_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_1_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_1_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_1_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_1_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_1_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_1_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_1_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_1_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_1_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_1_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_1_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_1_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_1_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_1_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_1_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_1_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_1_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_1_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_1_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_1_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_1_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_1_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_1_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_1_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_1_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_1_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_1_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_1_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_1_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_1_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_1_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_1_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_1_io_mod_state_id_mod),
    .io_mod_state_id(mau_1_io_mod_state_id),
    .io_mod_sram_w_cs(mau_1_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_1_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_1_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_1_io_mod_sram_w_data)
  );
  ParseModule mau_2 ( // @[parser.scala 21:25]
    .clock(mau_2_clock),
    .io_pipe_phv_in_data_0(mau_2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_2_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_2_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_2_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_2_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_2_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_2_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_2_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_2_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_2_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_2_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_2_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_2_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_2_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_2_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_2_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_2_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_2_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_2_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_2_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_2_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_2_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_2_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_2_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_2_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_2_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_2_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_2_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_2_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_2_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_2_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_2_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_2_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_2_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_2_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_2_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_2_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_2_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_2_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_2_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_2_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_2_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_2_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_2_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_2_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_2_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_2_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_2_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_2_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_2_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_2_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_2_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_2_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_2_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_2_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_2_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_2_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_2_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_2_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_2_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_2_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_2_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_2_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_2_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_2_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_2_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_2_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_2_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_2_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_2_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_2_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_2_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_2_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_2_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_2_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_2_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_2_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_2_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_2_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_2_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_2_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_2_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_2_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_2_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_2_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_2_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_2_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_2_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_2_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_2_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_2_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_2_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_2_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_2_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_2_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_2_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_2_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_2_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_2_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_2_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_2_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_2_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_2_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_2_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_2_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_2_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_2_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_2_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_2_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_2_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_2_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_2_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_2_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_2_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_2_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_2_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_2_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_2_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_2_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_2_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_2_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_2_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_2_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_2_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_2_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_2_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_2_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_2_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_2_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_2_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_2_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_2_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_2_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_2_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_2_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_2_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_2_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_2_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_2_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_2_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_2_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_2_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_2_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_2_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_2_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_2_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_2_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_2_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_2_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_2_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_2_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_2_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_2_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_2_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_2_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_2_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_2_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_2_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_2_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_2_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_2_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_2_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_2_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_2_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_2_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_2_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_2_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_2_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_2_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_2_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_2_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_2_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_2_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_2_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_2_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_2_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_2_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_2_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_2_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_2_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_2_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_2_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_2_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_2_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_2_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_2_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_2_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_2_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_2_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_2_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_2_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_2_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_2_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_2_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_2_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_2_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_2_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_2_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_2_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_2_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_2_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_2_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_2_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_2_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_2_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_2_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_2_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_2_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_2_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_2_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_2_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_2_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_2_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_2_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_2_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_2_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_2_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_2_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_2_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_2_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_2_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_2_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_2_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_2_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_2_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_2_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_2_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_2_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_2_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_2_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_2_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_2_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_2_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_2_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_2_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_2_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_2_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_2_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_2_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_2_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_2_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_2_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_2_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_2_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_2_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_2_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_2_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_2_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_2_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_2_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_2_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_2_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_2_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_2_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_2_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_2_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_2_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_2_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_2_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_2_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_2_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_2_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_2_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_2_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_2_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_2_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_2_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_2_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_2_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_2_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_2_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_2_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_2_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_2_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_2_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_2_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_2_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_2_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_2_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_2_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_2_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_2_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_2_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_2_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_2_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_2_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_2_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_2_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_2_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_2_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_2_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_2_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_2_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_2_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_2_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_2_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_2_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_2_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_2_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_2_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_2_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_2_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_2_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_2_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_2_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_2_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_2_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_2_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_2_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_2_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_2_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_2_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_2_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_2_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_2_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_2_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_2_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_2_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_2_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_2_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_2_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_2_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_2_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_2_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_2_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_2_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_2_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_2_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_2_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_2_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_2_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_2_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_2_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_2_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_2_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_2_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_2_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_2_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_2_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_2_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_2_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_2_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_2_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_2_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_2_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_2_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_2_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_2_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_2_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_2_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_2_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_2_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_2_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_2_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_2_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_2_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_2_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_2_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_2_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_2_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_2_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_2_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_2_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_2_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_2_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_2_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_2_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_2_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_2_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_2_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_2_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_2_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_2_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_2_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_2_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_2_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_2_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_2_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_2_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_2_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_2_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_2_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_2_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_2_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_2_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_2_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_2_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_2_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_2_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_2_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_2_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_2_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_2_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_2_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_2_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_2_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_2_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_2_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_2_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_2_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_2_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_2_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_2_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_2_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_2_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_2_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_2_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_2_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_2_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_2_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_2_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_2_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_2_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_2_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_2_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_2_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_2_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_2_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_2_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_2_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_2_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_2_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_2_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_2_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_2_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_2_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_2_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_2_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_2_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_2_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_2_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_2_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_2_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_2_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_2_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_2_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_2_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_2_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_2_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_2_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_2_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_2_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_2_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_2_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_2_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_2_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_2_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_2_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_2_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_2_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_2_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_2_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_2_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_2_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_2_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_2_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_2_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_2_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_2_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_2_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_2_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_2_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_2_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_2_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_2_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_2_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_2_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_2_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_2_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_2_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_2_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_2_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_2_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_2_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_2_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_2_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_2_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_2_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_2_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_2_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_2_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_2_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_2_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_2_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_2_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_2_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_2_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_2_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_2_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_2_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_2_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_2_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_2_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_2_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_2_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_2_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_2_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_2_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_2_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_2_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_2_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_2_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_2_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_2_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_2_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_2_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_2_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_2_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_2_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_2_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_2_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_2_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_2_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_2_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_2_io_mod_state_id_mod),
    .io_mod_state_id(mau_2_io_mod_state_id),
    .io_mod_sram_w_cs(mau_2_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_2_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_2_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_2_io_mod_sram_w_data)
  );
  ParseModule mau_3 ( // @[parser.scala 21:25]
    .clock(mau_3_clock),
    .io_pipe_phv_in_data_0(mau_3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(mau_3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(mau_3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(mau_3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(mau_3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(mau_3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(mau_3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(mau_3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(mau_3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(mau_3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(mau_3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(mau_3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(mau_3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(mau_3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(mau_3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(mau_3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(mau_3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(mau_3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(mau_3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(mau_3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(mau_3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(mau_3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(mau_3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(mau_3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(mau_3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(mau_3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(mau_3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(mau_3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(mau_3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(mau_3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(mau_3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(mau_3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(mau_3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(mau_3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(mau_3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(mau_3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(mau_3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(mau_3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(mau_3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(mau_3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(mau_3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(mau_3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(mau_3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(mau_3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(mau_3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(mau_3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(mau_3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(mau_3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(mau_3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(mau_3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(mau_3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(mau_3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(mau_3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(mau_3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(mau_3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(mau_3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(mau_3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(mau_3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(mau_3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(mau_3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(mau_3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(mau_3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(mau_3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(mau_3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(mau_3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(mau_3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(mau_3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(mau_3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(mau_3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(mau_3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(mau_3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(mau_3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(mau_3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(mau_3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(mau_3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(mau_3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(mau_3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(mau_3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(mau_3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(mau_3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(mau_3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(mau_3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(mau_3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(mau_3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(mau_3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(mau_3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(mau_3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(mau_3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(mau_3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(mau_3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(mau_3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(mau_3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(mau_3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(mau_3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(mau_3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(mau_3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(mau_3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(mau_3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(mau_3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(mau_3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(mau_3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(mau_3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(mau_3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(mau_3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(mau_3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(mau_3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(mau_3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(mau_3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(mau_3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(mau_3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(mau_3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(mau_3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(mau_3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(mau_3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(mau_3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(mau_3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(mau_3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(mau_3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(mau_3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(mau_3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(mau_3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(mau_3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(mau_3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(mau_3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(mau_3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(mau_3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(mau_3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(mau_3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(mau_3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(mau_3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(mau_3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(mau_3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(mau_3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(mau_3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(mau_3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(mau_3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(mau_3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(mau_3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(mau_3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(mau_3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(mau_3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(mau_3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(mau_3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(mau_3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(mau_3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(mau_3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(mau_3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(mau_3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(mau_3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(mau_3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(mau_3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(mau_3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(mau_3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(mau_3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(mau_3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(mau_3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(mau_3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(mau_3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(mau_3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(mau_3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(mau_3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(mau_3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(mau_3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(mau_3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(mau_3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(mau_3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(mau_3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(mau_3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(mau_3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(mau_3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(mau_3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(mau_3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(mau_3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(mau_3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(mau_3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(mau_3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(mau_3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(mau_3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(mau_3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(mau_3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(mau_3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(mau_3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(mau_3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(mau_3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(mau_3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(mau_3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(mau_3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(mau_3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(mau_3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(mau_3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(mau_3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(mau_3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(mau_3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(mau_3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(mau_3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(mau_3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(mau_3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(mau_3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(mau_3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(mau_3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(mau_3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(mau_3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(mau_3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(mau_3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(mau_3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(mau_3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(mau_3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(mau_3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(mau_3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(mau_3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(mau_3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(mau_3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(mau_3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(mau_3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(mau_3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(mau_3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(mau_3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(mau_3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(mau_3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(mau_3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(mau_3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(mau_3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(mau_3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(mau_3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(mau_3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(mau_3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(mau_3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(mau_3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(mau_3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(mau_3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(mau_3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(mau_3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(mau_3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(mau_3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(mau_3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(mau_3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(mau_3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(mau_3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(mau_3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(mau_3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(mau_3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(mau_3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(mau_3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(mau_3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(mau_3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(mau_3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(mau_3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(mau_3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(mau_3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(mau_3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(mau_3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(mau_3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(mau_3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(mau_3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(mau_3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(mau_3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(mau_3_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(mau_3_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(mau_3_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(mau_3_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(mau_3_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(mau_3_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(mau_3_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(mau_3_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(mau_3_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(mau_3_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(mau_3_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(mau_3_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(mau_3_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(mau_3_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(mau_3_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(mau_3_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(mau_3_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(mau_3_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(mau_3_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(mau_3_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(mau_3_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(mau_3_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(mau_3_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(mau_3_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(mau_3_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(mau_3_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(mau_3_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(mau_3_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(mau_3_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(mau_3_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(mau_3_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(mau_3_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(mau_3_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(mau_3_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(mau_3_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(mau_3_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(mau_3_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(mau_3_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(mau_3_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(mau_3_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(mau_3_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(mau_3_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(mau_3_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(mau_3_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(mau_3_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(mau_3_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(mau_3_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(mau_3_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(mau_3_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(mau_3_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(mau_3_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(mau_3_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(mau_3_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(mau_3_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(mau_3_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(mau_3_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(mau_3_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(mau_3_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(mau_3_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(mau_3_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(mau_3_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(mau_3_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(mau_3_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(mau_3_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(mau_3_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(mau_3_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(mau_3_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(mau_3_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(mau_3_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(mau_3_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(mau_3_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(mau_3_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(mau_3_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(mau_3_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(mau_3_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(mau_3_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(mau_3_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(mau_3_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(mau_3_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(mau_3_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(mau_3_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(mau_3_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(mau_3_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(mau_3_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(mau_3_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(mau_3_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(mau_3_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(mau_3_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(mau_3_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(mau_3_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(mau_3_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(mau_3_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(mau_3_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(mau_3_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(mau_3_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(mau_3_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(mau_3_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(mau_3_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(mau_3_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(mau_3_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(mau_3_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(mau_3_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(mau_3_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(mau_3_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(mau_3_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(mau_3_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(mau_3_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(mau_3_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(mau_3_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(mau_3_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(mau_3_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(mau_3_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(mau_3_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(mau_3_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(mau_3_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(mau_3_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(mau_3_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(mau_3_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(mau_3_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(mau_3_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(mau_3_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(mau_3_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(mau_3_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(mau_3_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(mau_3_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(mau_3_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(mau_3_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(mau_3_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(mau_3_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(mau_3_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(mau_3_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(mau_3_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(mau_3_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(mau_3_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(mau_3_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(mau_3_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(mau_3_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(mau_3_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(mau_3_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(mau_3_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(mau_3_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(mau_3_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(mau_3_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(mau_3_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(mau_3_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(mau_3_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(mau_3_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(mau_3_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(mau_3_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(mau_3_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(mau_3_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(mau_3_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(mau_3_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(mau_3_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(mau_3_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(mau_3_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(mau_3_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(mau_3_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(mau_3_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(mau_3_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(mau_3_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(mau_3_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(mau_3_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(mau_3_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(mau_3_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(mau_3_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(mau_3_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(mau_3_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(mau_3_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(mau_3_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(mau_3_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(mau_3_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(mau_3_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(mau_3_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(mau_3_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(mau_3_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(mau_3_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(mau_3_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(mau_3_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(mau_3_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(mau_3_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(mau_3_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(mau_3_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(mau_3_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(mau_3_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(mau_3_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(mau_3_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(mau_3_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(mau_3_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(mau_3_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(mau_3_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(mau_3_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(mau_3_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(mau_3_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(mau_3_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(mau_3_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(mau_3_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(mau_3_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(mau_3_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(mau_3_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(mau_3_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(mau_3_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(mau_3_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(mau_3_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(mau_3_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(mau_3_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(mau_3_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(mau_3_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(mau_3_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(mau_3_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(mau_3_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(mau_3_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(mau_3_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(mau_3_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(mau_3_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(mau_3_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(mau_3_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(mau_3_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(mau_3_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(mau_3_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(mau_3_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(mau_3_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(mau_3_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(mau_3_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(mau_3_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(mau_3_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(mau_3_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(mau_3_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(mau_3_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(mau_3_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(mau_3_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(mau_3_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(mau_3_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(mau_3_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(mau_3_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(mau_3_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(mau_3_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(mau_3_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(mau_3_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(mau_3_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(mau_3_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(mau_3_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(mau_3_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(mau_3_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(mau_3_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(mau_3_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(mau_3_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(mau_3_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(mau_3_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(mau_3_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(mau_3_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(mau_3_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(mau_3_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(mau_3_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(mau_3_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(mau_3_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(mau_3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(mau_3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(mau_3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(mau_3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(mau_3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(mau_3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(mau_3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(mau_3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(mau_3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(mau_3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(mau_3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(mau_3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(mau_3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(mau_3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(mau_3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(mau_3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(mau_3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(mau_3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(mau_3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(mau_3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(mau_3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(mau_3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(mau_3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(mau_3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(mau_3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(mau_3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(mau_3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(mau_3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(mau_3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(mau_3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(mau_3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(mau_3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(mau_3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(mau_3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(mau_3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(mau_3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(mau_3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(mau_3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(mau_3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(mau_3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(mau_3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(mau_3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(mau_3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(mau_3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(mau_3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(mau_3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(mau_3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(mau_3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(mau_3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(mau_3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(mau_3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(mau_3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(mau_3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(mau_3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(mau_3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(mau_3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(mau_3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(mau_3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(mau_3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(mau_3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(mau_3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(mau_3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(mau_3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(mau_3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(mau_3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(mau_3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(mau_3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(mau_3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(mau_3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(mau_3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(mau_3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(mau_3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(mau_3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(mau_3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(mau_3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(mau_3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(mau_3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(mau_3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(mau_3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(mau_3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(mau_3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(mau_3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(mau_3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(mau_3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(mau_3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(mau_3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(mau_3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(mau_3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(mau_3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(mau_3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(mau_3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(mau_3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(mau_3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(mau_3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(mau_3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(mau_3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(mau_3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(mau_3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(mau_3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(mau_3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(mau_3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(mau_3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(mau_3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(mau_3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(mau_3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(mau_3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(mau_3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(mau_3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(mau_3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(mau_3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(mau_3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(mau_3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(mau_3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(mau_3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(mau_3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(mau_3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(mau_3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(mau_3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(mau_3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(mau_3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(mau_3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(mau_3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(mau_3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(mau_3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(mau_3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(mau_3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(mau_3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(mau_3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(mau_3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(mau_3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(mau_3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(mau_3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(mau_3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(mau_3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(mau_3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(mau_3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(mau_3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(mau_3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(mau_3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(mau_3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(mau_3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(mau_3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(mau_3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(mau_3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(mau_3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(mau_3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(mau_3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(mau_3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(mau_3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(mau_3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(mau_3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(mau_3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(mau_3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(mau_3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(mau_3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(mau_3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(mau_3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(mau_3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(mau_3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(mau_3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(mau_3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(mau_3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(mau_3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(mau_3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(mau_3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(mau_3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(mau_3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(mau_3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(mau_3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(mau_3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(mau_3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(mau_3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(mau_3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(mau_3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(mau_3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(mau_3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(mau_3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(mau_3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(mau_3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(mau_3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(mau_3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(mau_3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(mau_3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(mau_3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(mau_3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(mau_3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(mau_3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(mau_3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(mau_3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(mau_3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(mau_3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(mau_3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(mau_3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(mau_3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(mau_3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(mau_3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(mau_3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(mau_3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(mau_3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(mau_3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(mau_3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(mau_3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(mau_3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(mau_3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(mau_3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(mau_3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(mau_3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(mau_3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(mau_3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(mau_3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(mau_3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(mau_3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(mau_3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(mau_3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(mau_3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(mau_3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(mau_3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(mau_3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(mau_3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(mau_3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(mau_3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(mau_3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(mau_3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(mau_3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(mau_3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(mau_3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(mau_3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(mau_3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(mau_3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(mau_3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(mau_3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(mau_3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(mau_3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(mau_3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(mau_3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(mau_3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(mau_3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(mau_3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(mau_3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(mau_3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(mau_3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(mau_3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(mau_3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(mau_3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(mau_3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(mau_3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(mau_3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(mau_3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(mau_3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(mau_3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(mau_3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(mau_3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(mau_3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(mau_3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(mau_3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(mau_3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(mau_3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(mau_3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(mau_3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(mau_3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(mau_3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(mau_3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(mau_3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(mau_3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(mau_3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(mau_3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(mau_3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(mau_3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(mau_3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(mau_3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(mau_3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(mau_3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(mau_3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(mau_3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(mau_3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(mau_3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(mau_3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(mau_3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(mau_3_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(mau_3_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(mau_3_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(mau_3_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(mau_3_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(mau_3_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(mau_3_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(mau_3_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(mau_3_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(mau_3_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(mau_3_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(mau_3_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(mau_3_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(mau_3_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(mau_3_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(mau_3_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(mau_3_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(mau_3_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(mau_3_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(mau_3_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(mau_3_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(mau_3_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(mau_3_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(mau_3_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(mau_3_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(mau_3_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(mau_3_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(mau_3_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(mau_3_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(mau_3_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(mau_3_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(mau_3_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(mau_3_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(mau_3_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(mau_3_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(mau_3_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(mau_3_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(mau_3_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(mau_3_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(mau_3_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(mau_3_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(mau_3_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(mau_3_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(mau_3_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(mau_3_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(mau_3_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(mau_3_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(mau_3_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(mau_3_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(mau_3_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(mau_3_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(mau_3_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(mau_3_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(mau_3_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(mau_3_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(mau_3_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(mau_3_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(mau_3_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(mau_3_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(mau_3_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(mau_3_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(mau_3_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(mau_3_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(mau_3_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(mau_3_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(mau_3_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(mau_3_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(mau_3_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(mau_3_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(mau_3_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(mau_3_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(mau_3_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(mau_3_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(mau_3_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(mau_3_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(mau_3_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(mau_3_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(mau_3_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(mau_3_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(mau_3_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(mau_3_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(mau_3_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(mau_3_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(mau_3_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(mau_3_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(mau_3_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(mau_3_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(mau_3_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(mau_3_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(mau_3_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(mau_3_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(mau_3_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(mau_3_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(mau_3_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(mau_3_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(mau_3_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(mau_3_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(mau_3_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(mau_3_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(mau_3_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(mau_3_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(mau_3_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(mau_3_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(mau_3_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(mau_3_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(mau_3_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(mau_3_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(mau_3_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(mau_3_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(mau_3_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(mau_3_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(mau_3_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(mau_3_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(mau_3_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(mau_3_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(mau_3_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(mau_3_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(mau_3_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(mau_3_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(mau_3_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(mau_3_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(mau_3_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(mau_3_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(mau_3_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(mau_3_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(mau_3_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(mau_3_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(mau_3_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(mau_3_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(mau_3_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(mau_3_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(mau_3_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(mau_3_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(mau_3_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(mau_3_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(mau_3_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(mau_3_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(mau_3_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(mau_3_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(mau_3_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(mau_3_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(mau_3_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(mau_3_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(mau_3_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(mau_3_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(mau_3_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(mau_3_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(mau_3_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(mau_3_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(mau_3_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(mau_3_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(mau_3_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(mau_3_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(mau_3_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(mau_3_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(mau_3_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(mau_3_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(mau_3_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(mau_3_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(mau_3_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(mau_3_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(mau_3_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(mau_3_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(mau_3_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(mau_3_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(mau_3_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(mau_3_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(mau_3_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(mau_3_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(mau_3_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(mau_3_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(mau_3_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(mau_3_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(mau_3_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(mau_3_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(mau_3_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(mau_3_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(mau_3_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(mau_3_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(mau_3_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(mau_3_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(mau_3_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(mau_3_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(mau_3_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(mau_3_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(mau_3_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(mau_3_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(mau_3_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(mau_3_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(mau_3_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(mau_3_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(mau_3_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(mau_3_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(mau_3_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(mau_3_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(mau_3_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(mau_3_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(mau_3_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(mau_3_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(mau_3_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(mau_3_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(mau_3_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(mau_3_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(mau_3_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(mau_3_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(mau_3_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(mau_3_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(mau_3_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(mau_3_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(mau_3_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(mau_3_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(mau_3_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(mau_3_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(mau_3_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(mau_3_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(mau_3_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(mau_3_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(mau_3_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(mau_3_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(mau_3_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(mau_3_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(mau_3_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(mau_3_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(mau_3_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(mau_3_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(mau_3_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(mau_3_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(mau_3_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(mau_3_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(mau_3_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(mau_3_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(mau_3_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(mau_3_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(mau_3_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(mau_3_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(mau_3_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(mau_3_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(mau_3_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(mau_3_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(mau_3_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(mau_3_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(mau_3_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(mau_3_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(mau_3_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(mau_3_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(mau_3_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(mau_3_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(mau_3_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(mau_3_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(mau_3_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(mau_3_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(mau_3_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(mau_3_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(mau_3_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(mau_3_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(mau_3_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(mau_3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(mau_3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(mau_3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(mau_3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(mau_3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(mau_3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(mau_3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(mau_3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(mau_3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(mau_3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(mau_3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(mau_3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(mau_3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(mau_3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(mau_3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(mau_3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(mau_3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(mau_3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(mau_3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(mau_3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(mau_3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(mau_3_io_pipe_phv_out_is_valid_processor),
    .io_mod_state_id_mod(mau_3_io_mod_state_id_mod),
    .io_mod_state_id(mau_3_io_mod_state_id),
    .io_mod_sram_w_cs(mau_3_io_mod_sram_w_cs),
    .io_mod_sram_w_en(mau_3_io_mod_sram_w_en),
    .io_mod_sram_w_addr(mau_3_io_mod_sram_w_addr),
    .io_mod_sram_w_data(mau_3_io_mod_sram_w_data)
  );
  assign io_pipe_phv_out_data_0 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_0 : _GEN_556; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_1 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_1 : _GEN_557; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_2 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_2 : _GEN_558; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_3 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_3 : _GEN_559; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_4 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_4 : _GEN_560; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_5 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_5 : _GEN_561; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_6 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_6 : _GEN_562; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_7 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_7 : _GEN_563; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_8 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_8 : _GEN_564; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_9 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_9 : _GEN_565; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_10 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_10 : _GEN_566; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_11 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_11 : _GEN_567; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_12 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_12 : _GEN_568; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_13 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_13 : _GEN_569; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_14 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_14 : _GEN_570; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_15 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_15 : _GEN_571; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_16 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_16 : _GEN_572; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_17 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_17 : _GEN_573; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_18 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_18 : _GEN_574; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_19 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_19 : _GEN_575; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_20 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_20 : _GEN_576; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_21 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_21 : _GEN_577; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_22 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_22 : _GEN_578; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_23 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_23 : _GEN_579; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_24 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_24 : _GEN_580; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_25 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_25 : _GEN_581; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_26 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_26 : _GEN_582; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_27 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_27 : _GEN_583; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_28 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_28 : _GEN_584; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_29 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_29 : _GEN_585; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_30 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_30 : _GEN_586; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_31 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_31 : _GEN_587; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_32 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_32 : _GEN_588; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_33 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_33 : _GEN_589; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_34 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_34 : _GEN_590; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_35 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_35 : _GEN_591; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_36 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_36 : _GEN_592; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_37 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_37 : _GEN_593; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_38 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_38 : _GEN_594; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_39 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_39 : _GEN_595; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_40 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_40 : _GEN_596; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_41 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_41 : _GEN_597; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_42 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_42 : _GEN_598; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_43 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_43 : _GEN_599; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_44 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_44 : _GEN_600; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_45 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_45 : _GEN_601; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_46 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_46 : _GEN_602; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_47 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_47 : _GEN_603; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_48 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_48 : _GEN_604; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_49 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_49 : _GEN_605; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_50 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_50 : _GEN_606; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_51 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_51 : _GEN_607; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_52 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_52 : _GEN_608; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_53 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_53 : _GEN_609; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_54 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_54 : _GEN_610; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_55 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_55 : _GEN_611; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_56 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_56 : _GEN_612; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_57 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_57 : _GEN_613; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_58 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_58 : _GEN_614; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_59 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_59 : _GEN_615; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_60 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_60 : _GEN_616; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_61 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_61 : _GEN_617; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_62 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_62 : _GEN_618; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_63 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_63 : _GEN_619; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_64 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_64 : _GEN_620; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_65 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_65 : _GEN_621; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_66 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_66 : _GEN_622; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_67 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_67 : _GEN_623; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_68 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_68 : _GEN_624; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_69 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_69 : _GEN_625; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_70 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_70 : _GEN_626; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_71 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_71 : _GEN_627; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_72 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_72 : _GEN_628; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_73 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_73 : _GEN_629; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_74 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_74 : _GEN_630; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_75 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_75 : _GEN_631; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_76 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_76 : _GEN_632; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_77 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_77 : _GEN_633; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_78 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_78 : _GEN_634; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_79 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_79 : _GEN_635; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_80 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_80 : _GEN_636; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_81 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_81 : _GEN_637; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_82 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_82 : _GEN_638; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_83 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_83 : _GEN_639; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_84 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_84 : _GEN_640; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_85 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_85 : _GEN_641; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_86 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_86 : _GEN_642; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_87 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_87 : _GEN_643; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_88 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_88 : _GEN_644; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_89 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_89 : _GEN_645; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_90 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_90 : _GEN_646; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_91 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_91 : _GEN_647; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_92 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_92 : _GEN_648; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_93 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_93 : _GEN_649; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_94 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_94 : _GEN_650; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_95 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_95 : _GEN_651; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_96 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_96 : _GEN_652; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_97 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_97 : _GEN_653; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_98 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_98 : _GEN_654; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_99 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_99 : _GEN_655; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_100 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_100 : _GEN_656; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_101 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_101 : _GEN_657; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_102 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_102 : _GEN_658; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_103 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_103 : _GEN_659; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_104 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_104 : _GEN_660; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_105 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_105 : _GEN_661; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_106 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_106 : _GEN_662; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_107 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_107 : _GEN_663; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_108 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_108 : _GEN_664; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_109 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_109 : _GEN_665; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_110 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_110 : _GEN_666; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_111 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_111 : _GEN_667; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_112 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_112 : _GEN_668; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_113 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_113 : _GEN_669; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_114 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_114 : _GEN_670; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_115 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_115 : _GEN_671; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_116 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_116 : _GEN_672; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_117 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_117 : _GEN_673; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_118 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_118 : _GEN_674; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_119 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_119 : _GEN_675; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_120 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_120 : _GEN_676; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_121 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_121 : _GEN_677; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_122 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_122 : _GEN_678; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_123 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_123 : _GEN_679; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_124 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_124 : _GEN_680; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_125 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_125 : _GEN_681; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_126 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_126 : _GEN_682; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_127 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_127 : _GEN_683; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_128 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_128 : _GEN_684; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_129 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_129 : _GEN_685; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_130 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_130 : _GEN_686; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_131 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_131 : _GEN_687; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_132 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_132 : _GEN_688; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_133 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_133 : _GEN_689; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_134 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_134 : _GEN_690; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_135 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_135 : _GEN_691; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_136 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_136 : _GEN_692; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_137 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_137 : _GEN_693; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_138 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_138 : _GEN_694; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_139 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_139 : _GEN_695; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_140 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_140 : _GEN_696; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_141 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_141 : _GEN_697; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_142 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_142 : _GEN_698; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_143 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_143 : _GEN_699; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_144 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_144 : _GEN_700; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_145 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_145 : _GEN_701; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_146 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_146 : _GEN_702; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_147 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_147 : _GEN_703; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_148 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_148 : _GEN_704; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_149 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_149 : _GEN_705; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_150 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_150 : _GEN_706; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_151 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_151 : _GEN_707; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_152 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_152 : _GEN_708; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_153 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_153 : _GEN_709; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_154 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_154 : _GEN_710; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_155 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_155 : _GEN_711; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_156 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_156 : _GEN_712; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_157 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_157 : _GEN_713; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_158 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_158 : _GEN_714; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_159 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_159 : _GEN_715; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_160 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_160 : _GEN_716; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_161 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_161 : _GEN_717; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_162 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_162 : _GEN_718; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_163 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_163 : _GEN_719; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_164 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_164 : _GEN_720; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_165 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_165 : _GEN_721; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_166 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_166 : _GEN_722; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_167 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_167 : _GEN_723; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_168 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_168 : _GEN_724; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_169 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_169 : _GEN_725; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_170 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_170 : _GEN_726; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_171 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_171 : _GEN_727; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_172 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_172 : _GEN_728; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_173 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_173 : _GEN_729; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_174 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_174 : _GEN_730; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_175 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_175 : _GEN_731; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_176 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_176 : _GEN_732; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_177 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_177 : _GEN_733; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_178 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_178 : _GEN_734; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_179 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_179 : _GEN_735; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_180 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_180 : _GEN_736; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_181 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_181 : _GEN_737; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_182 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_182 : _GEN_738; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_183 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_183 : _GEN_739; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_184 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_184 : _GEN_740; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_185 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_185 : _GEN_741; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_186 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_186 : _GEN_742; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_187 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_187 : _GEN_743; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_188 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_188 : _GEN_744; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_189 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_189 : _GEN_745; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_190 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_190 : _GEN_746; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_191 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_191 : _GEN_747; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_192 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_192 : _GEN_748; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_193 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_193 : _GEN_749; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_194 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_194 : _GEN_750; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_195 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_195 : _GEN_751; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_196 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_196 : _GEN_752; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_197 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_197 : _GEN_753; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_198 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_198 : _GEN_754; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_199 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_199 : _GEN_755; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_200 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_200 : _GEN_756; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_201 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_201 : _GEN_757; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_202 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_202 : _GEN_758; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_203 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_203 : _GEN_759; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_204 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_204 : _GEN_760; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_205 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_205 : _GEN_761; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_206 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_206 : _GEN_762; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_207 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_207 : _GEN_763; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_208 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_208 : _GEN_764; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_209 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_209 : _GEN_765; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_210 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_210 : _GEN_766; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_211 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_211 : _GEN_767; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_212 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_212 : _GEN_768; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_213 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_213 : _GEN_769; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_214 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_214 : _GEN_770; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_215 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_215 : _GEN_771; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_216 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_216 : _GEN_772; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_217 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_217 : _GEN_773; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_218 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_218 : _GEN_774; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_219 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_219 : _GEN_775; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_220 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_220 : _GEN_776; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_221 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_221 : _GEN_777; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_222 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_222 : _GEN_778; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_223 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_223 : _GEN_779; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_224 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_224 : _GEN_780; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_225 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_225 : _GEN_781; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_226 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_226 : _GEN_782; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_227 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_227 : _GEN_783; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_228 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_228 : _GEN_784; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_229 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_229 : _GEN_785; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_230 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_230 : _GEN_786; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_231 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_231 : _GEN_787; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_232 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_232 : _GEN_788; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_233 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_233 : _GEN_789; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_234 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_234 : _GEN_790; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_235 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_235 : _GEN_791; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_236 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_236 : _GEN_792; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_237 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_237 : _GEN_793; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_238 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_238 : _GEN_794; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_239 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_239 : _GEN_795; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_240 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_240 : _GEN_796; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_241 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_241 : _GEN_797; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_242 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_242 : _GEN_798; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_243 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_243 : _GEN_799; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_244 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_244 : _GEN_800; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_245 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_245 : _GEN_801; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_246 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_246 : _GEN_802; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_247 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_247 : _GEN_803; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_248 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_248 : _GEN_804; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_249 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_249 : _GEN_805; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_250 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_250 : _GEN_806; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_251 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_251 : _GEN_807; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_252 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_252 : _GEN_808; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_253 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_253 : _GEN_809; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_254 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_254 : _GEN_810; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_255 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_255 : _GEN_811; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_256 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_256 : _GEN_812; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_257 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_257 : _GEN_813; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_258 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_258 : _GEN_814; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_259 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_259 : _GEN_815; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_260 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_260 : _GEN_816; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_261 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_261 : _GEN_817; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_262 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_262 : _GEN_818; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_263 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_263 : _GEN_819; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_264 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_264 : _GEN_820; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_265 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_265 : _GEN_821; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_266 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_266 : _GEN_822; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_267 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_267 : _GEN_823; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_268 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_268 : _GEN_824; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_269 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_269 : _GEN_825; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_270 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_270 : _GEN_826; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_271 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_271 : _GEN_827; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_272 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_272 : _GEN_828; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_273 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_273 : _GEN_829; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_274 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_274 : _GEN_830; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_275 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_275 : _GEN_831; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_276 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_276 : _GEN_832; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_277 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_277 : _GEN_833; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_278 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_278 : _GEN_834; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_279 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_279 : _GEN_835; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_280 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_280 : _GEN_836; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_281 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_281 : _GEN_837; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_282 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_282 : _GEN_838; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_283 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_283 : _GEN_839; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_284 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_284 : _GEN_840; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_285 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_285 : _GEN_841; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_286 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_286 : _GEN_842; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_287 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_287 : _GEN_843; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_288 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_288 : _GEN_844; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_289 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_289 : _GEN_845; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_290 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_290 : _GEN_846; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_291 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_291 : _GEN_847; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_292 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_292 : _GEN_848; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_293 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_293 : _GEN_849; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_294 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_294 : _GEN_850; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_295 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_295 : _GEN_851; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_296 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_296 : _GEN_852; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_297 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_297 : _GEN_853; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_298 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_298 : _GEN_854; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_299 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_299 : _GEN_855; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_300 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_300 : _GEN_856; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_301 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_301 : _GEN_857; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_302 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_302 : _GEN_858; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_303 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_303 : _GEN_859; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_304 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_304 : _GEN_860; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_305 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_305 : _GEN_861; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_306 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_306 : _GEN_862; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_307 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_307 : _GEN_863; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_308 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_308 : _GEN_864; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_309 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_309 : _GEN_865; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_310 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_310 : _GEN_866; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_311 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_311 : _GEN_867; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_312 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_312 : _GEN_868; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_313 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_313 : _GEN_869; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_314 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_314 : _GEN_870; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_315 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_315 : _GEN_871; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_316 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_316 : _GEN_872; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_317 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_317 : _GEN_873; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_318 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_318 : _GEN_874; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_319 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_319 : _GEN_875; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_320 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_320 : _GEN_876; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_321 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_321 : _GEN_877; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_322 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_322 : _GEN_878; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_323 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_323 : _GEN_879; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_324 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_324 : _GEN_880; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_325 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_325 : _GEN_881; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_326 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_326 : _GEN_882; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_327 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_327 : _GEN_883; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_328 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_328 : _GEN_884; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_329 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_329 : _GEN_885; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_330 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_330 : _GEN_886; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_331 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_331 : _GEN_887; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_332 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_332 : _GEN_888; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_333 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_333 : _GEN_889; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_334 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_334 : _GEN_890; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_335 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_335 : _GEN_891; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_336 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_336 : _GEN_892; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_337 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_337 : _GEN_893; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_338 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_338 : _GEN_894; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_339 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_339 : _GEN_895; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_340 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_340 : _GEN_896; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_341 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_341 : _GEN_897; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_342 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_342 : _GEN_898; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_343 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_343 : _GEN_899; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_344 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_344 : _GEN_900; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_345 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_345 : _GEN_901; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_346 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_346 : _GEN_902; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_347 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_347 : _GEN_903; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_348 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_348 : _GEN_904; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_349 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_349 : _GEN_905; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_350 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_350 : _GEN_906; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_351 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_351 : _GEN_907; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_352 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_352 : _GEN_908; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_353 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_353 : _GEN_909; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_354 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_354 : _GEN_910; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_355 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_355 : _GEN_911; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_356 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_356 : _GEN_912; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_357 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_357 : _GEN_913; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_358 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_358 : _GEN_914; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_359 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_359 : _GEN_915; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_360 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_360 : _GEN_916; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_361 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_361 : _GEN_917; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_362 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_362 : _GEN_918; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_363 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_363 : _GEN_919; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_364 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_364 : _GEN_920; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_365 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_365 : _GEN_921; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_366 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_366 : _GEN_922; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_367 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_367 : _GEN_923; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_368 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_368 : _GEN_924; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_369 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_369 : _GEN_925; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_370 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_370 : _GEN_926; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_371 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_371 : _GEN_927; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_372 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_372 : _GEN_928; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_373 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_373 : _GEN_929; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_374 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_374 : _GEN_930; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_375 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_375 : _GEN_931; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_376 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_376 : _GEN_932; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_377 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_377 : _GEN_933; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_378 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_378 : _GEN_934; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_379 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_379 : _GEN_935; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_380 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_380 : _GEN_936; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_381 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_381 : _GEN_937; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_382 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_382 : _GEN_938; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_383 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_383 : _GEN_939; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_384 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_384 : _GEN_940; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_385 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_385 : _GEN_941; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_386 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_386 : _GEN_942; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_387 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_387 : _GEN_943; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_388 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_388 : _GEN_944; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_389 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_389 : _GEN_945; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_390 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_390 : _GEN_946; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_391 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_391 : _GEN_947; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_392 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_392 : _GEN_948; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_393 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_393 : _GEN_949; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_394 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_394 : _GEN_950; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_395 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_395 : _GEN_951; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_396 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_396 : _GEN_952; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_397 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_397 : _GEN_953; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_398 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_398 : _GEN_954; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_399 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_399 : _GEN_955; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_400 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_400 : _GEN_956; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_401 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_401 : _GEN_957; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_402 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_402 : _GEN_958; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_403 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_403 : _GEN_959; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_404 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_404 : _GEN_960; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_405 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_405 : _GEN_961; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_406 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_406 : _GEN_962; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_407 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_407 : _GEN_963; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_408 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_408 : _GEN_964; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_409 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_409 : _GEN_965; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_410 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_410 : _GEN_966; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_411 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_411 : _GEN_967; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_412 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_412 : _GEN_968; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_413 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_413 : _GEN_969; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_414 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_414 : _GEN_970; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_415 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_415 : _GEN_971; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_416 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_416 : _GEN_972; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_417 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_417 : _GEN_973; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_418 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_418 : _GEN_974; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_419 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_419 : _GEN_975; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_420 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_420 : _GEN_976; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_421 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_421 : _GEN_977; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_422 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_422 : _GEN_978; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_423 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_423 : _GEN_979; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_424 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_424 : _GEN_980; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_425 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_425 : _GEN_981; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_426 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_426 : _GEN_982; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_427 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_427 : _GEN_983; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_428 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_428 : _GEN_984; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_429 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_429 : _GEN_985; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_430 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_430 : _GEN_986; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_431 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_431 : _GEN_987; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_432 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_432 : _GEN_988; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_433 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_433 : _GEN_989; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_434 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_434 : _GEN_990; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_435 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_435 : _GEN_991; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_436 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_436 : _GEN_992; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_437 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_437 : _GEN_993; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_438 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_438 : _GEN_994; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_439 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_439 : _GEN_995; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_440 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_440 : _GEN_996; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_441 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_441 : _GEN_997; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_442 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_442 : _GEN_998; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_443 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_443 : _GEN_999; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_444 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_444 : _GEN_1000; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_445 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_445 : _GEN_1001; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_446 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_446 : _GEN_1002; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_447 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_447 : _GEN_1003; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_448 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_448 : _GEN_1004; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_449 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_449 : _GEN_1005; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_450 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_450 : _GEN_1006; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_451 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_451 : _GEN_1007; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_452 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_452 : _GEN_1008; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_453 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_453 : _GEN_1009; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_454 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_454 : _GEN_1010; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_455 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_455 : _GEN_1011; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_456 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_456 : _GEN_1012; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_457 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_457 : _GEN_1013; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_458 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_458 : _GEN_1014; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_459 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_459 : _GEN_1015; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_460 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_460 : _GEN_1016; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_461 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_461 : _GEN_1017; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_462 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_462 : _GEN_1018; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_463 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_463 : _GEN_1019; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_464 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_464 : _GEN_1020; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_465 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_465 : _GEN_1021; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_466 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_466 : _GEN_1022; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_467 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_467 : _GEN_1023; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_468 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_468 : _GEN_1024; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_469 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_469 : _GEN_1025; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_470 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_470 : _GEN_1026; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_471 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_471 : _GEN_1027; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_472 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_472 : _GEN_1028; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_473 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_473 : _GEN_1029; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_474 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_474 : _GEN_1030; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_475 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_475 : _GEN_1031; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_476 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_476 : _GEN_1032; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_477 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_477 : _GEN_1033; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_478 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_478 : _GEN_1034; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_479 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_479 : _GEN_1035; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_480 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_480 : _GEN_1036; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_481 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_481 : _GEN_1037; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_482 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_482 : _GEN_1038; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_483 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_483 : _GEN_1039; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_484 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_484 : _GEN_1040; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_485 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_485 : _GEN_1041; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_486 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_486 : _GEN_1042; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_487 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_487 : _GEN_1043; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_488 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_488 : _GEN_1044; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_489 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_489 : _GEN_1045; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_490 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_490 : _GEN_1046; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_491 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_491 : _GEN_1047; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_492 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_492 : _GEN_1048; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_493 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_493 : _GEN_1049; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_494 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_494 : _GEN_1050; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_495 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_495 : _GEN_1051; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_496 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_496 : _GEN_1052; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_497 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_497 : _GEN_1053; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_498 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_498 : _GEN_1054; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_499 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_499 : _GEN_1055; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_500 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_500 : _GEN_1056; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_501 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_501 : _GEN_1057; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_502 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_502 : _GEN_1058; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_503 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_503 : _GEN_1059; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_504 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_504 : _GEN_1060; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_505 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_505 : _GEN_1061; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_506 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_506 : _GEN_1062; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_507 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_507 : _GEN_1063; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_508 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_508 : _GEN_1064; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_509 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_509 : _GEN_1065; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_510 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_510 : _GEN_1066; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_data_511 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_data_511 : _GEN_1067; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_0 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_0 : _GEN_540; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_1 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_1 : _GEN_541; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_2 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_2 : _GEN_542; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_3 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_3 : _GEN_543; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_4 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_4 : _GEN_544; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_5 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_5 : _GEN_545; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_6 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_6 : _GEN_546; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_7 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_7 : _GEN_547; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_8 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_8 : _GEN_548; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_9 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_9 : _GEN_549; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_10 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_10 : _GEN_550; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_11 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_11 : _GEN_551; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_12 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_12 : _GEN_552; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_13 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_13 : _GEN_553; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_14 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_14 : _GEN_554; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_header_15 = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_header_15 : _GEN_555; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_current_state = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_parse_current_state :
    _GEN_539; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_current_offset = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_parse_current_offset :
    _GEN_538; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_parse_transition_field = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_parse_transition_field :
    _GEN_537; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_next_processor_id = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_processor_id : _GEN_536; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_next_config_id = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_next_config_id : _GEN_535; // @[parser.scala 33:62 parser.scala 34:35]
  assign io_pipe_phv_out_is_valid_processor = 3'h3 == last_mau_id ? mau_3_io_pipe_phv_out_is_valid_processor : _GEN_534; // @[parser.scala 33:62 parser.scala 34:35]
  assign mau_0_clock = clock;
  assign mau_0_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_256 = io_pipe_phv_in_data_256; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_257 = io_pipe_phv_in_data_257; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_258 = io_pipe_phv_in_data_258; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_259 = io_pipe_phv_in_data_259; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_260 = io_pipe_phv_in_data_260; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_261 = io_pipe_phv_in_data_261; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_262 = io_pipe_phv_in_data_262; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_263 = io_pipe_phv_in_data_263; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_264 = io_pipe_phv_in_data_264; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_265 = io_pipe_phv_in_data_265; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_266 = io_pipe_phv_in_data_266; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_267 = io_pipe_phv_in_data_267; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_268 = io_pipe_phv_in_data_268; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_269 = io_pipe_phv_in_data_269; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_270 = io_pipe_phv_in_data_270; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_271 = io_pipe_phv_in_data_271; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_272 = io_pipe_phv_in_data_272; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_273 = io_pipe_phv_in_data_273; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_274 = io_pipe_phv_in_data_274; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_275 = io_pipe_phv_in_data_275; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_276 = io_pipe_phv_in_data_276; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_277 = io_pipe_phv_in_data_277; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_278 = io_pipe_phv_in_data_278; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_279 = io_pipe_phv_in_data_279; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_280 = io_pipe_phv_in_data_280; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_281 = io_pipe_phv_in_data_281; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_282 = io_pipe_phv_in_data_282; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_283 = io_pipe_phv_in_data_283; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_284 = io_pipe_phv_in_data_284; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_285 = io_pipe_phv_in_data_285; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_286 = io_pipe_phv_in_data_286; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_287 = io_pipe_phv_in_data_287; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_288 = io_pipe_phv_in_data_288; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_289 = io_pipe_phv_in_data_289; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_290 = io_pipe_phv_in_data_290; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_291 = io_pipe_phv_in_data_291; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_292 = io_pipe_phv_in_data_292; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_293 = io_pipe_phv_in_data_293; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_294 = io_pipe_phv_in_data_294; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_295 = io_pipe_phv_in_data_295; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_296 = io_pipe_phv_in_data_296; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_297 = io_pipe_phv_in_data_297; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_298 = io_pipe_phv_in_data_298; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_299 = io_pipe_phv_in_data_299; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_300 = io_pipe_phv_in_data_300; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_301 = io_pipe_phv_in_data_301; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_302 = io_pipe_phv_in_data_302; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_303 = io_pipe_phv_in_data_303; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_304 = io_pipe_phv_in_data_304; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_305 = io_pipe_phv_in_data_305; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_306 = io_pipe_phv_in_data_306; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_307 = io_pipe_phv_in_data_307; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_308 = io_pipe_phv_in_data_308; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_309 = io_pipe_phv_in_data_309; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_310 = io_pipe_phv_in_data_310; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_311 = io_pipe_phv_in_data_311; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_312 = io_pipe_phv_in_data_312; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_313 = io_pipe_phv_in_data_313; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_314 = io_pipe_phv_in_data_314; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_315 = io_pipe_phv_in_data_315; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_316 = io_pipe_phv_in_data_316; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_317 = io_pipe_phv_in_data_317; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_318 = io_pipe_phv_in_data_318; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_319 = io_pipe_phv_in_data_319; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_320 = io_pipe_phv_in_data_320; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_321 = io_pipe_phv_in_data_321; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_322 = io_pipe_phv_in_data_322; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_323 = io_pipe_phv_in_data_323; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_324 = io_pipe_phv_in_data_324; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_325 = io_pipe_phv_in_data_325; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_326 = io_pipe_phv_in_data_326; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_327 = io_pipe_phv_in_data_327; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_328 = io_pipe_phv_in_data_328; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_329 = io_pipe_phv_in_data_329; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_330 = io_pipe_phv_in_data_330; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_331 = io_pipe_phv_in_data_331; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_332 = io_pipe_phv_in_data_332; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_333 = io_pipe_phv_in_data_333; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_334 = io_pipe_phv_in_data_334; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_335 = io_pipe_phv_in_data_335; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_336 = io_pipe_phv_in_data_336; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_337 = io_pipe_phv_in_data_337; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_338 = io_pipe_phv_in_data_338; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_339 = io_pipe_phv_in_data_339; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_340 = io_pipe_phv_in_data_340; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_341 = io_pipe_phv_in_data_341; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_342 = io_pipe_phv_in_data_342; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_343 = io_pipe_phv_in_data_343; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_344 = io_pipe_phv_in_data_344; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_345 = io_pipe_phv_in_data_345; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_346 = io_pipe_phv_in_data_346; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_347 = io_pipe_phv_in_data_347; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_348 = io_pipe_phv_in_data_348; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_349 = io_pipe_phv_in_data_349; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_350 = io_pipe_phv_in_data_350; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_351 = io_pipe_phv_in_data_351; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_352 = io_pipe_phv_in_data_352; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_353 = io_pipe_phv_in_data_353; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_354 = io_pipe_phv_in_data_354; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_355 = io_pipe_phv_in_data_355; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_356 = io_pipe_phv_in_data_356; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_357 = io_pipe_phv_in_data_357; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_358 = io_pipe_phv_in_data_358; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_359 = io_pipe_phv_in_data_359; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_360 = io_pipe_phv_in_data_360; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_361 = io_pipe_phv_in_data_361; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_362 = io_pipe_phv_in_data_362; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_363 = io_pipe_phv_in_data_363; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_364 = io_pipe_phv_in_data_364; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_365 = io_pipe_phv_in_data_365; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_366 = io_pipe_phv_in_data_366; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_367 = io_pipe_phv_in_data_367; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_368 = io_pipe_phv_in_data_368; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_369 = io_pipe_phv_in_data_369; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_370 = io_pipe_phv_in_data_370; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_371 = io_pipe_phv_in_data_371; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_372 = io_pipe_phv_in_data_372; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_373 = io_pipe_phv_in_data_373; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_374 = io_pipe_phv_in_data_374; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_375 = io_pipe_phv_in_data_375; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_376 = io_pipe_phv_in_data_376; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_377 = io_pipe_phv_in_data_377; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_378 = io_pipe_phv_in_data_378; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_379 = io_pipe_phv_in_data_379; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_380 = io_pipe_phv_in_data_380; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_381 = io_pipe_phv_in_data_381; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_382 = io_pipe_phv_in_data_382; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_383 = io_pipe_phv_in_data_383; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_384 = io_pipe_phv_in_data_384; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_385 = io_pipe_phv_in_data_385; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_386 = io_pipe_phv_in_data_386; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_387 = io_pipe_phv_in_data_387; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_388 = io_pipe_phv_in_data_388; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_389 = io_pipe_phv_in_data_389; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_390 = io_pipe_phv_in_data_390; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_391 = io_pipe_phv_in_data_391; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_392 = io_pipe_phv_in_data_392; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_393 = io_pipe_phv_in_data_393; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_394 = io_pipe_phv_in_data_394; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_395 = io_pipe_phv_in_data_395; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_396 = io_pipe_phv_in_data_396; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_397 = io_pipe_phv_in_data_397; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_398 = io_pipe_phv_in_data_398; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_399 = io_pipe_phv_in_data_399; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_400 = io_pipe_phv_in_data_400; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_401 = io_pipe_phv_in_data_401; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_402 = io_pipe_phv_in_data_402; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_403 = io_pipe_phv_in_data_403; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_404 = io_pipe_phv_in_data_404; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_405 = io_pipe_phv_in_data_405; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_406 = io_pipe_phv_in_data_406; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_407 = io_pipe_phv_in_data_407; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_408 = io_pipe_phv_in_data_408; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_409 = io_pipe_phv_in_data_409; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_410 = io_pipe_phv_in_data_410; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_411 = io_pipe_phv_in_data_411; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_412 = io_pipe_phv_in_data_412; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_413 = io_pipe_phv_in_data_413; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_414 = io_pipe_phv_in_data_414; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_415 = io_pipe_phv_in_data_415; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_416 = io_pipe_phv_in_data_416; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_417 = io_pipe_phv_in_data_417; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_418 = io_pipe_phv_in_data_418; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_419 = io_pipe_phv_in_data_419; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_420 = io_pipe_phv_in_data_420; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_421 = io_pipe_phv_in_data_421; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_422 = io_pipe_phv_in_data_422; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_423 = io_pipe_phv_in_data_423; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_424 = io_pipe_phv_in_data_424; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_425 = io_pipe_phv_in_data_425; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_426 = io_pipe_phv_in_data_426; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_427 = io_pipe_phv_in_data_427; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_428 = io_pipe_phv_in_data_428; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_429 = io_pipe_phv_in_data_429; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_430 = io_pipe_phv_in_data_430; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_431 = io_pipe_phv_in_data_431; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_432 = io_pipe_phv_in_data_432; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_433 = io_pipe_phv_in_data_433; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_434 = io_pipe_phv_in_data_434; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_435 = io_pipe_phv_in_data_435; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_436 = io_pipe_phv_in_data_436; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_437 = io_pipe_phv_in_data_437; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_438 = io_pipe_phv_in_data_438; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_439 = io_pipe_phv_in_data_439; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_440 = io_pipe_phv_in_data_440; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_441 = io_pipe_phv_in_data_441; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_442 = io_pipe_phv_in_data_442; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_443 = io_pipe_phv_in_data_443; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_444 = io_pipe_phv_in_data_444; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_445 = io_pipe_phv_in_data_445; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_446 = io_pipe_phv_in_data_446; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_447 = io_pipe_phv_in_data_447; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_448 = io_pipe_phv_in_data_448; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_449 = io_pipe_phv_in_data_449; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_450 = io_pipe_phv_in_data_450; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_451 = io_pipe_phv_in_data_451; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_452 = io_pipe_phv_in_data_452; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_453 = io_pipe_phv_in_data_453; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_454 = io_pipe_phv_in_data_454; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_455 = io_pipe_phv_in_data_455; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_456 = io_pipe_phv_in_data_456; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_457 = io_pipe_phv_in_data_457; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_458 = io_pipe_phv_in_data_458; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_459 = io_pipe_phv_in_data_459; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_460 = io_pipe_phv_in_data_460; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_461 = io_pipe_phv_in_data_461; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_462 = io_pipe_phv_in_data_462; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_463 = io_pipe_phv_in_data_463; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_464 = io_pipe_phv_in_data_464; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_465 = io_pipe_phv_in_data_465; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_466 = io_pipe_phv_in_data_466; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_467 = io_pipe_phv_in_data_467; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_468 = io_pipe_phv_in_data_468; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_469 = io_pipe_phv_in_data_469; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_470 = io_pipe_phv_in_data_470; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_471 = io_pipe_phv_in_data_471; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_472 = io_pipe_phv_in_data_472; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_473 = io_pipe_phv_in_data_473; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_474 = io_pipe_phv_in_data_474; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_475 = io_pipe_phv_in_data_475; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_476 = io_pipe_phv_in_data_476; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_477 = io_pipe_phv_in_data_477; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_478 = io_pipe_phv_in_data_478; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_479 = io_pipe_phv_in_data_479; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_480 = io_pipe_phv_in_data_480; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_481 = io_pipe_phv_in_data_481; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_482 = io_pipe_phv_in_data_482; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_483 = io_pipe_phv_in_data_483; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_484 = io_pipe_phv_in_data_484; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_485 = io_pipe_phv_in_data_485; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_486 = io_pipe_phv_in_data_486; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_487 = io_pipe_phv_in_data_487; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_488 = io_pipe_phv_in_data_488; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_489 = io_pipe_phv_in_data_489; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_490 = io_pipe_phv_in_data_490; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_491 = io_pipe_phv_in_data_491; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_492 = io_pipe_phv_in_data_492; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_493 = io_pipe_phv_in_data_493; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_494 = io_pipe_phv_in_data_494; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_495 = io_pipe_phv_in_data_495; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_496 = io_pipe_phv_in_data_496; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_497 = io_pipe_phv_in_data_497; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_498 = io_pipe_phv_in_data_498; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_499 = io_pipe_phv_in_data_499; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_500 = io_pipe_phv_in_data_500; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_501 = io_pipe_phv_in_data_501; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_502 = io_pipe_phv_in_data_502; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_503 = io_pipe_phv_in_data_503; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_504 = io_pipe_phv_in_data_504; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_505 = io_pipe_phv_in_data_505; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_506 = io_pipe_phv_in_data_506; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_507 = io_pipe_phv_in_data_507; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_508 = io_pipe_phv_in_data_508; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_509 = io_pipe_phv_in_data_509; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_510 = io_pipe_phv_in_data_510; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_data_511 = io_pipe_phv_in_data_511; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[parser.scala 30:35]
  assign mau_0_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[parser.scala 30:35]
  assign mau_0_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j : io_mod_module_mod_state_id_mod
    ; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_0_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_0_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_0_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_0_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_0_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  assign mau_1_clock = clock;
  assign mau_1_io_pipe_phv_in_data_0 = mau_0_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_1 = mau_0_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_2 = mau_0_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_3 = mau_0_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_4 = mau_0_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_5 = mau_0_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_6 = mau_0_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_7 = mau_0_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_8 = mau_0_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_9 = mau_0_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_10 = mau_0_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_11 = mau_0_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_12 = mau_0_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_13 = mau_0_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_14 = mau_0_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_15 = mau_0_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_16 = mau_0_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_17 = mau_0_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_18 = mau_0_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_19 = mau_0_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_20 = mau_0_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_21 = mau_0_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_22 = mau_0_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_23 = mau_0_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_24 = mau_0_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_25 = mau_0_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_26 = mau_0_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_27 = mau_0_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_28 = mau_0_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_29 = mau_0_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_30 = mau_0_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_31 = mau_0_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_32 = mau_0_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_33 = mau_0_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_34 = mau_0_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_35 = mau_0_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_36 = mau_0_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_37 = mau_0_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_38 = mau_0_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_39 = mau_0_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_40 = mau_0_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_41 = mau_0_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_42 = mau_0_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_43 = mau_0_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_44 = mau_0_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_45 = mau_0_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_46 = mau_0_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_47 = mau_0_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_48 = mau_0_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_49 = mau_0_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_50 = mau_0_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_51 = mau_0_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_52 = mau_0_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_53 = mau_0_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_54 = mau_0_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_55 = mau_0_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_56 = mau_0_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_57 = mau_0_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_58 = mau_0_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_59 = mau_0_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_60 = mau_0_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_61 = mau_0_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_62 = mau_0_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_63 = mau_0_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_64 = mau_0_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_65 = mau_0_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_66 = mau_0_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_67 = mau_0_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_68 = mau_0_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_69 = mau_0_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_70 = mau_0_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_71 = mau_0_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_72 = mau_0_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_73 = mau_0_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_74 = mau_0_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_75 = mau_0_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_76 = mau_0_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_77 = mau_0_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_78 = mau_0_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_79 = mau_0_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_80 = mau_0_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_81 = mau_0_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_82 = mau_0_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_83 = mau_0_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_84 = mau_0_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_85 = mau_0_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_86 = mau_0_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_87 = mau_0_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_88 = mau_0_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_89 = mau_0_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_90 = mau_0_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_91 = mau_0_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_92 = mau_0_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_93 = mau_0_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_94 = mau_0_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_95 = mau_0_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_96 = mau_0_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_97 = mau_0_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_98 = mau_0_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_99 = mau_0_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_100 = mau_0_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_101 = mau_0_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_102 = mau_0_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_103 = mau_0_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_104 = mau_0_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_105 = mau_0_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_106 = mau_0_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_107 = mau_0_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_108 = mau_0_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_109 = mau_0_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_110 = mau_0_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_111 = mau_0_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_112 = mau_0_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_113 = mau_0_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_114 = mau_0_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_115 = mau_0_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_116 = mau_0_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_117 = mau_0_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_118 = mau_0_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_119 = mau_0_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_120 = mau_0_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_121 = mau_0_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_122 = mau_0_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_123 = mau_0_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_124 = mau_0_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_125 = mau_0_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_126 = mau_0_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_127 = mau_0_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_128 = mau_0_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_129 = mau_0_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_130 = mau_0_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_131 = mau_0_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_132 = mau_0_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_133 = mau_0_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_134 = mau_0_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_135 = mau_0_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_136 = mau_0_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_137 = mau_0_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_138 = mau_0_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_139 = mau_0_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_140 = mau_0_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_141 = mau_0_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_142 = mau_0_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_143 = mau_0_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_144 = mau_0_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_145 = mau_0_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_146 = mau_0_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_147 = mau_0_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_148 = mau_0_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_149 = mau_0_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_150 = mau_0_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_151 = mau_0_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_152 = mau_0_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_153 = mau_0_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_154 = mau_0_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_155 = mau_0_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_156 = mau_0_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_157 = mau_0_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_158 = mau_0_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_159 = mau_0_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_160 = mau_0_io_pipe_phv_out_data_160; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_161 = mau_0_io_pipe_phv_out_data_161; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_162 = mau_0_io_pipe_phv_out_data_162; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_163 = mau_0_io_pipe_phv_out_data_163; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_164 = mau_0_io_pipe_phv_out_data_164; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_165 = mau_0_io_pipe_phv_out_data_165; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_166 = mau_0_io_pipe_phv_out_data_166; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_167 = mau_0_io_pipe_phv_out_data_167; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_168 = mau_0_io_pipe_phv_out_data_168; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_169 = mau_0_io_pipe_phv_out_data_169; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_170 = mau_0_io_pipe_phv_out_data_170; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_171 = mau_0_io_pipe_phv_out_data_171; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_172 = mau_0_io_pipe_phv_out_data_172; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_173 = mau_0_io_pipe_phv_out_data_173; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_174 = mau_0_io_pipe_phv_out_data_174; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_175 = mau_0_io_pipe_phv_out_data_175; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_176 = mau_0_io_pipe_phv_out_data_176; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_177 = mau_0_io_pipe_phv_out_data_177; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_178 = mau_0_io_pipe_phv_out_data_178; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_179 = mau_0_io_pipe_phv_out_data_179; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_180 = mau_0_io_pipe_phv_out_data_180; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_181 = mau_0_io_pipe_phv_out_data_181; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_182 = mau_0_io_pipe_phv_out_data_182; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_183 = mau_0_io_pipe_phv_out_data_183; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_184 = mau_0_io_pipe_phv_out_data_184; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_185 = mau_0_io_pipe_phv_out_data_185; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_186 = mau_0_io_pipe_phv_out_data_186; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_187 = mau_0_io_pipe_phv_out_data_187; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_188 = mau_0_io_pipe_phv_out_data_188; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_189 = mau_0_io_pipe_phv_out_data_189; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_190 = mau_0_io_pipe_phv_out_data_190; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_191 = mau_0_io_pipe_phv_out_data_191; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_192 = mau_0_io_pipe_phv_out_data_192; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_193 = mau_0_io_pipe_phv_out_data_193; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_194 = mau_0_io_pipe_phv_out_data_194; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_195 = mau_0_io_pipe_phv_out_data_195; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_196 = mau_0_io_pipe_phv_out_data_196; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_197 = mau_0_io_pipe_phv_out_data_197; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_198 = mau_0_io_pipe_phv_out_data_198; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_199 = mau_0_io_pipe_phv_out_data_199; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_200 = mau_0_io_pipe_phv_out_data_200; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_201 = mau_0_io_pipe_phv_out_data_201; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_202 = mau_0_io_pipe_phv_out_data_202; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_203 = mau_0_io_pipe_phv_out_data_203; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_204 = mau_0_io_pipe_phv_out_data_204; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_205 = mau_0_io_pipe_phv_out_data_205; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_206 = mau_0_io_pipe_phv_out_data_206; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_207 = mau_0_io_pipe_phv_out_data_207; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_208 = mau_0_io_pipe_phv_out_data_208; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_209 = mau_0_io_pipe_phv_out_data_209; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_210 = mau_0_io_pipe_phv_out_data_210; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_211 = mau_0_io_pipe_phv_out_data_211; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_212 = mau_0_io_pipe_phv_out_data_212; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_213 = mau_0_io_pipe_phv_out_data_213; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_214 = mau_0_io_pipe_phv_out_data_214; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_215 = mau_0_io_pipe_phv_out_data_215; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_216 = mau_0_io_pipe_phv_out_data_216; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_217 = mau_0_io_pipe_phv_out_data_217; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_218 = mau_0_io_pipe_phv_out_data_218; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_219 = mau_0_io_pipe_phv_out_data_219; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_220 = mau_0_io_pipe_phv_out_data_220; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_221 = mau_0_io_pipe_phv_out_data_221; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_222 = mau_0_io_pipe_phv_out_data_222; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_223 = mau_0_io_pipe_phv_out_data_223; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_224 = mau_0_io_pipe_phv_out_data_224; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_225 = mau_0_io_pipe_phv_out_data_225; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_226 = mau_0_io_pipe_phv_out_data_226; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_227 = mau_0_io_pipe_phv_out_data_227; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_228 = mau_0_io_pipe_phv_out_data_228; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_229 = mau_0_io_pipe_phv_out_data_229; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_230 = mau_0_io_pipe_phv_out_data_230; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_231 = mau_0_io_pipe_phv_out_data_231; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_232 = mau_0_io_pipe_phv_out_data_232; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_233 = mau_0_io_pipe_phv_out_data_233; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_234 = mau_0_io_pipe_phv_out_data_234; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_235 = mau_0_io_pipe_phv_out_data_235; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_236 = mau_0_io_pipe_phv_out_data_236; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_237 = mau_0_io_pipe_phv_out_data_237; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_238 = mau_0_io_pipe_phv_out_data_238; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_239 = mau_0_io_pipe_phv_out_data_239; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_240 = mau_0_io_pipe_phv_out_data_240; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_241 = mau_0_io_pipe_phv_out_data_241; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_242 = mau_0_io_pipe_phv_out_data_242; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_243 = mau_0_io_pipe_phv_out_data_243; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_244 = mau_0_io_pipe_phv_out_data_244; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_245 = mau_0_io_pipe_phv_out_data_245; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_246 = mau_0_io_pipe_phv_out_data_246; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_247 = mau_0_io_pipe_phv_out_data_247; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_248 = mau_0_io_pipe_phv_out_data_248; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_249 = mau_0_io_pipe_phv_out_data_249; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_250 = mau_0_io_pipe_phv_out_data_250; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_251 = mau_0_io_pipe_phv_out_data_251; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_252 = mau_0_io_pipe_phv_out_data_252; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_253 = mau_0_io_pipe_phv_out_data_253; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_254 = mau_0_io_pipe_phv_out_data_254; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_255 = mau_0_io_pipe_phv_out_data_255; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_256 = mau_0_io_pipe_phv_out_data_256; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_257 = mau_0_io_pipe_phv_out_data_257; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_258 = mau_0_io_pipe_phv_out_data_258; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_259 = mau_0_io_pipe_phv_out_data_259; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_260 = mau_0_io_pipe_phv_out_data_260; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_261 = mau_0_io_pipe_phv_out_data_261; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_262 = mau_0_io_pipe_phv_out_data_262; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_263 = mau_0_io_pipe_phv_out_data_263; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_264 = mau_0_io_pipe_phv_out_data_264; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_265 = mau_0_io_pipe_phv_out_data_265; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_266 = mau_0_io_pipe_phv_out_data_266; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_267 = mau_0_io_pipe_phv_out_data_267; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_268 = mau_0_io_pipe_phv_out_data_268; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_269 = mau_0_io_pipe_phv_out_data_269; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_270 = mau_0_io_pipe_phv_out_data_270; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_271 = mau_0_io_pipe_phv_out_data_271; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_272 = mau_0_io_pipe_phv_out_data_272; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_273 = mau_0_io_pipe_phv_out_data_273; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_274 = mau_0_io_pipe_phv_out_data_274; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_275 = mau_0_io_pipe_phv_out_data_275; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_276 = mau_0_io_pipe_phv_out_data_276; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_277 = mau_0_io_pipe_phv_out_data_277; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_278 = mau_0_io_pipe_phv_out_data_278; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_279 = mau_0_io_pipe_phv_out_data_279; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_280 = mau_0_io_pipe_phv_out_data_280; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_281 = mau_0_io_pipe_phv_out_data_281; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_282 = mau_0_io_pipe_phv_out_data_282; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_283 = mau_0_io_pipe_phv_out_data_283; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_284 = mau_0_io_pipe_phv_out_data_284; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_285 = mau_0_io_pipe_phv_out_data_285; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_286 = mau_0_io_pipe_phv_out_data_286; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_287 = mau_0_io_pipe_phv_out_data_287; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_288 = mau_0_io_pipe_phv_out_data_288; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_289 = mau_0_io_pipe_phv_out_data_289; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_290 = mau_0_io_pipe_phv_out_data_290; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_291 = mau_0_io_pipe_phv_out_data_291; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_292 = mau_0_io_pipe_phv_out_data_292; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_293 = mau_0_io_pipe_phv_out_data_293; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_294 = mau_0_io_pipe_phv_out_data_294; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_295 = mau_0_io_pipe_phv_out_data_295; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_296 = mau_0_io_pipe_phv_out_data_296; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_297 = mau_0_io_pipe_phv_out_data_297; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_298 = mau_0_io_pipe_phv_out_data_298; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_299 = mau_0_io_pipe_phv_out_data_299; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_300 = mau_0_io_pipe_phv_out_data_300; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_301 = mau_0_io_pipe_phv_out_data_301; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_302 = mau_0_io_pipe_phv_out_data_302; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_303 = mau_0_io_pipe_phv_out_data_303; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_304 = mau_0_io_pipe_phv_out_data_304; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_305 = mau_0_io_pipe_phv_out_data_305; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_306 = mau_0_io_pipe_phv_out_data_306; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_307 = mau_0_io_pipe_phv_out_data_307; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_308 = mau_0_io_pipe_phv_out_data_308; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_309 = mau_0_io_pipe_phv_out_data_309; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_310 = mau_0_io_pipe_phv_out_data_310; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_311 = mau_0_io_pipe_phv_out_data_311; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_312 = mau_0_io_pipe_phv_out_data_312; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_313 = mau_0_io_pipe_phv_out_data_313; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_314 = mau_0_io_pipe_phv_out_data_314; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_315 = mau_0_io_pipe_phv_out_data_315; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_316 = mau_0_io_pipe_phv_out_data_316; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_317 = mau_0_io_pipe_phv_out_data_317; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_318 = mau_0_io_pipe_phv_out_data_318; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_319 = mau_0_io_pipe_phv_out_data_319; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_320 = mau_0_io_pipe_phv_out_data_320; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_321 = mau_0_io_pipe_phv_out_data_321; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_322 = mau_0_io_pipe_phv_out_data_322; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_323 = mau_0_io_pipe_phv_out_data_323; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_324 = mau_0_io_pipe_phv_out_data_324; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_325 = mau_0_io_pipe_phv_out_data_325; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_326 = mau_0_io_pipe_phv_out_data_326; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_327 = mau_0_io_pipe_phv_out_data_327; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_328 = mau_0_io_pipe_phv_out_data_328; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_329 = mau_0_io_pipe_phv_out_data_329; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_330 = mau_0_io_pipe_phv_out_data_330; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_331 = mau_0_io_pipe_phv_out_data_331; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_332 = mau_0_io_pipe_phv_out_data_332; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_333 = mau_0_io_pipe_phv_out_data_333; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_334 = mau_0_io_pipe_phv_out_data_334; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_335 = mau_0_io_pipe_phv_out_data_335; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_336 = mau_0_io_pipe_phv_out_data_336; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_337 = mau_0_io_pipe_phv_out_data_337; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_338 = mau_0_io_pipe_phv_out_data_338; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_339 = mau_0_io_pipe_phv_out_data_339; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_340 = mau_0_io_pipe_phv_out_data_340; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_341 = mau_0_io_pipe_phv_out_data_341; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_342 = mau_0_io_pipe_phv_out_data_342; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_343 = mau_0_io_pipe_phv_out_data_343; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_344 = mau_0_io_pipe_phv_out_data_344; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_345 = mau_0_io_pipe_phv_out_data_345; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_346 = mau_0_io_pipe_phv_out_data_346; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_347 = mau_0_io_pipe_phv_out_data_347; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_348 = mau_0_io_pipe_phv_out_data_348; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_349 = mau_0_io_pipe_phv_out_data_349; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_350 = mau_0_io_pipe_phv_out_data_350; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_351 = mau_0_io_pipe_phv_out_data_351; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_352 = mau_0_io_pipe_phv_out_data_352; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_353 = mau_0_io_pipe_phv_out_data_353; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_354 = mau_0_io_pipe_phv_out_data_354; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_355 = mau_0_io_pipe_phv_out_data_355; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_356 = mau_0_io_pipe_phv_out_data_356; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_357 = mau_0_io_pipe_phv_out_data_357; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_358 = mau_0_io_pipe_phv_out_data_358; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_359 = mau_0_io_pipe_phv_out_data_359; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_360 = mau_0_io_pipe_phv_out_data_360; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_361 = mau_0_io_pipe_phv_out_data_361; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_362 = mau_0_io_pipe_phv_out_data_362; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_363 = mau_0_io_pipe_phv_out_data_363; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_364 = mau_0_io_pipe_phv_out_data_364; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_365 = mau_0_io_pipe_phv_out_data_365; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_366 = mau_0_io_pipe_phv_out_data_366; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_367 = mau_0_io_pipe_phv_out_data_367; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_368 = mau_0_io_pipe_phv_out_data_368; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_369 = mau_0_io_pipe_phv_out_data_369; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_370 = mau_0_io_pipe_phv_out_data_370; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_371 = mau_0_io_pipe_phv_out_data_371; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_372 = mau_0_io_pipe_phv_out_data_372; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_373 = mau_0_io_pipe_phv_out_data_373; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_374 = mau_0_io_pipe_phv_out_data_374; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_375 = mau_0_io_pipe_phv_out_data_375; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_376 = mau_0_io_pipe_phv_out_data_376; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_377 = mau_0_io_pipe_phv_out_data_377; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_378 = mau_0_io_pipe_phv_out_data_378; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_379 = mau_0_io_pipe_phv_out_data_379; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_380 = mau_0_io_pipe_phv_out_data_380; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_381 = mau_0_io_pipe_phv_out_data_381; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_382 = mau_0_io_pipe_phv_out_data_382; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_383 = mau_0_io_pipe_phv_out_data_383; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_384 = mau_0_io_pipe_phv_out_data_384; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_385 = mau_0_io_pipe_phv_out_data_385; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_386 = mau_0_io_pipe_phv_out_data_386; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_387 = mau_0_io_pipe_phv_out_data_387; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_388 = mau_0_io_pipe_phv_out_data_388; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_389 = mau_0_io_pipe_phv_out_data_389; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_390 = mau_0_io_pipe_phv_out_data_390; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_391 = mau_0_io_pipe_phv_out_data_391; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_392 = mau_0_io_pipe_phv_out_data_392; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_393 = mau_0_io_pipe_phv_out_data_393; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_394 = mau_0_io_pipe_phv_out_data_394; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_395 = mau_0_io_pipe_phv_out_data_395; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_396 = mau_0_io_pipe_phv_out_data_396; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_397 = mau_0_io_pipe_phv_out_data_397; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_398 = mau_0_io_pipe_phv_out_data_398; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_399 = mau_0_io_pipe_phv_out_data_399; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_400 = mau_0_io_pipe_phv_out_data_400; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_401 = mau_0_io_pipe_phv_out_data_401; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_402 = mau_0_io_pipe_phv_out_data_402; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_403 = mau_0_io_pipe_phv_out_data_403; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_404 = mau_0_io_pipe_phv_out_data_404; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_405 = mau_0_io_pipe_phv_out_data_405; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_406 = mau_0_io_pipe_phv_out_data_406; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_407 = mau_0_io_pipe_phv_out_data_407; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_408 = mau_0_io_pipe_phv_out_data_408; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_409 = mau_0_io_pipe_phv_out_data_409; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_410 = mau_0_io_pipe_phv_out_data_410; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_411 = mau_0_io_pipe_phv_out_data_411; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_412 = mau_0_io_pipe_phv_out_data_412; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_413 = mau_0_io_pipe_phv_out_data_413; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_414 = mau_0_io_pipe_phv_out_data_414; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_415 = mau_0_io_pipe_phv_out_data_415; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_416 = mau_0_io_pipe_phv_out_data_416; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_417 = mau_0_io_pipe_phv_out_data_417; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_418 = mau_0_io_pipe_phv_out_data_418; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_419 = mau_0_io_pipe_phv_out_data_419; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_420 = mau_0_io_pipe_phv_out_data_420; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_421 = mau_0_io_pipe_phv_out_data_421; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_422 = mau_0_io_pipe_phv_out_data_422; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_423 = mau_0_io_pipe_phv_out_data_423; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_424 = mau_0_io_pipe_phv_out_data_424; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_425 = mau_0_io_pipe_phv_out_data_425; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_426 = mau_0_io_pipe_phv_out_data_426; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_427 = mau_0_io_pipe_phv_out_data_427; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_428 = mau_0_io_pipe_phv_out_data_428; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_429 = mau_0_io_pipe_phv_out_data_429; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_430 = mau_0_io_pipe_phv_out_data_430; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_431 = mau_0_io_pipe_phv_out_data_431; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_432 = mau_0_io_pipe_phv_out_data_432; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_433 = mau_0_io_pipe_phv_out_data_433; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_434 = mau_0_io_pipe_phv_out_data_434; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_435 = mau_0_io_pipe_phv_out_data_435; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_436 = mau_0_io_pipe_phv_out_data_436; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_437 = mau_0_io_pipe_phv_out_data_437; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_438 = mau_0_io_pipe_phv_out_data_438; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_439 = mau_0_io_pipe_phv_out_data_439; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_440 = mau_0_io_pipe_phv_out_data_440; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_441 = mau_0_io_pipe_phv_out_data_441; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_442 = mau_0_io_pipe_phv_out_data_442; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_443 = mau_0_io_pipe_phv_out_data_443; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_444 = mau_0_io_pipe_phv_out_data_444; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_445 = mau_0_io_pipe_phv_out_data_445; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_446 = mau_0_io_pipe_phv_out_data_446; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_447 = mau_0_io_pipe_phv_out_data_447; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_448 = mau_0_io_pipe_phv_out_data_448; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_449 = mau_0_io_pipe_phv_out_data_449; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_450 = mau_0_io_pipe_phv_out_data_450; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_451 = mau_0_io_pipe_phv_out_data_451; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_452 = mau_0_io_pipe_phv_out_data_452; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_453 = mau_0_io_pipe_phv_out_data_453; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_454 = mau_0_io_pipe_phv_out_data_454; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_455 = mau_0_io_pipe_phv_out_data_455; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_456 = mau_0_io_pipe_phv_out_data_456; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_457 = mau_0_io_pipe_phv_out_data_457; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_458 = mau_0_io_pipe_phv_out_data_458; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_459 = mau_0_io_pipe_phv_out_data_459; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_460 = mau_0_io_pipe_phv_out_data_460; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_461 = mau_0_io_pipe_phv_out_data_461; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_462 = mau_0_io_pipe_phv_out_data_462; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_463 = mau_0_io_pipe_phv_out_data_463; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_464 = mau_0_io_pipe_phv_out_data_464; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_465 = mau_0_io_pipe_phv_out_data_465; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_466 = mau_0_io_pipe_phv_out_data_466; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_467 = mau_0_io_pipe_phv_out_data_467; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_468 = mau_0_io_pipe_phv_out_data_468; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_469 = mau_0_io_pipe_phv_out_data_469; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_470 = mau_0_io_pipe_phv_out_data_470; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_471 = mau_0_io_pipe_phv_out_data_471; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_472 = mau_0_io_pipe_phv_out_data_472; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_473 = mau_0_io_pipe_phv_out_data_473; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_474 = mau_0_io_pipe_phv_out_data_474; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_475 = mau_0_io_pipe_phv_out_data_475; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_476 = mau_0_io_pipe_phv_out_data_476; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_477 = mau_0_io_pipe_phv_out_data_477; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_478 = mau_0_io_pipe_phv_out_data_478; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_479 = mau_0_io_pipe_phv_out_data_479; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_480 = mau_0_io_pipe_phv_out_data_480; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_481 = mau_0_io_pipe_phv_out_data_481; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_482 = mau_0_io_pipe_phv_out_data_482; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_483 = mau_0_io_pipe_phv_out_data_483; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_484 = mau_0_io_pipe_phv_out_data_484; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_485 = mau_0_io_pipe_phv_out_data_485; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_486 = mau_0_io_pipe_phv_out_data_486; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_487 = mau_0_io_pipe_phv_out_data_487; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_488 = mau_0_io_pipe_phv_out_data_488; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_489 = mau_0_io_pipe_phv_out_data_489; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_490 = mau_0_io_pipe_phv_out_data_490; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_491 = mau_0_io_pipe_phv_out_data_491; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_492 = mau_0_io_pipe_phv_out_data_492; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_493 = mau_0_io_pipe_phv_out_data_493; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_494 = mau_0_io_pipe_phv_out_data_494; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_495 = mau_0_io_pipe_phv_out_data_495; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_496 = mau_0_io_pipe_phv_out_data_496; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_497 = mau_0_io_pipe_phv_out_data_497; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_498 = mau_0_io_pipe_phv_out_data_498; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_499 = mau_0_io_pipe_phv_out_data_499; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_500 = mau_0_io_pipe_phv_out_data_500; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_501 = mau_0_io_pipe_phv_out_data_501; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_502 = mau_0_io_pipe_phv_out_data_502; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_503 = mau_0_io_pipe_phv_out_data_503; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_504 = mau_0_io_pipe_phv_out_data_504; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_505 = mau_0_io_pipe_phv_out_data_505; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_506 = mau_0_io_pipe_phv_out_data_506; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_507 = mau_0_io_pipe_phv_out_data_507; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_508 = mau_0_io_pipe_phv_out_data_508; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_509 = mau_0_io_pipe_phv_out_data_509; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_510 = mau_0_io_pipe_phv_out_data_510; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_data_511 = mau_0_io_pipe_phv_out_data_511; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_0 = mau_0_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_1 = mau_0_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_2 = mau_0_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_3 = mau_0_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_4 = mau_0_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_5 = mau_0_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_6 = mau_0_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_7 = mau_0_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_8 = mau_0_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_9 = mau_0_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_10 = mau_0_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_11 = mau_0_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_12 = mau_0_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_13 = mau_0_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_14 = mau_0_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_header_15 = mau_0_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_current_state = mau_0_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_current_offset = mau_0_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_parse_transition_field = mau_0_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_next_processor_id = mau_0_io_pipe_phv_out_next_processor_id; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_next_config_id = mau_0_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_1_io_pipe_phv_in_is_valid_processor = mau_0_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_1_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_1 :
    io_mod_module_mod_state_id_mod; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_1_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_1_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_1_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_1 : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_1_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_1_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  assign mau_2_clock = clock;
  assign mau_2_io_pipe_phv_in_data_0 = mau_1_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_1 = mau_1_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_2 = mau_1_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_3 = mau_1_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_4 = mau_1_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_5 = mau_1_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_6 = mau_1_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_7 = mau_1_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_8 = mau_1_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_9 = mau_1_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_10 = mau_1_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_11 = mau_1_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_12 = mau_1_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_13 = mau_1_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_14 = mau_1_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_15 = mau_1_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_16 = mau_1_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_17 = mau_1_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_18 = mau_1_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_19 = mau_1_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_20 = mau_1_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_21 = mau_1_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_22 = mau_1_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_23 = mau_1_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_24 = mau_1_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_25 = mau_1_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_26 = mau_1_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_27 = mau_1_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_28 = mau_1_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_29 = mau_1_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_30 = mau_1_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_31 = mau_1_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_32 = mau_1_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_33 = mau_1_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_34 = mau_1_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_35 = mau_1_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_36 = mau_1_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_37 = mau_1_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_38 = mau_1_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_39 = mau_1_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_40 = mau_1_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_41 = mau_1_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_42 = mau_1_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_43 = mau_1_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_44 = mau_1_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_45 = mau_1_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_46 = mau_1_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_47 = mau_1_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_48 = mau_1_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_49 = mau_1_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_50 = mau_1_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_51 = mau_1_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_52 = mau_1_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_53 = mau_1_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_54 = mau_1_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_55 = mau_1_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_56 = mau_1_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_57 = mau_1_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_58 = mau_1_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_59 = mau_1_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_60 = mau_1_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_61 = mau_1_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_62 = mau_1_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_63 = mau_1_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_64 = mau_1_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_65 = mau_1_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_66 = mau_1_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_67 = mau_1_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_68 = mau_1_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_69 = mau_1_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_70 = mau_1_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_71 = mau_1_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_72 = mau_1_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_73 = mau_1_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_74 = mau_1_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_75 = mau_1_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_76 = mau_1_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_77 = mau_1_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_78 = mau_1_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_79 = mau_1_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_80 = mau_1_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_81 = mau_1_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_82 = mau_1_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_83 = mau_1_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_84 = mau_1_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_85 = mau_1_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_86 = mau_1_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_87 = mau_1_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_88 = mau_1_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_89 = mau_1_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_90 = mau_1_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_91 = mau_1_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_92 = mau_1_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_93 = mau_1_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_94 = mau_1_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_95 = mau_1_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_96 = mau_1_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_97 = mau_1_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_98 = mau_1_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_99 = mau_1_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_100 = mau_1_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_101 = mau_1_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_102 = mau_1_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_103 = mau_1_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_104 = mau_1_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_105 = mau_1_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_106 = mau_1_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_107 = mau_1_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_108 = mau_1_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_109 = mau_1_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_110 = mau_1_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_111 = mau_1_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_112 = mau_1_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_113 = mau_1_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_114 = mau_1_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_115 = mau_1_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_116 = mau_1_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_117 = mau_1_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_118 = mau_1_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_119 = mau_1_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_120 = mau_1_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_121 = mau_1_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_122 = mau_1_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_123 = mau_1_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_124 = mau_1_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_125 = mau_1_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_126 = mau_1_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_127 = mau_1_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_128 = mau_1_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_129 = mau_1_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_130 = mau_1_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_131 = mau_1_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_132 = mau_1_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_133 = mau_1_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_134 = mau_1_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_135 = mau_1_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_136 = mau_1_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_137 = mau_1_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_138 = mau_1_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_139 = mau_1_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_140 = mau_1_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_141 = mau_1_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_142 = mau_1_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_143 = mau_1_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_144 = mau_1_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_145 = mau_1_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_146 = mau_1_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_147 = mau_1_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_148 = mau_1_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_149 = mau_1_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_150 = mau_1_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_151 = mau_1_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_152 = mau_1_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_153 = mau_1_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_154 = mau_1_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_155 = mau_1_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_156 = mau_1_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_157 = mau_1_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_158 = mau_1_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_159 = mau_1_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_160 = mau_1_io_pipe_phv_out_data_160; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_161 = mau_1_io_pipe_phv_out_data_161; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_162 = mau_1_io_pipe_phv_out_data_162; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_163 = mau_1_io_pipe_phv_out_data_163; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_164 = mau_1_io_pipe_phv_out_data_164; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_165 = mau_1_io_pipe_phv_out_data_165; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_166 = mau_1_io_pipe_phv_out_data_166; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_167 = mau_1_io_pipe_phv_out_data_167; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_168 = mau_1_io_pipe_phv_out_data_168; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_169 = mau_1_io_pipe_phv_out_data_169; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_170 = mau_1_io_pipe_phv_out_data_170; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_171 = mau_1_io_pipe_phv_out_data_171; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_172 = mau_1_io_pipe_phv_out_data_172; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_173 = mau_1_io_pipe_phv_out_data_173; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_174 = mau_1_io_pipe_phv_out_data_174; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_175 = mau_1_io_pipe_phv_out_data_175; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_176 = mau_1_io_pipe_phv_out_data_176; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_177 = mau_1_io_pipe_phv_out_data_177; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_178 = mau_1_io_pipe_phv_out_data_178; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_179 = mau_1_io_pipe_phv_out_data_179; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_180 = mau_1_io_pipe_phv_out_data_180; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_181 = mau_1_io_pipe_phv_out_data_181; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_182 = mau_1_io_pipe_phv_out_data_182; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_183 = mau_1_io_pipe_phv_out_data_183; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_184 = mau_1_io_pipe_phv_out_data_184; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_185 = mau_1_io_pipe_phv_out_data_185; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_186 = mau_1_io_pipe_phv_out_data_186; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_187 = mau_1_io_pipe_phv_out_data_187; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_188 = mau_1_io_pipe_phv_out_data_188; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_189 = mau_1_io_pipe_phv_out_data_189; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_190 = mau_1_io_pipe_phv_out_data_190; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_191 = mau_1_io_pipe_phv_out_data_191; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_192 = mau_1_io_pipe_phv_out_data_192; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_193 = mau_1_io_pipe_phv_out_data_193; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_194 = mau_1_io_pipe_phv_out_data_194; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_195 = mau_1_io_pipe_phv_out_data_195; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_196 = mau_1_io_pipe_phv_out_data_196; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_197 = mau_1_io_pipe_phv_out_data_197; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_198 = mau_1_io_pipe_phv_out_data_198; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_199 = mau_1_io_pipe_phv_out_data_199; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_200 = mau_1_io_pipe_phv_out_data_200; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_201 = mau_1_io_pipe_phv_out_data_201; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_202 = mau_1_io_pipe_phv_out_data_202; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_203 = mau_1_io_pipe_phv_out_data_203; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_204 = mau_1_io_pipe_phv_out_data_204; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_205 = mau_1_io_pipe_phv_out_data_205; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_206 = mau_1_io_pipe_phv_out_data_206; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_207 = mau_1_io_pipe_phv_out_data_207; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_208 = mau_1_io_pipe_phv_out_data_208; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_209 = mau_1_io_pipe_phv_out_data_209; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_210 = mau_1_io_pipe_phv_out_data_210; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_211 = mau_1_io_pipe_phv_out_data_211; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_212 = mau_1_io_pipe_phv_out_data_212; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_213 = mau_1_io_pipe_phv_out_data_213; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_214 = mau_1_io_pipe_phv_out_data_214; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_215 = mau_1_io_pipe_phv_out_data_215; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_216 = mau_1_io_pipe_phv_out_data_216; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_217 = mau_1_io_pipe_phv_out_data_217; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_218 = mau_1_io_pipe_phv_out_data_218; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_219 = mau_1_io_pipe_phv_out_data_219; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_220 = mau_1_io_pipe_phv_out_data_220; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_221 = mau_1_io_pipe_phv_out_data_221; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_222 = mau_1_io_pipe_phv_out_data_222; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_223 = mau_1_io_pipe_phv_out_data_223; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_224 = mau_1_io_pipe_phv_out_data_224; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_225 = mau_1_io_pipe_phv_out_data_225; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_226 = mau_1_io_pipe_phv_out_data_226; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_227 = mau_1_io_pipe_phv_out_data_227; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_228 = mau_1_io_pipe_phv_out_data_228; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_229 = mau_1_io_pipe_phv_out_data_229; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_230 = mau_1_io_pipe_phv_out_data_230; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_231 = mau_1_io_pipe_phv_out_data_231; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_232 = mau_1_io_pipe_phv_out_data_232; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_233 = mau_1_io_pipe_phv_out_data_233; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_234 = mau_1_io_pipe_phv_out_data_234; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_235 = mau_1_io_pipe_phv_out_data_235; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_236 = mau_1_io_pipe_phv_out_data_236; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_237 = mau_1_io_pipe_phv_out_data_237; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_238 = mau_1_io_pipe_phv_out_data_238; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_239 = mau_1_io_pipe_phv_out_data_239; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_240 = mau_1_io_pipe_phv_out_data_240; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_241 = mau_1_io_pipe_phv_out_data_241; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_242 = mau_1_io_pipe_phv_out_data_242; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_243 = mau_1_io_pipe_phv_out_data_243; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_244 = mau_1_io_pipe_phv_out_data_244; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_245 = mau_1_io_pipe_phv_out_data_245; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_246 = mau_1_io_pipe_phv_out_data_246; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_247 = mau_1_io_pipe_phv_out_data_247; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_248 = mau_1_io_pipe_phv_out_data_248; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_249 = mau_1_io_pipe_phv_out_data_249; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_250 = mau_1_io_pipe_phv_out_data_250; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_251 = mau_1_io_pipe_phv_out_data_251; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_252 = mau_1_io_pipe_phv_out_data_252; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_253 = mau_1_io_pipe_phv_out_data_253; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_254 = mau_1_io_pipe_phv_out_data_254; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_255 = mau_1_io_pipe_phv_out_data_255; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_256 = mau_1_io_pipe_phv_out_data_256; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_257 = mau_1_io_pipe_phv_out_data_257; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_258 = mau_1_io_pipe_phv_out_data_258; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_259 = mau_1_io_pipe_phv_out_data_259; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_260 = mau_1_io_pipe_phv_out_data_260; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_261 = mau_1_io_pipe_phv_out_data_261; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_262 = mau_1_io_pipe_phv_out_data_262; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_263 = mau_1_io_pipe_phv_out_data_263; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_264 = mau_1_io_pipe_phv_out_data_264; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_265 = mau_1_io_pipe_phv_out_data_265; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_266 = mau_1_io_pipe_phv_out_data_266; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_267 = mau_1_io_pipe_phv_out_data_267; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_268 = mau_1_io_pipe_phv_out_data_268; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_269 = mau_1_io_pipe_phv_out_data_269; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_270 = mau_1_io_pipe_phv_out_data_270; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_271 = mau_1_io_pipe_phv_out_data_271; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_272 = mau_1_io_pipe_phv_out_data_272; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_273 = mau_1_io_pipe_phv_out_data_273; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_274 = mau_1_io_pipe_phv_out_data_274; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_275 = mau_1_io_pipe_phv_out_data_275; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_276 = mau_1_io_pipe_phv_out_data_276; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_277 = mau_1_io_pipe_phv_out_data_277; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_278 = mau_1_io_pipe_phv_out_data_278; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_279 = mau_1_io_pipe_phv_out_data_279; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_280 = mau_1_io_pipe_phv_out_data_280; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_281 = mau_1_io_pipe_phv_out_data_281; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_282 = mau_1_io_pipe_phv_out_data_282; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_283 = mau_1_io_pipe_phv_out_data_283; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_284 = mau_1_io_pipe_phv_out_data_284; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_285 = mau_1_io_pipe_phv_out_data_285; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_286 = mau_1_io_pipe_phv_out_data_286; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_287 = mau_1_io_pipe_phv_out_data_287; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_288 = mau_1_io_pipe_phv_out_data_288; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_289 = mau_1_io_pipe_phv_out_data_289; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_290 = mau_1_io_pipe_phv_out_data_290; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_291 = mau_1_io_pipe_phv_out_data_291; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_292 = mau_1_io_pipe_phv_out_data_292; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_293 = mau_1_io_pipe_phv_out_data_293; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_294 = mau_1_io_pipe_phv_out_data_294; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_295 = mau_1_io_pipe_phv_out_data_295; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_296 = mau_1_io_pipe_phv_out_data_296; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_297 = mau_1_io_pipe_phv_out_data_297; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_298 = mau_1_io_pipe_phv_out_data_298; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_299 = mau_1_io_pipe_phv_out_data_299; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_300 = mau_1_io_pipe_phv_out_data_300; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_301 = mau_1_io_pipe_phv_out_data_301; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_302 = mau_1_io_pipe_phv_out_data_302; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_303 = mau_1_io_pipe_phv_out_data_303; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_304 = mau_1_io_pipe_phv_out_data_304; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_305 = mau_1_io_pipe_phv_out_data_305; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_306 = mau_1_io_pipe_phv_out_data_306; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_307 = mau_1_io_pipe_phv_out_data_307; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_308 = mau_1_io_pipe_phv_out_data_308; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_309 = mau_1_io_pipe_phv_out_data_309; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_310 = mau_1_io_pipe_phv_out_data_310; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_311 = mau_1_io_pipe_phv_out_data_311; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_312 = mau_1_io_pipe_phv_out_data_312; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_313 = mau_1_io_pipe_phv_out_data_313; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_314 = mau_1_io_pipe_phv_out_data_314; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_315 = mau_1_io_pipe_phv_out_data_315; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_316 = mau_1_io_pipe_phv_out_data_316; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_317 = mau_1_io_pipe_phv_out_data_317; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_318 = mau_1_io_pipe_phv_out_data_318; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_319 = mau_1_io_pipe_phv_out_data_319; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_320 = mau_1_io_pipe_phv_out_data_320; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_321 = mau_1_io_pipe_phv_out_data_321; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_322 = mau_1_io_pipe_phv_out_data_322; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_323 = mau_1_io_pipe_phv_out_data_323; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_324 = mau_1_io_pipe_phv_out_data_324; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_325 = mau_1_io_pipe_phv_out_data_325; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_326 = mau_1_io_pipe_phv_out_data_326; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_327 = mau_1_io_pipe_phv_out_data_327; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_328 = mau_1_io_pipe_phv_out_data_328; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_329 = mau_1_io_pipe_phv_out_data_329; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_330 = mau_1_io_pipe_phv_out_data_330; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_331 = mau_1_io_pipe_phv_out_data_331; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_332 = mau_1_io_pipe_phv_out_data_332; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_333 = mau_1_io_pipe_phv_out_data_333; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_334 = mau_1_io_pipe_phv_out_data_334; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_335 = mau_1_io_pipe_phv_out_data_335; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_336 = mau_1_io_pipe_phv_out_data_336; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_337 = mau_1_io_pipe_phv_out_data_337; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_338 = mau_1_io_pipe_phv_out_data_338; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_339 = mau_1_io_pipe_phv_out_data_339; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_340 = mau_1_io_pipe_phv_out_data_340; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_341 = mau_1_io_pipe_phv_out_data_341; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_342 = mau_1_io_pipe_phv_out_data_342; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_343 = mau_1_io_pipe_phv_out_data_343; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_344 = mau_1_io_pipe_phv_out_data_344; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_345 = mau_1_io_pipe_phv_out_data_345; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_346 = mau_1_io_pipe_phv_out_data_346; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_347 = mau_1_io_pipe_phv_out_data_347; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_348 = mau_1_io_pipe_phv_out_data_348; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_349 = mau_1_io_pipe_phv_out_data_349; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_350 = mau_1_io_pipe_phv_out_data_350; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_351 = mau_1_io_pipe_phv_out_data_351; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_352 = mau_1_io_pipe_phv_out_data_352; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_353 = mau_1_io_pipe_phv_out_data_353; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_354 = mau_1_io_pipe_phv_out_data_354; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_355 = mau_1_io_pipe_phv_out_data_355; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_356 = mau_1_io_pipe_phv_out_data_356; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_357 = mau_1_io_pipe_phv_out_data_357; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_358 = mau_1_io_pipe_phv_out_data_358; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_359 = mau_1_io_pipe_phv_out_data_359; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_360 = mau_1_io_pipe_phv_out_data_360; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_361 = mau_1_io_pipe_phv_out_data_361; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_362 = mau_1_io_pipe_phv_out_data_362; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_363 = mau_1_io_pipe_phv_out_data_363; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_364 = mau_1_io_pipe_phv_out_data_364; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_365 = mau_1_io_pipe_phv_out_data_365; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_366 = mau_1_io_pipe_phv_out_data_366; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_367 = mau_1_io_pipe_phv_out_data_367; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_368 = mau_1_io_pipe_phv_out_data_368; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_369 = mau_1_io_pipe_phv_out_data_369; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_370 = mau_1_io_pipe_phv_out_data_370; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_371 = mau_1_io_pipe_phv_out_data_371; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_372 = mau_1_io_pipe_phv_out_data_372; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_373 = mau_1_io_pipe_phv_out_data_373; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_374 = mau_1_io_pipe_phv_out_data_374; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_375 = mau_1_io_pipe_phv_out_data_375; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_376 = mau_1_io_pipe_phv_out_data_376; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_377 = mau_1_io_pipe_phv_out_data_377; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_378 = mau_1_io_pipe_phv_out_data_378; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_379 = mau_1_io_pipe_phv_out_data_379; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_380 = mau_1_io_pipe_phv_out_data_380; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_381 = mau_1_io_pipe_phv_out_data_381; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_382 = mau_1_io_pipe_phv_out_data_382; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_383 = mau_1_io_pipe_phv_out_data_383; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_384 = mau_1_io_pipe_phv_out_data_384; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_385 = mau_1_io_pipe_phv_out_data_385; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_386 = mau_1_io_pipe_phv_out_data_386; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_387 = mau_1_io_pipe_phv_out_data_387; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_388 = mau_1_io_pipe_phv_out_data_388; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_389 = mau_1_io_pipe_phv_out_data_389; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_390 = mau_1_io_pipe_phv_out_data_390; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_391 = mau_1_io_pipe_phv_out_data_391; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_392 = mau_1_io_pipe_phv_out_data_392; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_393 = mau_1_io_pipe_phv_out_data_393; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_394 = mau_1_io_pipe_phv_out_data_394; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_395 = mau_1_io_pipe_phv_out_data_395; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_396 = mau_1_io_pipe_phv_out_data_396; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_397 = mau_1_io_pipe_phv_out_data_397; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_398 = mau_1_io_pipe_phv_out_data_398; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_399 = mau_1_io_pipe_phv_out_data_399; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_400 = mau_1_io_pipe_phv_out_data_400; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_401 = mau_1_io_pipe_phv_out_data_401; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_402 = mau_1_io_pipe_phv_out_data_402; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_403 = mau_1_io_pipe_phv_out_data_403; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_404 = mau_1_io_pipe_phv_out_data_404; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_405 = mau_1_io_pipe_phv_out_data_405; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_406 = mau_1_io_pipe_phv_out_data_406; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_407 = mau_1_io_pipe_phv_out_data_407; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_408 = mau_1_io_pipe_phv_out_data_408; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_409 = mau_1_io_pipe_phv_out_data_409; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_410 = mau_1_io_pipe_phv_out_data_410; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_411 = mau_1_io_pipe_phv_out_data_411; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_412 = mau_1_io_pipe_phv_out_data_412; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_413 = mau_1_io_pipe_phv_out_data_413; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_414 = mau_1_io_pipe_phv_out_data_414; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_415 = mau_1_io_pipe_phv_out_data_415; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_416 = mau_1_io_pipe_phv_out_data_416; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_417 = mau_1_io_pipe_phv_out_data_417; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_418 = mau_1_io_pipe_phv_out_data_418; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_419 = mau_1_io_pipe_phv_out_data_419; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_420 = mau_1_io_pipe_phv_out_data_420; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_421 = mau_1_io_pipe_phv_out_data_421; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_422 = mau_1_io_pipe_phv_out_data_422; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_423 = mau_1_io_pipe_phv_out_data_423; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_424 = mau_1_io_pipe_phv_out_data_424; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_425 = mau_1_io_pipe_phv_out_data_425; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_426 = mau_1_io_pipe_phv_out_data_426; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_427 = mau_1_io_pipe_phv_out_data_427; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_428 = mau_1_io_pipe_phv_out_data_428; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_429 = mau_1_io_pipe_phv_out_data_429; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_430 = mau_1_io_pipe_phv_out_data_430; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_431 = mau_1_io_pipe_phv_out_data_431; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_432 = mau_1_io_pipe_phv_out_data_432; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_433 = mau_1_io_pipe_phv_out_data_433; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_434 = mau_1_io_pipe_phv_out_data_434; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_435 = mau_1_io_pipe_phv_out_data_435; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_436 = mau_1_io_pipe_phv_out_data_436; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_437 = mau_1_io_pipe_phv_out_data_437; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_438 = mau_1_io_pipe_phv_out_data_438; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_439 = mau_1_io_pipe_phv_out_data_439; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_440 = mau_1_io_pipe_phv_out_data_440; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_441 = mau_1_io_pipe_phv_out_data_441; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_442 = mau_1_io_pipe_phv_out_data_442; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_443 = mau_1_io_pipe_phv_out_data_443; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_444 = mau_1_io_pipe_phv_out_data_444; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_445 = mau_1_io_pipe_phv_out_data_445; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_446 = mau_1_io_pipe_phv_out_data_446; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_447 = mau_1_io_pipe_phv_out_data_447; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_448 = mau_1_io_pipe_phv_out_data_448; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_449 = mau_1_io_pipe_phv_out_data_449; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_450 = mau_1_io_pipe_phv_out_data_450; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_451 = mau_1_io_pipe_phv_out_data_451; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_452 = mau_1_io_pipe_phv_out_data_452; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_453 = mau_1_io_pipe_phv_out_data_453; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_454 = mau_1_io_pipe_phv_out_data_454; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_455 = mau_1_io_pipe_phv_out_data_455; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_456 = mau_1_io_pipe_phv_out_data_456; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_457 = mau_1_io_pipe_phv_out_data_457; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_458 = mau_1_io_pipe_phv_out_data_458; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_459 = mau_1_io_pipe_phv_out_data_459; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_460 = mau_1_io_pipe_phv_out_data_460; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_461 = mau_1_io_pipe_phv_out_data_461; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_462 = mau_1_io_pipe_phv_out_data_462; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_463 = mau_1_io_pipe_phv_out_data_463; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_464 = mau_1_io_pipe_phv_out_data_464; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_465 = mau_1_io_pipe_phv_out_data_465; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_466 = mau_1_io_pipe_phv_out_data_466; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_467 = mau_1_io_pipe_phv_out_data_467; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_468 = mau_1_io_pipe_phv_out_data_468; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_469 = mau_1_io_pipe_phv_out_data_469; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_470 = mau_1_io_pipe_phv_out_data_470; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_471 = mau_1_io_pipe_phv_out_data_471; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_472 = mau_1_io_pipe_phv_out_data_472; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_473 = mau_1_io_pipe_phv_out_data_473; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_474 = mau_1_io_pipe_phv_out_data_474; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_475 = mau_1_io_pipe_phv_out_data_475; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_476 = mau_1_io_pipe_phv_out_data_476; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_477 = mau_1_io_pipe_phv_out_data_477; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_478 = mau_1_io_pipe_phv_out_data_478; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_479 = mau_1_io_pipe_phv_out_data_479; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_480 = mau_1_io_pipe_phv_out_data_480; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_481 = mau_1_io_pipe_phv_out_data_481; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_482 = mau_1_io_pipe_phv_out_data_482; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_483 = mau_1_io_pipe_phv_out_data_483; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_484 = mau_1_io_pipe_phv_out_data_484; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_485 = mau_1_io_pipe_phv_out_data_485; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_486 = mau_1_io_pipe_phv_out_data_486; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_487 = mau_1_io_pipe_phv_out_data_487; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_488 = mau_1_io_pipe_phv_out_data_488; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_489 = mau_1_io_pipe_phv_out_data_489; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_490 = mau_1_io_pipe_phv_out_data_490; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_491 = mau_1_io_pipe_phv_out_data_491; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_492 = mau_1_io_pipe_phv_out_data_492; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_493 = mau_1_io_pipe_phv_out_data_493; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_494 = mau_1_io_pipe_phv_out_data_494; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_495 = mau_1_io_pipe_phv_out_data_495; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_496 = mau_1_io_pipe_phv_out_data_496; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_497 = mau_1_io_pipe_phv_out_data_497; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_498 = mau_1_io_pipe_phv_out_data_498; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_499 = mau_1_io_pipe_phv_out_data_499; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_500 = mau_1_io_pipe_phv_out_data_500; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_501 = mau_1_io_pipe_phv_out_data_501; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_502 = mau_1_io_pipe_phv_out_data_502; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_503 = mau_1_io_pipe_phv_out_data_503; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_504 = mau_1_io_pipe_phv_out_data_504; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_505 = mau_1_io_pipe_phv_out_data_505; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_506 = mau_1_io_pipe_phv_out_data_506; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_507 = mau_1_io_pipe_phv_out_data_507; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_508 = mau_1_io_pipe_phv_out_data_508; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_509 = mau_1_io_pipe_phv_out_data_509; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_510 = mau_1_io_pipe_phv_out_data_510; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_data_511 = mau_1_io_pipe_phv_out_data_511; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_0 = mau_1_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_1 = mau_1_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_2 = mau_1_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_3 = mau_1_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_4 = mau_1_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_5 = mau_1_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_6 = mau_1_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_7 = mau_1_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_8 = mau_1_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_9 = mau_1_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_10 = mau_1_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_11 = mau_1_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_12 = mau_1_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_13 = mau_1_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_14 = mau_1_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_header_15 = mau_1_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_current_state = mau_1_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_current_offset = mau_1_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_parse_transition_field = mau_1_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_next_processor_id = mau_1_io_pipe_phv_out_next_processor_id; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_next_config_id = mau_1_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_2_io_pipe_phv_in_is_valid_processor = mau_1_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_2_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_2 :
    io_mod_module_mod_state_id_mod; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_2_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_2_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_2_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_2 : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_2_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_2_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  assign mau_3_clock = clock;
  assign mau_3_io_pipe_phv_in_data_0 = mau_2_io_pipe_phv_out_data_0; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_1 = mau_2_io_pipe_phv_out_data_1; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_2 = mau_2_io_pipe_phv_out_data_2; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_3 = mau_2_io_pipe_phv_out_data_3; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_4 = mau_2_io_pipe_phv_out_data_4; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_5 = mau_2_io_pipe_phv_out_data_5; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_6 = mau_2_io_pipe_phv_out_data_6; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_7 = mau_2_io_pipe_phv_out_data_7; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_8 = mau_2_io_pipe_phv_out_data_8; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_9 = mau_2_io_pipe_phv_out_data_9; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_10 = mau_2_io_pipe_phv_out_data_10; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_11 = mau_2_io_pipe_phv_out_data_11; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_12 = mau_2_io_pipe_phv_out_data_12; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_13 = mau_2_io_pipe_phv_out_data_13; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_14 = mau_2_io_pipe_phv_out_data_14; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_15 = mau_2_io_pipe_phv_out_data_15; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_16 = mau_2_io_pipe_phv_out_data_16; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_17 = mau_2_io_pipe_phv_out_data_17; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_18 = mau_2_io_pipe_phv_out_data_18; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_19 = mau_2_io_pipe_phv_out_data_19; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_20 = mau_2_io_pipe_phv_out_data_20; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_21 = mau_2_io_pipe_phv_out_data_21; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_22 = mau_2_io_pipe_phv_out_data_22; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_23 = mau_2_io_pipe_phv_out_data_23; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_24 = mau_2_io_pipe_phv_out_data_24; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_25 = mau_2_io_pipe_phv_out_data_25; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_26 = mau_2_io_pipe_phv_out_data_26; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_27 = mau_2_io_pipe_phv_out_data_27; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_28 = mau_2_io_pipe_phv_out_data_28; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_29 = mau_2_io_pipe_phv_out_data_29; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_30 = mau_2_io_pipe_phv_out_data_30; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_31 = mau_2_io_pipe_phv_out_data_31; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_32 = mau_2_io_pipe_phv_out_data_32; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_33 = mau_2_io_pipe_phv_out_data_33; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_34 = mau_2_io_pipe_phv_out_data_34; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_35 = mau_2_io_pipe_phv_out_data_35; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_36 = mau_2_io_pipe_phv_out_data_36; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_37 = mau_2_io_pipe_phv_out_data_37; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_38 = mau_2_io_pipe_phv_out_data_38; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_39 = mau_2_io_pipe_phv_out_data_39; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_40 = mau_2_io_pipe_phv_out_data_40; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_41 = mau_2_io_pipe_phv_out_data_41; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_42 = mau_2_io_pipe_phv_out_data_42; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_43 = mau_2_io_pipe_phv_out_data_43; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_44 = mau_2_io_pipe_phv_out_data_44; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_45 = mau_2_io_pipe_phv_out_data_45; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_46 = mau_2_io_pipe_phv_out_data_46; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_47 = mau_2_io_pipe_phv_out_data_47; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_48 = mau_2_io_pipe_phv_out_data_48; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_49 = mau_2_io_pipe_phv_out_data_49; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_50 = mau_2_io_pipe_phv_out_data_50; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_51 = mau_2_io_pipe_phv_out_data_51; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_52 = mau_2_io_pipe_phv_out_data_52; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_53 = mau_2_io_pipe_phv_out_data_53; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_54 = mau_2_io_pipe_phv_out_data_54; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_55 = mau_2_io_pipe_phv_out_data_55; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_56 = mau_2_io_pipe_phv_out_data_56; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_57 = mau_2_io_pipe_phv_out_data_57; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_58 = mau_2_io_pipe_phv_out_data_58; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_59 = mau_2_io_pipe_phv_out_data_59; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_60 = mau_2_io_pipe_phv_out_data_60; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_61 = mau_2_io_pipe_phv_out_data_61; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_62 = mau_2_io_pipe_phv_out_data_62; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_63 = mau_2_io_pipe_phv_out_data_63; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_64 = mau_2_io_pipe_phv_out_data_64; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_65 = mau_2_io_pipe_phv_out_data_65; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_66 = mau_2_io_pipe_phv_out_data_66; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_67 = mau_2_io_pipe_phv_out_data_67; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_68 = mau_2_io_pipe_phv_out_data_68; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_69 = mau_2_io_pipe_phv_out_data_69; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_70 = mau_2_io_pipe_phv_out_data_70; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_71 = mau_2_io_pipe_phv_out_data_71; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_72 = mau_2_io_pipe_phv_out_data_72; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_73 = mau_2_io_pipe_phv_out_data_73; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_74 = mau_2_io_pipe_phv_out_data_74; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_75 = mau_2_io_pipe_phv_out_data_75; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_76 = mau_2_io_pipe_phv_out_data_76; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_77 = mau_2_io_pipe_phv_out_data_77; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_78 = mau_2_io_pipe_phv_out_data_78; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_79 = mau_2_io_pipe_phv_out_data_79; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_80 = mau_2_io_pipe_phv_out_data_80; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_81 = mau_2_io_pipe_phv_out_data_81; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_82 = mau_2_io_pipe_phv_out_data_82; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_83 = mau_2_io_pipe_phv_out_data_83; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_84 = mau_2_io_pipe_phv_out_data_84; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_85 = mau_2_io_pipe_phv_out_data_85; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_86 = mau_2_io_pipe_phv_out_data_86; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_87 = mau_2_io_pipe_phv_out_data_87; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_88 = mau_2_io_pipe_phv_out_data_88; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_89 = mau_2_io_pipe_phv_out_data_89; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_90 = mau_2_io_pipe_phv_out_data_90; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_91 = mau_2_io_pipe_phv_out_data_91; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_92 = mau_2_io_pipe_phv_out_data_92; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_93 = mau_2_io_pipe_phv_out_data_93; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_94 = mau_2_io_pipe_phv_out_data_94; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_95 = mau_2_io_pipe_phv_out_data_95; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_96 = mau_2_io_pipe_phv_out_data_96; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_97 = mau_2_io_pipe_phv_out_data_97; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_98 = mau_2_io_pipe_phv_out_data_98; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_99 = mau_2_io_pipe_phv_out_data_99; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_100 = mau_2_io_pipe_phv_out_data_100; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_101 = mau_2_io_pipe_phv_out_data_101; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_102 = mau_2_io_pipe_phv_out_data_102; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_103 = mau_2_io_pipe_phv_out_data_103; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_104 = mau_2_io_pipe_phv_out_data_104; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_105 = mau_2_io_pipe_phv_out_data_105; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_106 = mau_2_io_pipe_phv_out_data_106; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_107 = mau_2_io_pipe_phv_out_data_107; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_108 = mau_2_io_pipe_phv_out_data_108; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_109 = mau_2_io_pipe_phv_out_data_109; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_110 = mau_2_io_pipe_phv_out_data_110; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_111 = mau_2_io_pipe_phv_out_data_111; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_112 = mau_2_io_pipe_phv_out_data_112; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_113 = mau_2_io_pipe_phv_out_data_113; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_114 = mau_2_io_pipe_phv_out_data_114; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_115 = mau_2_io_pipe_phv_out_data_115; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_116 = mau_2_io_pipe_phv_out_data_116; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_117 = mau_2_io_pipe_phv_out_data_117; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_118 = mau_2_io_pipe_phv_out_data_118; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_119 = mau_2_io_pipe_phv_out_data_119; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_120 = mau_2_io_pipe_phv_out_data_120; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_121 = mau_2_io_pipe_phv_out_data_121; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_122 = mau_2_io_pipe_phv_out_data_122; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_123 = mau_2_io_pipe_phv_out_data_123; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_124 = mau_2_io_pipe_phv_out_data_124; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_125 = mau_2_io_pipe_phv_out_data_125; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_126 = mau_2_io_pipe_phv_out_data_126; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_127 = mau_2_io_pipe_phv_out_data_127; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_128 = mau_2_io_pipe_phv_out_data_128; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_129 = mau_2_io_pipe_phv_out_data_129; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_130 = mau_2_io_pipe_phv_out_data_130; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_131 = mau_2_io_pipe_phv_out_data_131; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_132 = mau_2_io_pipe_phv_out_data_132; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_133 = mau_2_io_pipe_phv_out_data_133; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_134 = mau_2_io_pipe_phv_out_data_134; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_135 = mau_2_io_pipe_phv_out_data_135; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_136 = mau_2_io_pipe_phv_out_data_136; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_137 = mau_2_io_pipe_phv_out_data_137; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_138 = mau_2_io_pipe_phv_out_data_138; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_139 = mau_2_io_pipe_phv_out_data_139; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_140 = mau_2_io_pipe_phv_out_data_140; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_141 = mau_2_io_pipe_phv_out_data_141; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_142 = mau_2_io_pipe_phv_out_data_142; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_143 = mau_2_io_pipe_phv_out_data_143; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_144 = mau_2_io_pipe_phv_out_data_144; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_145 = mau_2_io_pipe_phv_out_data_145; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_146 = mau_2_io_pipe_phv_out_data_146; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_147 = mau_2_io_pipe_phv_out_data_147; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_148 = mau_2_io_pipe_phv_out_data_148; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_149 = mau_2_io_pipe_phv_out_data_149; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_150 = mau_2_io_pipe_phv_out_data_150; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_151 = mau_2_io_pipe_phv_out_data_151; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_152 = mau_2_io_pipe_phv_out_data_152; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_153 = mau_2_io_pipe_phv_out_data_153; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_154 = mau_2_io_pipe_phv_out_data_154; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_155 = mau_2_io_pipe_phv_out_data_155; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_156 = mau_2_io_pipe_phv_out_data_156; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_157 = mau_2_io_pipe_phv_out_data_157; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_158 = mau_2_io_pipe_phv_out_data_158; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_159 = mau_2_io_pipe_phv_out_data_159; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_160 = mau_2_io_pipe_phv_out_data_160; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_161 = mau_2_io_pipe_phv_out_data_161; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_162 = mau_2_io_pipe_phv_out_data_162; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_163 = mau_2_io_pipe_phv_out_data_163; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_164 = mau_2_io_pipe_phv_out_data_164; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_165 = mau_2_io_pipe_phv_out_data_165; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_166 = mau_2_io_pipe_phv_out_data_166; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_167 = mau_2_io_pipe_phv_out_data_167; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_168 = mau_2_io_pipe_phv_out_data_168; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_169 = mau_2_io_pipe_phv_out_data_169; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_170 = mau_2_io_pipe_phv_out_data_170; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_171 = mau_2_io_pipe_phv_out_data_171; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_172 = mau_2_io_pipe_phv_out_data_172; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_173 = mau_2_io_pipe_phv_out_data_173; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_174 = mau_2_io_pipe_phv_out_data_174; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_175 = mau_2_io_pipe_phv_out_data_175; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_176 = mau_2_io_pipe_phv_out_data_176; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_177 = mau_2_io_pipe_phv_out_data_177; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_178 = mau_2_io_pipe_phv_out_data_178; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_179 = mau_2_io_pipe_phv_out_data_179; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_180 = mau_2_io_pipe_phv_out_data_180; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_181 = mau_2_io_pipe_phv_out_data_181; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_182 = mau_2_io_pipe_phv_out_data_182; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_183 = mau_2_io_pipe_phv_out_data_183; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_184 = mau_2_io_pipe_phv_out_data_184; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_185 = mau_2_io_pipe_phv_out_data_185; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_186 = mau_2_io_pipe_phv_out_data_186; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_187 = mau_2_io_pipe_phv_out_data_187; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_188 = mau_2_io_pipe_phv_out_data_188; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_189 = mau_2_io_pipe_phv_out_data_189; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_190 = mau_2_io_pipe_phv_out_data_190; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_191 = mau_2_io_pipe_phv_out_data_191; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_192 = mau_2_io_pipe_phv_out_data_192; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_193 = mau_2_io_pipe_phv_out_data_193; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_194 = mau_2_io_pipe_phv_out_data_194; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_195 = mau_2_io_pipe_phv_out_data_195; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_196 = mau_2_io_pipe_phv_out_data_196; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_197 = mau_2_io_pipe_phv_out_data_197; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_198 = mau_2_io_pipe_phv_out_data_198; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_199 = mau_2_io_pipe_phv_out_data_199; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_200 = mau_2_io_pipe_phv_out_data_200; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_201 = mau_2_io_pipe_phv_out_data_201; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_202 = mau_2_io_pipe_phv_out_data_202; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_203 = mau_2_io_pipe_phv_out_data_203; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_204 = mau_2_io_pipe_phv_out_data_204; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_205 = mau_2_io_pipe_phv_out_data_205; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_206 = mau_2_io_pipe_phv_out_data_206; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_207 = mau_2_io_pipe_phv_out_data_207; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_208 = mau_2_io_pipe_phv_out_data_208; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_209 = mau_2_io_pipe_phv_out_data_209; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_210 = mau_2_io_pipe_phv_out_data_210; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_211 = mau_2_io_pipe_phv_out_data_211; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_212 = mau_2_io_pipe_phv_out_data_212; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_213 = mau_2_io_pipe_phv_out_data_213; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_214 = mau_2_io_pipe_phv_out_data_214; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_215 = mau_2_io_pipe_phv_out_data_215; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_216 = mau_2_io_pipe_phv_out_data_216; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_217 = mau_2_io_pipe_phv_out_data_217; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_218 = mau_2_io_pipe_phv_out_data_218; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_219 = mau_2_io_pipe_phv_out_data_219; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_220 = mau_2_io_pipe_phv_out_data_220; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_221 = mau_2_io_pipe_phv_out_data_221; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_222 = mau_2_io_pipe_phv_out_data_222; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_223 = mau_2_io_pipe_phv_out_data_223; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_224 = mau_2_io_pipe_phv_out_data_224; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_225 = mau_2_io_pipe_phv_out_data_225; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_226 = mau_2_io_pipe_phv_out_data_226; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_227 = mau_2_io_pipe_phv_out_data_227; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_228 = mau_2_io_pipe_phv_out_data_228; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_229 = mau_2_io_pipe_phv_out_data_229; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_230 = mau_2_io_pipe_phv_out_data_230; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_231 = mau_2_io_pipe_phv_out_data_231; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_232 = mau_2_io_pipe_phv_out_data_232; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_233 = mau_2_io_pipe_phv_out_data_233; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_234 = mau_2_io_pipe_phv_out_data_234; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_235 = mau_2_io_pipe_phv_out_data_235; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_236 = mau_2_io_pipe_phv_out_data_236; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_237 = mau_2_io_pipe_phv_out_data_237; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_238 = mau_2_io_pipe_phv_out_data_238; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_239 = mau_2_io_pipe_phv_out_data_239; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_240 = mau_2_io_pipe_phv_out_data_240; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_241 = mau_2_io_pipe_phv_out_data_241; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_242 = mau_2_io_pipe_phv_out_data_242; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_243 = mau_2_io_pipe_phv_out_data_243; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_244 = mau_2_io_pipe_phv_out_data_244; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_245 = mau_2_io_pipe_phv_out_data_245; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_246 = mau_2_io_pipe_phv_out_data_246; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_247 = mau_2_io_pipe_phv_out_data_247; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_248 = mau_2_io_pipe_phv_out_data_248; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_249 = mau_2_io_pipe_phv_out_data_249; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_250 = mau_2_io_pipe_phv_out_data_250; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_251 = mau_2_io_pipe_phv_out_data_251; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_252 = mau_2_io_pipe_phv_out_data_252; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_253 = mau_2_io_pipe_phv_out_data_253; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_254 = mau_2_io_pipe_phv_out_data_254; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_255 = mau_2_io_pipe_phv_out_data_255; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_256 = mau_2_io_pipe_phv_out_data_256; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_257 = mau_2_io_pipe_phv_out_data_257; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_258 = mau_2_io_pipe_phv_out_data_258; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_259 = mau_2_io_pipe_phv_out_data_259; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_260 = mau_2_io_pipe_phv_out_data_260; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_261 = mau_2_io_pipe_phv_out_data_261; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_262 = mau_2_io_pipe_phv_out_data_262; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_263 = mau_2_io_pipe_phv_out_data_263; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_264 = mau_2_io_pipe_phv_out_data_264; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_265 = mau_2_io_pipe_phv_out_data_265; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_266 = mau_2_io_pipe_phv_out_data_266; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_267 = mau_2_io_pipe_phv_out_data_267; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_268 = mau_2_io_pipe_phv_out_data_268; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_269 = mau_2_io_pipe_phv_out_data_269; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_270 = mau_2_io_pipe_phv_out_data_270; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_271 = mau_2_io_pipe_phv_out_data_271; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_272 = mau_2_io_pipe_phv_out_data_272; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_273 = mau_2_io_pipe_phv_out_data_273; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_274 = mau_2_io_pipe_phv_out_data_274; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_275 = mau_2_io_pipe_phv_out_data_275; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_276 = mau_2_io_pipe_phv_out_data_276; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_277 = mau_2_io_pipe_phv_out_data_277; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_278 = mau_2_io_pipe_phv_out_data_278; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_279 = mau_2_io_pipe_phv_out_data_279; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_280 = mau_2_io_pipe_phv_out_data_280; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_281 = mau_2_io_pipe_phv_out_data_281; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_282 = mau_2_io_pipe_phv_out_data_282; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_283 = mau_2_io_pipe_phv_out_data_283; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_284 = mau_2_io_pipe_phv_out_data_284; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_285 = mau_2_io_pipe_phv_out_data_285; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_286 = mau_2_io_pipe_phv_out_data_286; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_287 = mau_2_io_pipe_phv_out_data_287; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_288 = mau_2_io_pipe_phv_out_data_288; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_289 = mau_2_io_pipe_phv_out_data_289; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_290 = mau_2_io_pipe_phv_out_data_290; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_291 = mau_2_io_pipe_phv_out_data_291; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_292 = mau_2_io_pipe_phv_out_data_292; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_293 = mau_2_io_pipe_phv_out_data_293; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_294 = mau_2_io_pipe_phv_out_data_294; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_295 = mau_2_io_pipe_phv_out_data_295; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_296 = mau_2_io_pipe_phv_out_data_296; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_297 = mau_2_io_pipe_phv_out_data_297; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_298 = mau_2_io_pipe_phv_out_data_298; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_299 = mau_2_io_pipe_phv_out_data_299; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_300 = mau_2_io_pipe_phv_out_data_300; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_301 = mau_2_io_pipe_phv_out_data_301; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_302 = mau_2_io_pipe_phv_out_data_302; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_303 = mau_2_io_pipe_phv_out_data_303; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_304 = mau_2_io_pipe_phv_out_data_304; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_305 = mau_2_io_pipe_phv_out_data_305; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_306 = mau_2_io_pipe_phv_out_data_306; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_307 = mau_2_io_pipe_phv_out_data_307; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_308 = mau_2_io_pipe_phv_out_data_308; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_309 = mau_2_io_pipe_phv_out_data_309; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_310 = mau_2_io_pipe_phv_out_data_310; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_311 = mau_2_io_pipe_phv_out_data_311; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_312 = mau_2_io_pipe_phv_out_data_312; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_313 = mau_2_io_pipe_phv_out_data_313; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_314 = mau_2_io_pipe_phv_out_data_314; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_315 = mau_2_io_pipe_phv_out_data_315; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_316 = mau_2_io_pipe_phv_out_data_316; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_317 = mau_2_io_pipe_phv_out_data_317; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_318 = mau_2_io_pipe_phv_out_data_318; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_319 = mau_2_io_pipe_phv_out_data_319; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_320 = mau_2_io_pipe_phv_out_data_320; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_321 = mau_2_io_pipe_phv_out_data_321; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_322 = mau_2_io_pipe_phv_out_data_322; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_323 = mau_2_io_pipe_phv_out_data_323; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_324 = mau_2_io_pipe_phv_out_data_324; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_325 = mau_2_io_pipe_phv_out_data_325; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_326 = mau_2_io_pipe_phv_out_data_326; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_327 = mau_2_io_pipe_phv_out_data_327; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_328 = mau_2_io_pipe_phv_out_data_328; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_329 = mau_2_io_pipe_phv_out_data_329; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_330 = mau_2_io_pipe_phv_out_data_330; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_331 = mau_2_io_pipe_phv_out_data_331; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_332 = mau_2_io_pipe_phv_out_data_332; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_333 = mau_2_io_pipe_phv_out_data_333; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_334 = mau_2_io_pipe_phv_out_data_334; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_335 = mau_2_io_pipe_phv_out_data_335; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_336 = mau_2_io_pipe_phv_out_data_336; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_337 = mau_2_io_pipe_phv_out_data_337; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_338 = mau_2_io_pipe_phv_out_data_338; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_339 = mau_2_io_pipe_phv_out_data_339; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_340 = mau_2_io_pipe_phv_out_data_340; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_341 = mau_2_io_pipe_phv_out_data_341; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_342 = mau_2_io_pipe_phv_out_data_342; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_343 = mau_2_io_pipe_phv_out_data_343; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_344 = mau_2_io_pipe_phv_out_data_344; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_345 = mau_2_io_pipe_phv_out_data_345; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_346 = mau_2_io_pipe_phv_out_data_346; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_347 = mau_2_io_pipe_phv_out_data_347; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_348 = mau_2_io_pipe_phv_out_data_348; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_349 = mau_2_io_pipe_phv_out_data_349; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_350 = mau_2_io_pipe_phv_out_data_350; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_351 = mau_2_io_pipe_phv_out_data_351; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_352 = mau_2_io_pipe_phv_out_data_352; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_353 = mau_2_io_pipe_phv_out_data_353; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_354 = mau_2_io_pipe_phv_out_data_354; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_355 = mau_2_io_pipe_phv_out_data_355; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_356 = mau_2_io_pipe_phv_out_data_356; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_357 = mau_2_io_pipe_phv_out_data_357; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_358 = mau_2_io_pipe_phv_out_data_358; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_359 = mau_2_io_pipe_phv_out_data_359; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_360 = mau_2_io_pipe_phv_out_data_360; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_361 = mau_2_io_pipe_phv_out_data_361; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_362 = mau_2_io_pipe_phv_out_data_362; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_363 = mau_2_io_pipe_phv_out_data_363; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_364 = mau_2_io_pipe_phv_out_data_364; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_365 = mau_2_io_pipe_phv_out_data_365; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_366 = mau_2_io_pipe_phv_out_data_366; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_367 = mau_2_io_pipe_phv_out_data_367; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_368 = mau_2_io_pipe_phv_out_data_368; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_369 = mau_2_io_pipe_phv_out_data_369; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_370 = mau_2_io_pipe_phv_out_data_370; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_371 = mau_2_io_pipe_phv_out_data_371; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_372 = mau_2_io_pipe_phv_out_data_372; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_373 = mau_2_io_pipe_phv_out_data_373; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_374 = mau_2_io_pipe_phv_out_data_374; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_375 = mau_2_io_pipe_phv_out_data_375; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_376 = mau_2_io_pipe_phv_out_data_376; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_377 = mau_2_io_pipe_phv_out_data_377; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_378 = mau_2_io_pipe_phv_out_data_378; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_379 = mau_2_io_pipe_phv_out_data_379; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_380 = mau_2_io_pipe_phv_out_data_380; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_381 = mau_2_io_pipe_phv_out_data_381; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_382 = mau_2_io_pipe_phv_out_data_382; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_383 = mau_2_io_pipe_phv_out_data_383; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_384 = mau_2_io_pipe_phv_out_data_384; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_385 = mau_2_io_pipe_phv_out_data_385; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_386 = mau_2_io_pipe_phv_out_data_386; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_387 = mau_2_io_pipe_phv_out_data_387; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_388 = mau_2_io_pipe_phv_out_data_388; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_389 = mau_2_io_pipe_phv_out_data_389; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_390 = mau_2_io_pipe_phv_out_data_390; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_391 = mau_2_io_pipe_phv_out_data_391; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_392 = mau_2_io_pipe_phv_out_data_392; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_393 = mau_2_io_pipe_phv_out_data_393; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_394 = mau_2_io_pipe_phv_out_data_394; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_395 = mau_2_io_pipe_phv_out_data_395; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_396 = mau_2_io_pipe_phv_out_data_396; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_397 = mau_2_io_pipe_phv_out_data_397; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_398 = mau_2_io_pipe_phv_out_data_398; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_399 = mau_2_io_pipe_phv_out_data_399; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_400 = mau_2_io_pipe_phv_out_data_400; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_401 = mau_2_io_pipe_phv_out_data_401; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_402 = mau_2_io_pipe_phv_out_data_402; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_403 = mau_2_io_pipe_phv_out_data_403; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_404 = mau_2_io_pipe_phv_out_data_404; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_405 = mau_2_io_pipe_phv_out_data_405; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_406 = mau_2_io_pipe_phv_out_data_406; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_407 = mau_2_io_pipe_phv_out_data_407; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_408 = mau_2_io_pipe_phv_out_data_408; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_409 = mau_2_io_pipe_phv_out_data_409; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_410 = mau_2_io_pipe_phv_out_data_410; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_411 = mau_2_io_pipe_phv_out_data_411; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_412 = mau_2_io_pipe_phv_out_data_412; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_413 = mau_2_io_pipe_phv_out_data_413; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_414 = mau_2_io_pipe_phv_out_data_414; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_415 = mau_2_io_pipe_phv_out_data_415; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_416 = mau_2_io_pipe_phv_out_data_416; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_417 = mau_2_io_pipe_phv_out_data_417; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_418 = mau_2_io_pipe_phv_out_data_418; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_419 = mau_2_io_pipe_phv_out_data_419; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_420 = mau_2_io_pipe_phv_out_data_420; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_421 = mau_2_io_pipe_phv_out_data_421; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_422 = mau_2_io_pipe_phv_out_data_422; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_423 = mau_2_io_pipe_phv_out_data_423; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_424 = mau_2_io_pipe_phv_out_data_424; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_425 = mau_2_io_pipe_phv_out_data_425; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_426 = mau_2_io_pipe_phv_out_data_426; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_427 = mau_2_io_pipe_phv_out_data_427; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_428 = mau_2_io_pipe_phv_out_data_428; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_429 = mau_2_io_pipe_phv_out_data_429; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_430 = mau_2_io_pipe_phv_out_data_430; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_431 = mau_2_io_pipe_phv_out_data_431; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_432 = mau_2_io_pipe_phv_out_data_432; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_433 = mau_2_io_pipe_phv_out_data_433; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_434 = mau_2_io_pipe_phv_out_data_434; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_435 = mau_2_io_pipe_phv_out_data_435; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_436 = mau_2_io_pipe_phv_out_data_436; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_437 = mau_2_io_pipe_phv_out_data_437; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_438 = mau_2_io_pipe_phv_out_data_438; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_439 = mau_2_io_pipe_phv_out_data_439; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_440 = mau_2_io_pipe_phv_out_data_440; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_441 = mau_2_io_pipe_phv_out_data_441; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_442 = mau_2_io_pipe_phv_out_data_442; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_443 = mau_2_io_pipe_phv_out_data_443; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_444 = mau_2_io_pipe_phv_out_data_444; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_445 = mau_2_io_pipe_phv_out_data_445; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_446 = mau_2_io_pipe_phv_out_data_446; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_447 = mau_2_io_pipe_phv_out_data_447; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_448 = mau_2_io_pipe_phv_out_data_448; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_449 = mau_2_io_pipe_phv_out_data_449; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_450 = mau_2_io_pipe_phv_out_data_450; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_451 = mau_2_io_pipe_phv_out_data_451; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_452 = mau_2_io_pipe_phv_out_data_452; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_453 = mau_2_io_pipe_phv_out_data_453; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_454 = mau_2_io_pipe_phv_out_data_454; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_455 = mau_2_io_pipe_phv_out_data_455; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_456 = mau_2_io_pipe_phv_out_data_456; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_457 = mau_2_io_pipe_phv_out_data_457; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_458 = mau_2_io_pipe_phv_out_data_458; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_459 = mau_2_io_pipe_phv_out_data_459; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_460 = mau_2_io_pipe_phv_out_data_460; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_461 = mau_2_io_pipe_phv_out_data_461; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_462 = mau_2_io_pipe_phv_out_data_462; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_463 = mau_2_io_pipe_phv_out_data_463; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_464 = mau_2_io_pipe_phv_out_data_464; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_465 = mau_2_io_pipe_phv_out_data_465; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_466 = mau_2_io_pipe_phv_out_data_466; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_467 = mau_2_io_pipe_phv_out_data_467; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_468 = mau_2_io_pipe_phv_out_data_468; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_469 = mau_2_io_pipe_phv_out_data_469; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_470 = mau_2_io_pipe_phv_out_data_470; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_471 = mau_2_io_pipe_phv_out_data_471; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_472 = mau_2_io_pipe_phv_out_data_472; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_473 = mau_2_io_pipe_phv_out_data_473; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_474 = mau_2_io_pipe_phv_out_data_474; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_475 = mau_2_io_pipe_phv_out_data_475; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_476 = mau_2_io_pipe_phv_out_data_476; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_477 = mau_2_io_pipe_phv_out_data_477; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_478 = mau_2_io_pipe_phv_out_data_478; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_479 = mau_2_io_pipe_phv_out_data_479; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_480 = mau_2_io_pipe_phv_out_data_480; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_481 = mau_2_io_pipe_phv_out_data_481; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_482 = mau_2_io_pipe_phv_out_data_482; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_483 = mau_2_io_pipe_phv_out_data_483; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_484 = mau_2_io_pipe_phv_out_data_484; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_485 = mau_2_io_pipe_phv_out_data_485; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_486 = mau_2_io_pipe_phv_out_data_486; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_487 = mau_2_io_pipe_phv_out_data_487; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_488 = mau_2_io_pipe_phv_out_data_488; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_489 = mau_2_io_pipe_phv_out_data_489; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_490 = mau_2_io_pipe_phv_out_data_490; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_491 = mau_2_io_pipe_phv_out_data_491; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_492 = mau_2_io_pipe_phv_out_data_492; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_493 = mau_2_io_pipe_phv_out_data_493; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_494 = mau_2_io_pipe_phv_out_data_494; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_495 = mau_2_io_pipe_phv_out_data_495; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_496 = mau_2_io_pipe_phv_out_data_496; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_497 = mau_2_io_pipe_phv_out_data_497; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_498 = mau_2_io_pipe_phv_out_data_498; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_499 = mau_2_io_pipe_phv_out_data_499; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_500 = mau_2_io_pipe_phv_out_data_500; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_501 = mau_2_io_pipe_phv_out_data_501; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_502 = mau_2_io_pipe_phv_out_data_502; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_503 = mau_2_io_pipe_phv_out_data_503; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_504 = mau_2_io_pipe_phv_out_data_504; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_505 = mau_2_io_pipe_phv_out_data_505; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_506 = mau_2_io_pipe_phv_out_data_506; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_507 = mau_2_io_pipe_phv_out_data_507; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_508 = mau_2_io_pipe_phv_out_data_508; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_509 = mau_2_io_pipe_phv_out_data_509; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_510 = mau_2_io_pipe_phv_out_data_510; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_data_511 = mau_2_io_pipe_phv_out_data_511; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_0 = mau_2_io_pipe_phv_out_header_0; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_1 = mau_2_io_pipe_phv_out_header_1; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_2 = mau_2_io_pipe_phv_out_header_2; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_3 = mau_2_io_pipe_phv_out_header_3; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_4 = mau_2_io_pipe_phv_out_header_4; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_5 = mau_2_io_pipe_phv_out_header_5; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_6 = mau_2_io_pipe_phv_out_header_6; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_7 = mau_2_io_pipe_phv_out_header_7; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_8 = mau_2_io_pipe_phv_out_header_8; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_9 = mau_2_io_pipe_phv_out_header_9; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_10 = mau_2_io_pipe_phv_out_header_10; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_11 = mau_2_io_pipe_phv_out_header_11; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_12 = mau_2_io_pipe_phv_out_header_12; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_13 = mau_2_io_pipe_phv_out_header_13; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_14 = mau_2_io_pipe_phv_out_header_14; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_header_15 = mau_2_io_pipe_phv_out_header_15; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_current_state = mau_2_io_pipe_phv_out_parse_current_state; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_current_offset = mau_2_io_pipe_phv_out_parse_current_offset; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_parse_transition_field = mau_2_io_pipe_phv_out_parse_transition_field; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_next_processor_id = mau_2_io_pipe_phv_out_next_processor_id; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_next_config_id = mau_2_io_pipe_phv_out_next_config_id; // @[parser.scala 32:35]
  assign mau_3_io_pipe_phv_in_is_valid_processor = mau_2_io_pipe_phv_out_is_valid_processor; // @[parser.scala 32:35]
  assign mau_3_io_mod_state_id_mod = io_mod_en ? io_mod_module_mod_state_id_mod & mod_j_3 :
    io_mod_module_mod_state_id_mod; // @[parser.scala 41:22 parser.scala 48:40 parser.scala 37:23]
  assign mau_3_io_mod_state_id = io_mod_module_mod_state_id; // @[parser.scala 37:23]
  assign mau_3_io_mod_sram_w_cs = io_mod_module_mod_sram_w_cs; // @[parser.scala 37:23]
  assign mau_3_io_mod_sram_w_en = io_mod_en ? io_mod_module_mod_sram_w_en & mod_j_3 : io_mod_module_mod_sram_w_en; // @[parser.scala 41:22 parser.scala 47:40 parser.scala 37:23]
  assign mau_3_io_mod_sram_w_addr = io_mod_module_mod_sram_w_addr; // @[parser.scala 37:23]
  assign mau_3_io_mod_sram_w_data = io_mod_module_mod_sram_w_data; // @[parser.scala 37:23]
  always @(posedge clock) begin
    if (io_mod_en) begin // @[parser.scala 41:22]
      if (io_mod_last_mau_id_mod) begin // @[parser.scala 42:39]
        last_mau_id <= {{1'd0}, io_mod_last_mau_id}; // @[parser.scala 43:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  last_mau_id = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
