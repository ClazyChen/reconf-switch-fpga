module Matcher(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  input         io_pipe_phv_in_valid,
  input         io_pipe_phv_in_last,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  output        io_pipe_phv_out_valid,
  output        io_pipe_phv_out_last
);
  wire  pipe1_clock; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 343:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_valid; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_in_last; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 343:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 343:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 343:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_valid; // @[matcher.scala 343:23]
  wire  pipe1_io_pipe_phv_out_last; // @[matcher.scala 343:23]
  wire  pipe2_clock; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 344:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_valid; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_in_last; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 344:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 344:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 344:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_valid; // @[matcher.scala 344:23]
  wire  pipe2_io_pipe_phv_out_last; // @[matcher.scala 344:23]
  wire  pipe3to8_clock; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_0; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_1; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_2; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_3; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_4; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_5; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_6; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_7; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_8; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_9; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_10; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_11; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_12; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_13; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_14; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_16; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_17; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_18; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_19; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_20; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_21; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_22; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_23; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_24; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_25; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_26; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_27; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_28; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_29; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_30; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_31; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_32; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_33; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_34; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_35; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_36; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_37; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_38; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_39; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_40; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_41; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_42; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_43; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_44; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_45; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_46; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_47; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_48; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_49; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_50; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_51; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_52; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_53; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_54; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_55; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_56; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_57; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_58; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_59; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_60; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_61; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_62; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_63; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_64; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_65; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_66; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_67; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_68; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_69; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_70; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_71; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_72; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_73; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_74; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_75; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_76; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_77; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_78; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_79; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_80; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_81; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_82; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_83; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_84; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_85; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_86; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_87; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_88; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_89; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_90; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_91; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_92; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_93; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_94; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_95; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_96; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_97; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_98; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_99; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_100; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_101; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_102; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_103; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_104; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_105; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_106; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_107; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_108; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_109; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_110; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_111; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_112; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_113; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_114; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_115; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_116; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_117; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_118; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_119; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_120; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_121; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_122; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_123; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_124; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_125; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_126; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_127; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_128; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_129; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_130; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_131; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_132; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_133; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_134; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_135; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_136; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_137; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_138; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_139; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_140; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_141; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_142; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_143; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_144; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_145; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_146; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_147; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_148; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_149; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_150; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_151; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_152; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_153; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_154; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_155; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_156; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_157; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_158; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_data_159; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_0; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_1; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_2; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_3; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_4; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_5; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_6; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_7; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_8; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_9; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_10; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_11; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_12; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_13; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_14; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_header_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_state; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 345:26]
  wire [3:0] pipe3to8_io_pipe_phv_in_next_processor_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_next_config_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_valid; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_in_last; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_96; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_97; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_98; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_99; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_100; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_101; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_102; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_103; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_104; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_105; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_106; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_107; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_108; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_109; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_110; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_111; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_112; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_113; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_114; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_115; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_116; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_117; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_118; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_119; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_120; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_121; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_122; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_123; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_124; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_125; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_126; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_127; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_128; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_129; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_130; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_131; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_132; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_133; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_134; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_135; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_136; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_137; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_138; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_139; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_140; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_141; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_142; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_143; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_144; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_145; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_146; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_147; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_148; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_149; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_150; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_151; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_152; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_153; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_154; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_155; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_156; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_157; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_158; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_data_159; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 345:26]
  wire [7:0] pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 345:26]
  wire [15:0] pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 345:26]
  wire [3:0] pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_valid; // @[matcher.scala 345:26]
  wire  pipe3to8_io_pipe_phv_out_last; // @[matcher.scala 345:26]
  wire  pipe9_clock; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_0; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_1; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_2; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_3; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_4; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_5; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_6; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_7; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_8; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_9; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_10; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_11; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_12; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_13; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_14; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_16; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_17; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_18; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_19; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_20; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_21; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_22; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_23; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_24; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_25; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_26; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_27; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_28; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_29; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_30; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_31; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_32; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_33; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_34; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_35; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_36; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_37; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_38; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_39; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_40; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_41; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_42; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_43; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_44; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_45; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_46; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_47; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_48; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_49; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_50; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_51; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_52; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_53; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_54; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_55; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_56; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_57; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_58; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_59; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_60; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_61; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_62; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_63; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_64; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_65; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_66; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_67; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_68; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_69; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_70; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_71; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_72; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_73; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_74; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_75; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_76; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_77; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_78; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_79; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_80; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_81; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_82; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_83; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_84; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_85; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_86; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_87; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_88; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_89; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_90; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_91; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_92; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_93; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_94; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_95; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_96; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_97; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_98; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_99; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_100; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_101; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_102; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_103; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_104; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_105; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_106; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_107; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_108; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_109; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_110; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_111; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_112; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_113; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_114; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_115; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_116; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_117; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_118; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_119; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_120; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_121; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_122; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_123; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_124; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_125; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_126; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_127; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_128; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_129; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_130; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_131; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_132; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_133; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_134; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_135; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_136; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_137; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_138; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_139; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_140; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_141; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_142; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_143; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_144; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_145; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_146; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_147; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_148; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_149; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_150; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_151; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_152; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_153; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_154; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_155; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_156; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_157; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_158; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_data_159; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_0; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_1; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_2; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_3; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_4; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_5; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_6; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_7; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_8; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_9; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_10; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_11; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_12; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_13; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_14; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_header_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_state; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 346:23]
  wire [3:0] pipe9_io_pipe_phv_in_next_processor_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_next_config_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_valid; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_in_last; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_96; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_97; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_98; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_99; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_100; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_101; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_102; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_103; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_104; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_105; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_106; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_107; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_108; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_109; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_110; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_111; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_112; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_113; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_114; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_115; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_116; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_117; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_118; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_119; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_120; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_121; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_122; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_123; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_124; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_125; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_126; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_127; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_128; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_129; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_130; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_131; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_132; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_133; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_134; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_135; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_136; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_137; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_138; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_139; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_140; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_141; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_142; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_143; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_144; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_145; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_146; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_147; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_148; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_149; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_150; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_151; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_152; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_153; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_154; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_155; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_156; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_157; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_158; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_data_159; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 346:23]
  wire [7:0] pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 346:23]
  wire [15:0] pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 346:23]
  wire [3:0] pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_valid; // @[matcher.scala 346:23]
  wire  pipe9_io_pipe_phv_out_last; // @[matcher.scala 346:23]
  wire  pipe10_clock; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_0; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_1; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_2; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_3; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_4; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_5; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_6; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_7; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_8; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_9; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_10; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_11; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_12; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_13; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_14; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_16; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_17; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_18; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_19; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_20; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_21; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_22; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_23; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_24; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_25; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_26; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_27; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_28; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_29; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_30; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_31; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_32; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_33; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_34; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_35; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_36; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_37; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_38; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_39; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_40; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_41; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_42; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_43; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_44; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_45; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_46; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_47; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_48; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_49; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_50; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_51; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_52; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_53; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_54; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_55; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_56; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_57; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_58; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_59; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_60; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_61; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_62; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_63; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_64; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_65; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_66; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_67; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_68; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_69; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_70; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_71; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_72; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_73; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_74; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_75; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_76; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_77; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_78; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_79; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_80; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_81; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_82; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_83; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_84; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_85; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_86; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_87; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_88; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_89; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_90; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_91; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_92; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_93; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_94; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_95; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_96; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_97; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_98; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_99; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_100; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_101; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_102; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_103; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_104; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_105; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_106; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_107; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_108; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_109; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_110; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_111; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_112; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_113; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_114; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_115; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_116; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_117; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_118; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_119; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_120; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_121; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_122; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_123; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_124; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_125; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_126; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_127; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_128; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_129; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_130; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_131; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_132; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_133; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_134; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_135; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_136; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_137; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_138; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_139; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_140; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_141; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_142; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_143; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_144; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_145; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_146; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_147; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_148; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_149; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_150; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_151; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_152; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_153; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_154; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_155; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_156; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_157; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_158; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_data_159; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_0; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_1; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_2; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_3; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_4; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_5; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_6; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_7; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_8; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_9; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_10; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_11; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_12; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_13; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_14; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_header_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_state; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 347:24]
  wire [3:0] pipe10_io_pipe_phv_in_next_processor_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_next_config_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_valid; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_in_last; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_96; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_97; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_98; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_99; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_100; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_101; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_102; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_103; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_104; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_105; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_106; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_107; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_108; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_109; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_110; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_111; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_112; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_113; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_114; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_115; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_116; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_117; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_118; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_119; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_120; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_121; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_122; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_123; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_124; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_125; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_126; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_127; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_128; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_129; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_130; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_131; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_132; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_133; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_134; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_135; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_136; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_137; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_138; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_139; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_140; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_141; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_142; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_143; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_144; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_145; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_146; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_147; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_148; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_149; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_150; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_151; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_152; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_153; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_154; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_155; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_156; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_157; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_158; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_data_159; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 347:24]
  wire [7:0] pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 347:24]
  wire [15:0] pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 347:24]
  wire [3:0] pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_valid; // @[matcher.scala 347:24]
  wire  pipe10_io_pipe_phv_out_last; // @[matcher.scala 347:24]
  wire  pipe11_clock; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_0; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_1; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_2; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_3; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_4; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_5; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_6; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_7; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_8; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_9; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_10; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_11; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_12; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_13; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_14; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_16; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_17; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_18; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_19; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_20; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_21; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_22; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_23; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_24; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_25; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_26; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_27; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_28; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_29; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_30; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_31; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_32; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_33; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_34; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_35; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_36; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_37; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_38; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_39; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_40; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_41; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_42; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_43; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_44; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_45; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_46; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_47; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_48; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_49; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_50; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_51; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_52; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_53; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_54; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_55; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_56; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_57; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_58; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_59; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_60; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_61; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_62; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_63; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_64; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_65; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_66; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_67; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_68; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_69; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_70; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_71; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_72; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_73; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_74; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_75; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_76; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_77; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_78; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_79; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_80; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_81; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_82; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_83; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_84; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_85; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_86; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_87; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_88; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_89; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_90; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_91; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_92; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_93; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_94; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_95; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_96; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_97; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_98; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_99; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_100; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_101; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_102; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_103; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_104; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_105; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_106; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_107; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_108; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_109; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_110; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_111; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_112; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_113; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_114; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_115; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_116; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_117; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_118; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_119; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_120; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_121; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_122; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_123; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_124; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_125; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_126; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_127; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_128; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_129; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_130; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_131; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_132; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_133; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_134; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_135; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_136; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_137; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_138; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_139; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_140; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_141; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_142; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_143; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_144; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_145; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_146; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_147; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_148; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_149; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_150; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_151; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_152; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_153; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_154; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_155; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_156; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_157; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_158; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_data_159; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_0; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_1; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_2; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_3; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_4; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_5; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_6; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_7; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_8; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_9; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_10; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_11; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_12; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_13; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_14; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_header_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_state; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 348:24]
  wire [3:0] pipe11_io_pipe_phv_in_next_processor_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_next_config_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_valid; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_in_last; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_96; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_97; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_98; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_99; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_100; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_101; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_102; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_103; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_104; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_105; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_106; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_107; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_108; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_109; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_110; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_111; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_112; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_113; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_114; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_115; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_116; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_117; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_118; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_119; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_120; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_121; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_122; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_123; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_124; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_125; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_126; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_127; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_128; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_129; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_130; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_131; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_132; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_133; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_134; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_135; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_136; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_137; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_138; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_139; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_140; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_141; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_142; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_143; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_144; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_145; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_146; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_147; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_148; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_149; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_150; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_151; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_152; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_153; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_154; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_155; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_156; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_157; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_158; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_data_159; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 348:24]
  wire [7:0] pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 348:24]
  wire [15:0] pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 348:24]
  wire [3:0] pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_valid; // @[matcher.scala 348:24]
  wire  pipe11_io_pipe_phv_out_last; // @[matcher.scala 348:24]
  wire  pipe12_clock; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_0; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_1; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_2; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_3; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_4; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_5; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_6; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_7; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_8; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_9; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_10; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_11; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_12; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_13; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_14; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_16; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_17; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_18; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_19; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_20; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_21; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_22; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_23; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_24; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_25; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_26; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_27; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_28; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_29; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_30; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_31; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_32; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_33; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_34; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_35; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_36; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_37; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_38; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_39; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_40; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_41; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_42; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_43; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_44; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_45; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_46; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_47; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_48; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_49; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_50; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_51; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_52; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_53; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_54; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_55; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_56; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_57; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_58; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_59; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_60; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_61; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_62; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_63; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_64; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_65; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_66; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_67; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_68; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_69; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_70; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_71; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_72; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_73; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_74; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_75; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_76; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_77; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_78; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_79; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_80; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_81; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_82; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_83; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_84; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_85; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_86; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_87; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_88; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_89; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_90; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_91; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_92; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_93; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_94; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_95; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_96; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_97; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_98; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_99; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_100; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_101; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_102; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_103; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_104; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_105; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_106; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_107; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_108; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_109; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_110; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_111; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_112; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_113; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_114; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_115; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_116; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_117; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_118; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_119; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_120; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_121; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_122; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_123; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_124; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_125; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_126; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_127; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_128; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_129; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_130; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_131; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_132; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_133; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_134; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_135; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_136; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_137; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_138; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_139; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_140; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_141; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_142; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_143; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_144; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_145; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_146; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_147; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_148; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_149; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_150; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_151; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_152; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_153; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_154; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_155; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_156; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_157; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_158; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_data_159; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_0; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_1; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_2; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_3; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_4; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_5; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_6; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_7; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_8; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_9; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_10; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_11; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_12; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_13; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_14; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_header_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_state; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_in_parse_current_offset; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_in_parse_transition_field; // @[matcher.scala 349:24]
  wire [3:0] pipe12_io_pipe_phv_in_next_processor_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_next_config_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_is_valid_processor; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_valid; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_in_last; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_96; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_97; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_98; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_99; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_100; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_101; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_102; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_103; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_104; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_105; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_106; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_107; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_108; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_109; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_110; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_111; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_112; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_113; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_114; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_115; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_116; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_117; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_118; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_119; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_120; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_121; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_122; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_123; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_124; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_125; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_126; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_127; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_128; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_129; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_130; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_131; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_132; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_133; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_134; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_135; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_136; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_137; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_138; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_139; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_140; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_141; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_142; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_143; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_144; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_145; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_146; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_147; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_148; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_149; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_150; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_151; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_152; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_153; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_154; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_155; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_156; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_157; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_158; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_data_159; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 349:24]
  wire [7:0] pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 349:24]
  wire [15:0] pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 349:24]
  wire [3:0] pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_valid; // @[matcher.scala 349:24]
  wire  pipe12_io_pipe_phv_out_last; // @[matcher.scala 349:24]
  MatchGetOffset pipe1 ( // @[matcher.scala 343:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(pipe1_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(pipe1_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(pipe1_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(pipe1_io_pipe_phv_out_last)
  );
  MatchGetKey pipe2 ( // @[matcher.scala 344:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(pipe2_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(pipe2_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(pipe2_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(pipe2_io_pipe_phv_out_last)
  );
  Hash pipe3to8 ( // @[matcher.scala 345:26]
    .clock(pipe3to8_clock),
    .io_pipe_phv_in_data_0(pipe3to8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3to8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3to8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3to8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3to8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3to8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3to8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3to8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3to8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3to8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3to8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3to8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3to8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3to8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3to8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3to8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3to8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3to8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3to8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3to8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3to8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3to8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3to8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3to8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3to8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3to8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3to8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3to8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3to8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3to8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3to8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3to8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3to8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3to8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3to8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3to8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3to8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3to8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3to8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3to8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3to8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3to8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3to8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3to8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3to8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3to8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3to8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3to8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3to8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3to8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3to8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3to8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3to8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3to8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3to8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3to8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3to8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3to8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3to8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3to8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3to8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3to8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3to8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3to8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3to8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3to8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3to8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3to8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3to8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3to8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3to8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3to8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3to8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3to8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3to8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3to8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3to8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3to8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3to8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3to8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3to8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3to8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3to8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3to8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3to8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3to8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3to8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3to8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3to8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3to8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3to8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3to8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3to8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3to8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3to8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3to8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3to8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3to8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3to8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3to8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3to8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3to8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3to8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3to8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3to8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3to8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3to8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3to8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3to8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3to8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3to8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3to8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3to8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3to8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3to8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3to8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3to8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3to8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3to8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3to8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3to8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3to8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3to8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3to8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3to8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3to8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3to8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3to8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3to8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3to8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3to8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3to8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3to8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3to8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3to8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3to8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3to8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3to8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3to8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3to8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3to8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3to8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3to8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3to8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3to8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3to8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3to8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3to8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3to8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3to8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3to8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3to8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3to8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3to8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3to8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3to8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3to8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3to8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3to8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3to8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe3to8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3to8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3to8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3to8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3to8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3to8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3to8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3to8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3to8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3to8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3to8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3to8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3to8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3to8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3to8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3to8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3to8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3to8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3to8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3to8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3to8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3to8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(pipe3to8_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(pipe3to8_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(pipe3to8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3to8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3to8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3to8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3to8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3to8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3to8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3to8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3to8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3to8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3to8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3to8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3to8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3to8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3to8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3to8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3to8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3to8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3to8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3to8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3to8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3to8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3to8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3to8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3to8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3to8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3to8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3to8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3to8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3to8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3to8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3to8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3to8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3to8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3to8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3to8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3to8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3to8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3to8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3to8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3to8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3to8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3to8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3to8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3to8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3to8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3to8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3to8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3to8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3to8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3to8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3to8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3to8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3to8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3to8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3to8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3to8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3to8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3to8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3to8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3to8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3to8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3to8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3to8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3to8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3to8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3to8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3to8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3to8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3to8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3to8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3to8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3to8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3to8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3to8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3to8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3to8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3to8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3to8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3to8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3to8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3to8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3to8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3to8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3to8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3to8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3to8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3to8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3to8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3to8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3to8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3to8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3to8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3to8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3to8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3to8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3to8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3to8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3to8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3to8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3to8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3to8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3to8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3to8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3to8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3to8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3to8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3to8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3to8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3to8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3to8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3to8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3to8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3to8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3to8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3to8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3to8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3to8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3to8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3to8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3to8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3to8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3to8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3to8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3to8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3to8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3to8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3to8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3to8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3to8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3to8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3to8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3to8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3to8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3to8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3to8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3to8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3to8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3to8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3to8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3to8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3to8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3to8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3to8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3to8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3to8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3to8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3to8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3to8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3to8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3to8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3to8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3to8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3to8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3to8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3to8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3to8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3to8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3to8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3to8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe3to8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3to8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3to8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3to8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3to8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3to8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3to8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3to8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3to8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3to8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3to8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3to8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3to8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3to8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3to8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3to8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3to8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3to8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3to8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3to8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3to8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3to8_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(pipe3to8_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(pipe3to8_io_pipe_phv_out_last)
  );
  MatchGetCs pipe9 ( // @[matcher.scala 346:23]
    .clock(pipe9_clock),
    .io_pipe_phv_in_data_0(pipe9_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe9_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe9_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe9_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe9_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe9_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe9_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe9_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe9_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe9_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe9_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe9_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe9_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe9_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe9_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe9_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe9_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe9_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe9_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe9_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe9_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe9_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe9_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe9_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe9_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe9_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe9_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe9_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe9_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe9_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe9_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe9_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe9_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe9_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe9_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe9_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe9_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe9_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe9_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe9_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe9_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe9_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe9_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe9_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe9_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe9_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe9_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe9_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe9_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe9_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe9_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe9_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe9_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe9_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe9_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe9_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe9_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe9_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe9_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe9_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe9_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe9_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe9_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe9_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe9_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe9_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe9_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe9_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe9_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe9_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe9_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe9_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe9_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe9_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe9_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe9_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe9_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe9_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe9_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe9_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe9_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe9_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe9_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe9_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe9_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe9_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe9_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe9_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe9_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe9_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe9_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe9_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe9_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe9_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe9_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe9_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe9_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe9_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe9_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe9_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe9_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe9_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe9_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe9_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe9_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe9_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe9_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe9_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe9_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe9_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe9_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe9_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe9_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe9_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe9_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe9_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe9_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe9_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe9_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe9_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe9_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe9_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe9_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe9_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe9_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe9_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe9_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe9_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe9_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe9_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe9_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe9_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe9_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe9_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe9_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe9_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe9_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe9_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe9_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe9_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe9_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe9_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe9_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe9_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe9_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe9_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe9_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe9_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe9_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe9_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe9_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe9_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe9_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe9_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe9_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe9_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe9_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe9_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe9_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe9_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe9_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe9_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe9_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe9_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe9_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe9_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe9_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe9_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe9_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe9_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe9_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe9_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe9_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe9_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe9_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe9_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe9_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe9_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe9_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe9_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe9_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe9_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(pipe9_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(pipe9_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(pipe9_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe9_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe9_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe9_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe9_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe9_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe9_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe9_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe9_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe9_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe9_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe9_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe9_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe9_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe9_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe9_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe9_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe9_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe9_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe9_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe9_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe9_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe9_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe9_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe9_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe9_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe9_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe9_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe9_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe9_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe9_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe9_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe9_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe9_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe9_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe9_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe9_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe9_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe9_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe9_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe9_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe9_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe9_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe9_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe9_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe9_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe9_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe9_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe9_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe9_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe9_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe9_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe9_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe9_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe9_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe9_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe9_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe9_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe9_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe9_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe9_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe9_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe9_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe9_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe9_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe9_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe9_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe9_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe9_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe9_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe9_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe9_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe9_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe9_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe9_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe9_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe9_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe9_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe9_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe9_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe9_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe9_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe9_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe9_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe9_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe9_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe9_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe9_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe9_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe9_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe9_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe9_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe9_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe9_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe9_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe9_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe9_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe9_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe9_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe9_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe9_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe9_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe9_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe9_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe9_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe9_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe9_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe9_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe9_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe9_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe9_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe9_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe9_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe9_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe9_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe9_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe9_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe9_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe9_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe9_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe9_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe9_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe9_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe9_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe9_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe9_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe9_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe9_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe9_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe9_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe9_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe9_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe9_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe9_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe9_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe9_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe9_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe9_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe9_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe9_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe9_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe9_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe9_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe9_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe9_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe9_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe9_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe9_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe9_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe9_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe9_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe9_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe9_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe9_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe9_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe9_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe9_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe9_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe9_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe9_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe9_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe9_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe9_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe9_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe9_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe9_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe9_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe9_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe9_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe9_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe9_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe9_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe9_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe9_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe9_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe9_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe9_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe9_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe9_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe9_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe9_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe9_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(pipe9_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(pipe9_io_pipe_phv_out_last)
  );
  MatchReadData pipe10 ( // @[matcher.scala 347:24]
    .clock(pipe10_clock),
    .io_pipe_phv_in_data_0(pipe10_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe10_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe10_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe10_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe10_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe10_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe10_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe10_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe10_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe10_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe10_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe10_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe10_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe10_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe10_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe10_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe10_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe10_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe10_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe10_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe10_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe10_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe10_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe10_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe10_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe10_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe10_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe10_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe10_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe10_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe10_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe10_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe10_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe10_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe10_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe10_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe10_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe10_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe10_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe10_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe10_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe10_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe10_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe10_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe10_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe10_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe10_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe10_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe10_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe10_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe10_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe10_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe10_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe10_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe10_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe10_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe10_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe10_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe10_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe10_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe10_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe10_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe10_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe10_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe10_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe10_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe10_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe10_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe10_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe10_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe10_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe10_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe10_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe10_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe10_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe10_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe10_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe10_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe10_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe10_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe10_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe10_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe10_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe10_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe10_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe10_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe10_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe10_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe10_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe10_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe10_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe10_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe10_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe10_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe10_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe10_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe10_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe10_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe10_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe10_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe10_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe10_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe10_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe10_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe10_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe10_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe10_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe10_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe10_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe10_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe10_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe10_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe10_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe10_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe10_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe10_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe10_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe10_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe10_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe10_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe10_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe10_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe10_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe10_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe10_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe10_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe10_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe10_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe10_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe10_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe10_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe10_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe10_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe10_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe10_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe10_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe10_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe10_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe10_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe10_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe10_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe10_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe10_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe10_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe10_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe10_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe10_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe10_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe10_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe10_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe10_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe10_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe10_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe10_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe10_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe10_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe10_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe10_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe10_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe10_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe10_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe10_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe10_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe10_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe10_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe10_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe10_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe10_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe10_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe10_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe10_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe10_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe10_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe10_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe10_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe10_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe10_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe10_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe10_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe10_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe10_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe10_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(pipe10_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(pipe10_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(pipe10_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe10_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe10_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe10_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe10_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe10_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe10_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe10_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe10_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe10_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe10_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe10_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe10_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe10_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe10_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe10_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe10_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe10_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe10_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe10_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe10_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe10_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe10_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe10_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe10_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe10_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe10_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe10_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe10_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe10_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe10_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe10_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe10_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe10_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe10_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe10_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe10_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe10_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe10_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe10_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe10_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe10_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe10_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe10_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe10_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe10_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe10_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe10_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe10_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe10_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe10_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe10_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe10_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe10_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe10_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe10_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe10_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe10_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe10_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe10_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe10_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe10_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe10_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe10_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe10_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe10_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe10_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe10_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe10_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe10_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe10_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe10_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe10_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe10_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe10_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe10_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe10_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe10_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe10_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe10_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe10_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe10_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe10_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe10_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe10_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe10_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe10_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe10_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe10_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe10_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe10_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe10_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe10_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe10_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe10_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe10_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe10_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe10_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe10_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe10_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe10_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe10_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe10_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe10_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe10_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe10_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe10_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe10_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe10_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe10_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe10_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe10_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe10_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe10_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe10_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe10_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe10_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe10_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe10_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe10_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe10_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe10_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe10_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe10_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe10_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe10_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe10_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe10_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe10_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe10_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe10_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe10_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe10_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe10_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe10_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe10_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe10_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe10_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe10_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe10_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe10_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe10_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe10_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe10_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe10_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe10_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe10_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe10_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe10_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe10_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe10_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe10_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe10_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe10_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe10_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe10_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe10_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe10_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe10_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe10_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe10_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe10_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe10_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe10_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe10_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe10_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe10_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe10_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe10_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe10_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe10_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe10_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe10_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe10_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe10_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe10_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe10_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe10_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe10_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe10_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe10_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe10_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(pipe10_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(pipe10_io_pipe_phv_out_last)
  );
  MatchDataReshape pipe11 ( // @[matcher.scala 348:24]
    .clock(pipe11_clock),
    .io_pipe_phv_in_data_0(pipe11_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe11_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe11_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe11_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe11_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe11_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe11_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe11_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe11_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe11_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe11_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe11_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe11_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe11_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe11_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe11_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe11_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe11_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe11_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe11_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe11_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe11_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe11_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe11_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe11_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe11_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe11_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe11_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe11_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe11_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe11_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe11_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe11_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe11_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe11_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe11_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe11_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe11_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe11_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe11_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe11_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe11_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe11_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe11_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe11_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe11_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe11_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe11_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe11_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe11_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe11_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe11_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe11_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe11_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe11_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe11_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe11_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe11_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe11_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe11_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe11_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe11_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe11_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe11_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe11_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe11_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe11_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe11_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe11_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe11_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe11_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe11_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe11_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe11_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe11_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe11_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe11_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe11_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe11_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe11_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe11_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe11_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe11_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe11_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe11_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe11_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe11_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe11_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe11_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe11_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe11_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe11_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe11_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe11_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe11_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe11_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe11_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe11_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe11_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe11_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe11_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe11_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe11_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe11_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe11_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe11_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe11_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe11_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe11_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe11_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe11_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe11_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe11_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe11_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe11_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe11_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe11_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe11_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe11_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe11_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe11_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe11_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe11_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe11_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe11_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe11_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe11_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe11_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe11_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe11_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe11_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe11_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe11_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe11_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe11_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe11_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe11_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe11_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe11_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe11_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe11_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe11_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe11_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe11_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe11_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe11_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe11_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe11_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe11_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe11_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe11_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe11_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe11_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe11_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe11_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe11_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe11_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe11_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe11_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe11_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe11_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe11_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe11_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe11_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe11_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe11_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe11_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe11_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe11_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe11_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe11_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe11_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe11_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe11_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe11_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe11_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe11_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe11_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe11_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe11_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe11_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe11_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(pipe11_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(pipe11_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(pipe11_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe11_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe11_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe11_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe11_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe11_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe11_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe11_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe11_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe11_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe11_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe11_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe11_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe11_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe11_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe11_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe11_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe11_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe11_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe11_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe11_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe11_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe11_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe11_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe11_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe11_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe11_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe11_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe11_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe11_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe11_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe11_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe11_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe11_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe11_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe11_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe11_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe11_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe11_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe11_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe11_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe11_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe11_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe11_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe11_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe11_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe11_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe11_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe11_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe11_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe11_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe11_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe11_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe11_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe11_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe11_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe11_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe11_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe11_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe11_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe11_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe11_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe11_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe11_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe11_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe11_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe11_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe11_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe11_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe11_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe11_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe11_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe11_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe11_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe11_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe11_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe11_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe11_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe11_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe11_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe11_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe11_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe11_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe11_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe11_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe11_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe11_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe11_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe11_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe11_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe11_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe11_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe11_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe11_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe11_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe11_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe11_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe11_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe11_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe11_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe11_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe11_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe11_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe11_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe11_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe11_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe11_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe11_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe11_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe11_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe11_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe11_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe11_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe11_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe11_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe11_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe11_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe11_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe11_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe11_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe11_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe11_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe11_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe11_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe11_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe11_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe11_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe11_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe11_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe11_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe11_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe11_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe11_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe11_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe11_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe11_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe11_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe11_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe11_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe11_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe11_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe11_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe11_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe11_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe11_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe11_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe11_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe11_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe11_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe11_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe11_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe11_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe11_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe11_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe11_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe11_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe11_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe11_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe11_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe11_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe11_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe11_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe11_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe11_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe11_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe11_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe11_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe11_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe11_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe11_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe11_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe11_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe11_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe11_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe11_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe11_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe11_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe11_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe11_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe11_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe11_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe11_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(pipe11_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(pipe11_io_pipe_phv_out_last)
  );
  MatchResult pipe12 ( // @[matcher.scala 349:24]
    .clock(pipe12_clock),
    .io_pipe_phv_in_data_0(pipe12_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe12_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe12_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe12_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe12_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe12_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe12_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe12_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe12_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe12_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe12_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe12_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe12_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe12_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe12_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe12_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe12_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe12_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe12_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe12_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe12_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe12_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe12_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe12_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe12_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe12_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe12_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe12_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe12_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe12_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe12_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe12_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe12_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe12_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe12_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe12_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe12_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe12_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe12_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe12_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe12_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe12_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe12_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe12_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe12_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe12_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe12_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe12_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe12_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe12_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe12_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe12_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe12_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe12_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe12_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe12_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe12_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe12_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe12_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe12_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe12_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe12_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe12_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe12_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe12_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe12_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe12_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe12_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe12_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe12_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe12_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe12_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe12_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe12_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe12_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe12_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe12_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe12_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe12_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe12_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe12_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe12_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe12_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe12_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe12_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe12_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe12_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe12_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe12_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe12_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe12_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe12_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe12_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe12_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe12_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe12_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe12_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe12_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe12_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe12_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe12_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe12_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe12_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe12_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe12_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe12_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe12_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe12_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe12_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe12_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe12_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe12_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe12_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe12_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe12_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe12_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe12_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe12_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe12_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe12_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe12_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe12_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe12_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe12_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe12_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe12_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe12_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe12_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe12_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe12_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe12_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe12_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe12_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe12_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe12_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe12_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe12_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe12_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe12_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe12_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe12_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe12_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe12_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe12_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe12_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe12_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe12_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe12_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe12_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe12_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe12_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe12_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe12_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe12_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe12_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe12_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe12_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe12_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe12_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe12_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe12_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe12_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe12_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe12_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe12_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe12_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe12_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe12_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe12_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe12_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe12_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe12_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe12_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe12_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe12_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe12_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe12_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe12_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe12_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe12_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe12_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe12_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(pipe12_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(pipe12_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(pipe12_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe12_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe12_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe12_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe12_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe12_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe12_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe12_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe12_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe12_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe12_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe12_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe12_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe12_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe12_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe12_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe12_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe12_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe12_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe12_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe12_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe12_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe12_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe12_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe12_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe12_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe12_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe12_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe12_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe12_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe12_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe12_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe12_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe12_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe12_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe12_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe12_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe12_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe12_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe12_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe12_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe12_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe12_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe12_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe12_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe12_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe12_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe12_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe12_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe12_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe12_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe12_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe12_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe12_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe12_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe12_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe12_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe12_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe12_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe12_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe12_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe12_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe12_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe12_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe12_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe12_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe12_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe12_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe12_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe12_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe12_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe12_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe12_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe12_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe12_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe12_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe12_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe12_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe12_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe12_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe12_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe12_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe12_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe12_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe12_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe12_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe12_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe12_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe12_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe12_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe12_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe12_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe12_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe12_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe12_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe12_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe12_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe12_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe12_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe12_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe12_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe12_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe12_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe12_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe12_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe12_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe12_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe12_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe12_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe12_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe12_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe12_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe12_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe12_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe12_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe12_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe12_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe12_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe12_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe12_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe12_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe12_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe12_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe12_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe12_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe12_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe12_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe12_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe12_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe12_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe12_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe12_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe12_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe12_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe12_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe12_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe12_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe12_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe12_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe12_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe12_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe12_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe12_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe12_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe12_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe12_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe12_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe12_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe12_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe12_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe12_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe12_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe12_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe12_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe12_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe12_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe12_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe12_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe12_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe12_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe12_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe12_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe12_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe12_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe12_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe12_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe12_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe12_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe12_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe12_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe12_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe12_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe12_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe12_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe12_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe12_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe12_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe12_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe12_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe12_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe12_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe12_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(pipe12_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(pipe12_io_pipe_phv_out_last)
  );
  assign io_pipe_phv_out_data_0 = pipe12_io_pipe_phv_out_data_0; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_1 = pipe12_io_pipe_phv_out_data_1; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_2 = pipe12_io_pipe_phv_out_data_2; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_3 = pipe12_io_pipe_phv_out_data_3; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_4 = pipe12_io_pipe_phv_out_data_4; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_5 = pipe12_io_pipe_phv_out_data_5; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_6 = pipe12_io_pipe_phv_out_data_6; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_7 = pipe12_io_pipe_phv_out_data_7; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_8 = pipe12_io_pipe_phv_out_data_8; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_9 = pipe12_io_pipe_phv_out_data_9; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_10 = pipe12_io_pipe_phv_out_data_10; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_11 = pipe12_io_pipe_phv_out_data_11; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_12 = pipe12_io_pipe_phv_out_data_12; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_13 = pipe12_io_pipe_phv_out_data_13; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_14 = pipe12_io_pipe_phv_out_data_14; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_15 = pipe12_io_pipe_phv_out_data_15; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_16 = pipe12_io_pipe_phv_out_data_16; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_17 = pipe12_io_pipe_phv_out_data_17; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_18 = pipe12_io_pipe_phv_out_data_18; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_19 = pipe12_io_pipe_phv_out_data_19; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_20 = pipe12_io_pipe_phv_out_data_20; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_21 = pipe12_io_pipe_phv_out_data_21; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_22 = pipe12_io_pipe_phv_out_data_22; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_23 = pipe12_io_pipe_phv_out_data_23; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_24 = pipe12_io_pipe_phv_out_data_24; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_25 = pipe12_io_pipe_phv_out_data_25; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_26 = pipe12_io_pipe_phv_out_data_26; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_27 = pipe12_io_pipe_phv_out_data_27; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_28 = pipe12_io_pipe_phv_out_data_28; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_29 = pipe12_io_pipe_phv_out_data_29; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_30 = pipe12_io_pipe_phv_out_data_30; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_31 = pipe12_io_pipe_phv_out_data_31; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_32 = pipe12_io_pipe_phv_out_data_32; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_33 = pipe12_io_pipe_phv_out_data_33; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_34 = pipe12_io_pipe_phv_out_data_34; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_35 = pipe12_io_pipe_phv_out_data_35; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_36 = pipe12_io_pipe_phv_out_data_36; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_37 = pipe12_io_pipe_phv_out_data_37; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_38 = pipe12_io_pipe_phv_out_data_38; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_39 = pipe12_io_pipe_phv_out_data_39; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_40 = pipe12_io_pipe_phv_out_data_40; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_41 = pipe12_io_pipe_phv_out_data_41; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_42 = pipe12_io_pipe_phv_out_data_42; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_43 = pipe12_io_pipe_phv_out_data_43; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_44 = pipe12_io_pipe_phv_out_data_44; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_45 = pipe12_io_pipe_phv_out_data_45; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_46 = pipe12_io_pipe_phv_out_data_46; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_47 = pipe12_io_pipe_phv_out_data_47; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_48 = pipe12_io_pipe_phv_out_data_48; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_49 = pipe12_io_pipe_phv_out_data_49; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_50 = pipe12_io_pipe_phv_out_data_50; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_51 = pipe12_io_pipe_phv_out_data_51; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_52 = pipe12_io_pipe_phv_out_data_52; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_53 = pipe12_io_pipe_phv_out_data_53; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_54 = pipe12_io_pipe_phv_out_data_54; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_55 = pipe12_io_pipe_phv_out_data_55; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_56 = pipe12_io_pipe_phv_out_data_56; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_57 = pipe12_io_pipe_phv_out_data_57; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_58 = pipe12_io_pipe_phv_out_data_58; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_59 = pipe12_io_pipe_phv_out_data_59; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_60 = pipe12_io_pipe_phv_out_data_60; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_61 = pipe12_io_pipe_phv_out_data_61; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_62 = pipe12_io_pipe_phv_out_data_62; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_63 = pipe12_io_pipe_phv_out_data_63; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_64 = pipe12_io_pipe_phv_out_data_64; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_65 = pipe12_io_pipe_phv_out_data_65; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_66 = pipe12_io_pipe_phv_out_data_66; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_67 = pipe12_io_pipe_phv_out_data_67; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_68 = pipe12_io_pipe_phv_out_data_68; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_69 = pipe12_io_pipe_phv_out_data_69; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_70 = pipe12_io_pipe_phv_out_data_70; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_71 = pipe12_io_pipe_phv_out_data_71; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_72 = pipe12_io_pipe_phv_out_data_72; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_73 = pipe12_io_pipe_phv_out_data_73; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_74 = pipe12_io_pipe_phv_out_data_74; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_75 = pipe12_io_pipe_phv_out_data_75; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_76 = pipe12_io_pipe_phv_out_data_76; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_77 = pipe12_io_pipe_phv_out_data_77; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_78 = pipe12_io_pipe_phv_out_data_78; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_79 = pipe12_io_pipe_phv_out_data_79; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_80 = pipe12_io_pipe_phv_out_data_80; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_81 = pipe12_io_pipe_phv_out_data_81; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_82 = pipe12_io_pipe_phv_out_data_82; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_83 = pipe12_io_pipe_phv_out_data_83; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_84 = pipe12_io_pipe_phv_out_data_84; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_85 = pipe12_io_pipe_phv_out_data_85; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_86 = pipe12_io_pipe_phv_out_data_86; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_87 = pipe12_io_pipe_phv_out_data_87; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_88 = pipe12_io_pipe_phv_out_data_88; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_89 = pipe12_io_pipe_phv_out_data_89; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_90 = pipe12_io_pipe_phv_out_data_90; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_91 = pipe12_io_pipe_phv_out_data_91; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_92 = pipe12_io_pipe_phv_out_data_92; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_93 = pipe12_io_pipe_phv_out_data_93; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_94 = pipe12_io_pipe_phv_out_data_94; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_95 = pipe12_io_pipe_phv_out_data_95; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_96 = pipe12_io_pipe_phv_out_data_96; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_97 = pipe12_io_pipe_phv_out_data_97; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_98 = pipe12_io_pipe_phv_out_data_98; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_99 = pipe12_io_pipe_phv_out_data_99; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_100 = pipe12_io_pipe_phv_out_data_100; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_101 = pipe12_io_pipe_phv_out_data_101; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_102 = pipe12_io_pipe_phv_out_data_102; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_103 = pipe12_io_pipe_phv_out_data_103; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_104 = pipe12_io_pipe_phv_out_data_104; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_105 = pipe12_io_pipe_phv_out_data_105; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_106 = pipe12_io_pipe_phv_out_data_106; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_107 = pipe12_io_pipe_phv_out_data_107; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_108 = pipe12_io_pipe_phv_out_data_108; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_109 = pipe12_io_pipe_phv_out_data_109; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_110 = pipe12_io_pipe_phv_out_data_110; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_111 = pipe12_io_pipe_phv_out_data_111; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_112 = pipe12_io_pipe_phv_out_data_112; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_113 = pipe12_io_pipe_phv_out_data_113; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_114 = pipe12_io_pipe_phv_out_data_114; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_115 = pipe12_io_pipe_phv_out_data_115; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_116 = pipe12_io_pipe_phv_out_data_116; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_117 = pipe12_io_pipe_phv_out_data_117; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_118 = pipe12_io_pipe_phv_out_data_118; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_119 = pipe12_io_pipe_phv_out_data_119; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_120 = pipe12_io_pipe_phv_out_data_120; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_121 = pipe12_io_pipe_phv_out_data_121; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_122 = pipe12_io_pipe_phv_out_data_122; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_123 = pipe12_io_pipe_phv_out_data_123; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_124 = pipe12_io_pipe_phv_out_data_124; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_125 = pipe12_io_pipe_phv_out_data_125; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_126 = pipe12_io_pipe_phv_out_data_126; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_127 = pipe12_io_pipe_phv_out_data_127; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_128 = pipe12_io_pipe_phv_out_data_128; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_129 = pipe12_io_pipe_phv_out_data_129; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_130 = pipe12_io_pipe_phv_out_data_130; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_131 = pipe12_io_pipe_phv_out_data_131; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_132 = pipe12_io_pipe_phv_out_data_132; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_133 = pipe12_io_pipe_phv_out_data_133; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_134 = pipe12_io_pipe_phv_out_data_134; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_135 = pipe12_io_pipe_phv_out_data_135; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_136 = pipe12_io_pipe_phv_out_data_136; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_137 = pipe12_io_pipe_phv_out_data_137; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_138 = pipe12_io_pipe_phv_out_data_138; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_139 = pipe12_io_pipe_phv_out_data_139; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_140 = pipe12_io_pipe_phv_out_data_140; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_141 = pipe12_io_pipe_phv_out_data_141; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_142 = pipe12_io_pipe_phv_out_data_142; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_143 = pipe12_io_pipe_phv_out_data_143; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_144 = pipe12_io_pipe_phv_out_data_144; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_145 = pipe12_io_pipe_phv_out_data_145; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_146 = pipe12_io_pipe_phv_out_data_146; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_147 = pipe12_io_pipe_phv_out_data_147; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_148 = pipe12_io_pipe_phv_out_data_148; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_149 = pipe12_io_pipe_phv_out_data_149; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_150 = pipe12_io_pipe_phv_out_data_150; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_151 = pipe12_io_pipe_phv_out_data_151; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_152 = pipe12_io_pipe_phv_out_data_152; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_153 = pipe12_io_pipe_phv_out_data_153; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_154 = pipe12_io_pipe_phv_out_data_154; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_155 = pipe12_io_pipe_phv_out_data_155; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_156 = pipe12_io_pipe_phv_out_data_156; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_157 = pipe12_io_pipe_phv_out_data_157; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_158 = pipe12_io_pipe_phv_out_data_158; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_data_159 = pipe12_io_pipe_phv_out_data_159; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_0 = pipe12_io_pipe_phv_out_header_0; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_1 = pipe12_io_pipe_phv_out_header_1; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_2 = pipe12_io_pipe_phv_out_header_2; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_3 = pipe12_io_pipe_phv_out_header_3; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_4 = pipe12_io_pipe_phv_out_header_4; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_5 = pipe12_io_pipe_phv_out_header_5; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_6 = pipe12_io_pipe_phv_out_header_6; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_7 = pipe12_io_pipe_phv_out_header_7; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_8 = pipe12_io_pipe_phv_out_header_8; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_9 = pipe12_io_pipe_phv_out_header_9; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_10 = pipe12_io_pipe_phv_out_header_10; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_11 = pipe12_io_pipe_phv_out_header_11; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_12 = pipe12_io_pipe_phv_out_header_12; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_13 = pipe12_io_pipe_phv_out_header_13; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_14 = pipe12_io_pipe_phv_out_header_14; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_header_15 = pipe12_io_pipe_phv_out_header_15; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_current_state = pipe12_io_pipe_phv_out_parse_current_state; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_current_offset = pipe12_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_parse_transition_field = pipe12_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_next_processor_id = pipe12_io_pipe_phv_out_next_processor_id; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_next_config_id = pipe12_io_pipe_phv_out_next_config_id; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_is_valid_processor = pipe12_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_valid = pipe12_io_pipe_phv_out_valid; // @[matcher.scala 388:27]
  assign io_pipe_phv_out_last = pipe12_io_pipe_phv_out_last; // @[matcher.scala 388:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_valid = io_pipe_phv_in_valid; // @[matcher.scala 351:26]
  assign pipe1_io_pipe_phv_in_last = io_pipe_phv_in_last; // @[matcher.scala 351:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_valid = pipe1_io_pipe_phv_out_valid; // @[matcher.scala 354:26]
  assign pipe2_io_pipe_phv_in_last = pipe1_io_pipe_phv_out_last; // @[matcher.scala 354:26]
  assign pipe3to8_clock = clock;
  assign pipe3to8_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_valid = pipe2_io_pipe_phv_out_valid; // @[matcher.scala 358:29]
  assign pipe3to8_io_pipe_phv_in_last = pipe2_io_pipe_phv_out_last; // @[matcher.scala 358:29]
  assign pipe9_clock = clock;
  assign pipe9_io_pipe_phv_in_data_0 = pipe3to8_io_pipe_phv_out_data_0; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_1 = pipe3to8_io_pipe_phv_out_data_1; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_2 = pipe3to8_io_pipe_phv_out_data_2; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_3 = pipe3to8_io_pipe_phv_out_data_3; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_4 = pipe3to8_io_pipe_phv_out_data_4; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_5 = pipe3to8_io_pipe_phv_out_data_5; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_6 = pipe3to8_io_pipe_phv_out_data_6; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_7 = pipe3to8_io_pipe_phv_out_data_7; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_8 = pipe3to8_io_pipe_phv_out_data_8; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_9 = pipe3to8_io_pipe_phv_out_data_9; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_10 = pipe3to8_io_pipe_phv_out_data_10; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_11 = pipe3to8_io_pipe_phv_out_data_11; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_12 = pipe3to8_io_pipe_phv_out_data_12; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_13 = pipe3to8_io_pipe_phv_out_data_13; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_14 = pipe3to8_io_pipe_phv_out_data_14; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_15 = pipe3to8_io_pipe_phv_out_data_15; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_16 = pipe3to8_io_pipe_phv_out_data_16; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_17 = pipe3to8_io_pipe_phv_out_data_17; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_18 = pipe3to8_io_pipe_phv_out_data_18; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_19 = pipe3to8_io_pipe_phv_out_data_19; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_20 = pipe3to8_io_pipe_phv_out_data_20; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_21 = pipe3to8_io_pipe_phv_out_data_21; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_22 = pipe3to8_io_pipe_phv_out_data_22; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_23 = pipe3to8_io_pipe_phv_out_data_23; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_24 = pipe3to8_io_pipe_phv_out_data_24; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_25 = pipe3to8_io_pipe_phv_out_data_25; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_26 = pipe3to8_io_pipe_phv_out_data_26; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_27 = pipe3to8_io_pipe_phv_out_data_27; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_28 = pipe3to8_io_pipe_phv_out_data_28; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_29 = pipe3to8_io_pipe_phv_out_data_29; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_30 = pipe3to8_io_pipe_phv_out_data_30; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_31 = pipe3to8_io_pipe_phv_out_data_31; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_32 = pipe3to8_io_pipe_phv_out_data_32; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_33 = pipe3to8_io_pipe_phv_out_data_33; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_34 = pipe3to8_io_pipe_phv_out_data_34; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_35 = pipe3to8_io_pipe_phv_out_data_35; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_36 = pipe3to8_io_pipe_phv_out_data_36; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_37 = pipe3to8_io_pipe_phv_out_data_37; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_38 = pipe3to8_io_pipe_phv_out_data_38; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_39 = pipe3to8_io_pipe_phv_out_data_39; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_40 = pipe3to8_io_pipe_phv_out_data_40; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_41 = pipe3to8_io_pipe_phv_out_data_41; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_42 = pipe3to8_io_pipe_phv_out_data_42; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_43 = pipe3to8_io_pipe_phv_out_data_43; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_44 = pipe3to8_io_pipe_phv_out_data_44; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_45 = pipe3to8_io_pipe_phv_out_data_45; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_46 = pipe3to8_io_pipe_phv_out_data_46; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_47 = pipe3to8_io_pipe_phv_out_data_47; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_48 = pipe3to8_io_pipe_phv_out_data_48; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_49 = pipe3to8_io_pipe_phv_out_data_49; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_50 = pipe3to8_io_pipe_phv_out_data_50; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_51 = pipe3to8_io_pipe_phv_out_data_51; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_52 = pipe3to8_io_pipe_phv_out_data_52; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_53 = pipe3to8_io_pipe_phv_out_data_53; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_54 = pipe3to8_io_pipe_phv_out_data_54; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_55 = pipe3to8_io_pipe_phv_out_data_55; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_56 = pipe3to8_io_pipe_phv_out_data_56; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_57 = pipe3to8_io_pipe_phv_out_data_57; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_58 = pipe3to8_io_pipe_phv_out_data_58; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_59 = pipe3to8_io_pipe_phv_out_data_59; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_60 = pipe3to8_io_pipe_phv_out_data_60; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_61 = pipe3to8_io_pipe_phv_out_data_61; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_62 = pipe3to8_io_pipe_phv_out_data_62; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_63 = pipe3to8_io_pipe_phv_out_data_63; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_64 = pipe3to8_io_pipe_phv_out_data_64; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_65 = pipe3to8_io_pipe_phv_out_data_65; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_66 = pipe3to8_io_pipe_phv_out_data_66; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_67 = pipe3to8_io_pipe_phv_out_data_67; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_68 = pipe3to8_io_pipe_phv_out_data_68; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_69 = pipe3to8_io_pipe_phv_out_data_69; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_70 = pipe3to8_io_pipe_phv_out_data_70; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_71 = pipe3to8_io_pipe_phv_out_data_71; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_72 = pipe3to8_io_pipe_phv_out_data_72; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_73 = pipe3to8_io_pipe_phv_out_data_73; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_74 = pipe3to8_io_pipe_phv_out_data_74; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_75 = pipe3to8_io_pipe_phv_out_data_75; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_76 = pipe3to8_io_pipe_phv_out_data_76; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_77 = pipe3to8_io_pipe_phv_out_data_77; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_78 = pipe3to8_io_pipe_phv_out_data_78; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_79 = pipe3to8_io_pipe_phv_out_data_79; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_80 = pipe3to8_io_pipe_phv_out_data_80; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_81 = pipe3to8_io_pipe_phv_out_data_81; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_82 = pipe3to8_io_pipe_phv_out_data_82; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_83 = pipe3to8_io_pipe_phv_out_data_83; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_84 = pipe3to8_io_pipe_phv_out_data_84; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_85 = pipe3to8_io_pipe_phv_out_data_85; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_86 = pipe3to8_io_pipe_phv_out_data_86; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_87 = pipe3to8_io_pipe_phv_out_data_87; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_88 = pipe3to8_io_pipe_phv_out_data_88; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_89 = pipe3to8_io_pipe_phv_out_data_89; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_90 = pipe3to8_io_pipe_phv_out_data_90; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_91 = pipe3to8_io_pipe_phv_out_data_91; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_92 = pipe3to8_io_pipe_phv_out_data_92; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_93 = pipe3to8_io_pipe_phv_out_data_93; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_94 = pipe3to8_io_pipe_phv_out_data_94; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_95 = pipe3to8_io_pipe_phv_out_data_95; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_96 = pipe3to8_io_pipe_phv_out_data_96; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_97 = pipe3to8_io_pipe_phv_out_data_97; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_98 = pipe3to8_io_pipe_phv_out_data_98; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_99 = pipe3to8_io_pipe_phv_out_data_99; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_100 = pipe3to8_io_pipe_phv_out_data_100; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_101 = pipe3to8_io_pipe_phv_out_data_101; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_102 = pipe3to8_io_pipe_phv_out_data_102; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_103 = pipe3to8_io_pipe_phv_out_data_103; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_104 = pipe3to8_io_pipe_phv_out_data_104; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_105 = pipe3to8_io_pipe_phv_out_data_105; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_106 = pipe3to8_io_pipe_phv_out_data_106; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_107 = pipe3to8_io_pipe_phv_out_data_107; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_108 = pipe3to8_io_pipe_phv_out_data_108; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_109 = pipe3to8_io_pipe_phv_out_data_109; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_110 = pipe3to8_io_pipe_phv_out_data_110; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_111 = pipe3to8_io_pipe_phv_out_data_111; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_112 = pipe3to8_io_pipe_phv_out_data_112; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_113 = pipe3to8_io_pipe_phv_out_data_113; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_114 = pipe3to8_io_pipe_phv_out_data_114; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_115 = pipe3to8_io_pipe_phv_out_data_115; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_116 = pipe3to8_io_pipe_phv_out_data_116; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_117 = pipe3to8_io_pipe_phv_out_data_117; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_118 = pipe3to8_io_pipe_phv_out_data_118; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_119 = pipe3to8_io_pipe_phv_out_data_119; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_120 = pipe3to8_io_pipe_phv_out_data_120; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_121 = pipe3to8_io_pipe_phv_out_data_121; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_122 = pipe3to8_io_pipe_phv_out_data_122; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_123 = pipe3to8_io_pipe_phv_out_data_123; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_124 = pipe3to8_io_pipe_phv_out_data_124; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_125 = pipe3to8_io_pipe_phv_out_data_125; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_126 = pipe3to8_io_pipe_phv_out_data_126; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_127 = pipe3to8_io_pipe_phv_out_data_127; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_128 = pipe3to8_io_pipe_phv_out_data_128; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_129 = pipe3to8_io_pipe_phv_out_data_129; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_130 = pipe3to8_io_pipe_phv_out_data_130; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_131 = pipe3to8_io_pipe_phv_out_data_131; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_132 = pipe3to8_io_pipe_phv_out_data_132; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_133 = pipe3to8_io_pipe_phv_out_data_133; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_134 = pipe3to8_io_pipe_phv_out_data_134; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_135 = pipe3to8_io_pipe_phv_out_data_135; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_136 = pipe3to8_io_pipe_phv_out_data_136; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_137 = pipe3to8_io_pipe_phv_out_data_137; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_138 = pipe3to8_io_pipe_phv_out_data_138; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_139 = pipe3to8_io_pipe_phv_out_data_139; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_140 = pipe3to8_io_pipe_phv_out_data_140; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_141 = pipe3to8_io_pipe_phv_out_data_141; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_142 = pipe3to8_io_pipe_phv_out_data_142; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_143 = pipe3to8_io_pipe_phv_out_data_143; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_144 = pipe3to8_io_pipe_phv_out_data_144; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_145 = pipe3to8_io_pipe_phv_out_data_145; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_146 = pipe3to8_io_pipe_phv_out_data_146; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_147 = pipe3to8_io_pipe_phv_out_data_147; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_148 = pipe3to8_io_pipe_phv_out_data_148; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_149 = pipe3to8_io_pipe_phv_out_data_149; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_150 = pipe3to8_io_pipe_phv_out_data_150; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_151 = pipe3to8_io_pipe_phv_out_data_151; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_152 = pipe3to8_io_pipe_phv_out_data_152; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_153 = pipe3to8_io_pipe_phv_out_data_153; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_154 = pipe3to8_io_pipe_phv_out_data_154; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_155 = pipe3to8_io_pipe_phv_out_data_155; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_156 = pipe3to8_io_pipe_phv_out_data_156; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_157 = pipe3to8_io_pipe_phv_out_data_157; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_158 = pipe3to8_io_pipe_phv_out_data_158; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_data_159 = pipe3to8_io_pipe_phv_out_data_159; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_0 = pipe3to8_io_pipe_phv_out_header_0; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_1 = pipe3to8_io_pipe_phv_out_header_1; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_2 = pipe3to8_io_pipe_phv_out_header_2; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_3 = pipe3to8_io_pipe_phv_out_header_3; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_4 = pipe3to8_io_pipe_phv_out_header_4; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_5 = pipe3to8_io_pipe_phv_out_header_5; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_6 = pipe3to8_io_pipe_phv_out_header_6; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_7 = pipe3to8_io_pipe_phv_out_header_7; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_8 = pipe3to8_io_pipe_phv_out_header_8; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_9 = pipe3to8_io_pipe_phv_out_header_9; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_10 = pipe3to8_io_pipe_phv_out_header_10; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_11 = pipe3to8_io_pipe_phv_out_header_11; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_12 = pipe3to8_io_pipe_phv_out_header_12; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_13 = pipe3to8_io_pipe_phv_out_header_13; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_14 = pipe3to8_io_pipe_phv_out_header_14; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_header_15 = pipe3to8_io_pipe_phv_out_header_15; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_current_state = pipe3to8_io_pipe_phv_out_parse_current_state; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_current_offset = pipe3to8_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_parse_transition_field = pipe3to8_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_next_processor_id = pipe3to8_io_pipe_phv_out_next_processor_id; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_next_config_id = pipe3to8_io_pipe_phv_out_next_config_id; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_is_valid_processor = pipe3to8_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_valid = pipe3to8_io_pipe_phv_out_valid; // @[matcher.scala 364:27]
  assign pipe9_io_pipe_phv_in_last = pipe3to8_io_pipe_phv_out_last; // @[matcher.scala 364:27]
  assign pipe10_clock = clock;
  assign pipe10_io_pipe_phv_in_data_0 = pipe9_io_pipe_phv_out_data_0; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_1 = pipe9_io_pipe_phv_out_data_1; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_2 = pipe9_io_pipe_phv_out_data_2; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_3 = pipe9_io_pipe_phv_out_data_3; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_4 = pipe9_io_pipe_phv_out_data_4; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_5 = pipe9_io_pipe_phv_out_data_5; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_6 = pipe9_io_pipe_phv_out_data_6; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_7 = pipe9_io_pipe_phv_out_data_7; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_8 = pipe9_io_pipe_phv_out_data_8; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_9 = pipe9_io_pipe_phv_out_data_9; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_10 = pipe9_io_pipe_phv_out_data_10; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_11 = pipe9_io_pipe_phv_out_data_11; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_12 = pipe9_io_pipe_phv_out_data_12; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_13 = pipe9_io_pipe_phv_out_data_13; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_14 = pipe9_io_pipe_phv_out_data_14; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_15 = pipe9_io_pipe_phv_out_data_15; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_16 = pipe9_io_pipe_phv_out_data_16; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_17 = pipe9_io_pipe_phv_out_data_17; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_18 = pipe9_io_pipe_phv_out_data_18; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_19 = pipe9_io_pipe_phv_out_data_19; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_20 = pipe9_io_pipe_phv_out_data_20; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_21 = pipe9_io_pipe_phv_out_data_21; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_22 = pipe9_io_pipe_phv_out_data_22; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_23 = pipe9_io_pipe_phv_out_data_23; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_24 = pipe9_io_pipe_phv_out_data_24; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_25 = pipe9_io_pipe_phv_out_data_25; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_26 = pipe9_io_pipe_phv_out_data_26; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_27 = pipe9_io_pipe_phv_out_data_27; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_28 = pipe9_io_pipe_phv_out_data_28; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_29 = pipe9_io_pipe_phv_out_data_29; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_30 = pipe9_io_pipe_phv_out_data_30; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_31 = pipe9_io_pipe_phv_out_data_31; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_32 = pipe9_io_pipe_phv_out_data_32; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_33 = pipe9_io_pipe_phv_out_data_33; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_34 = pipe9_io_pipe_phv_out_data_34; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_35 = pipe9_io_pipe_phv_out_data_35; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_36 = pipe9_io_pipe_phv_out_data_36; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_37 = pipe9_io_pipe_phv_out_data_37; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_38 = pipe9_io_pipe_phv_out_data_38; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_39 = pipe9_io_pipe_phv_out_data_39; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_40 = pipe9_io_pipe_phv_out_data_40; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_41 = pipe9_io_pipe_phv_out_data_41; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_42 = pipe9_io_pipe_phv_out_data_42; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_43 = pipe9_io_pipe_phv_out_data_43; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_44 = pipe9_io_pipe_phv_out_data_44; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_45 = pipe9_io_pipe_phv_out_data_45; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_46 = pipe9_io_pipe_phv_out_data_46; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_47 = pipe9_io_pipe_phv_out_data_47; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_48 = pipe9_io_pipe_phv_out_data_48; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_49 = pipe9_io_pipe_phv_out_data_49; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_50 = pipe9_io_pipe_phv_out_data_50; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_51 = pipe9_io_pipe_phv_out_data_51; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_52 = pipe9_io_pipe_phv_out_data_52; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_53 = pipe9_io_pipe_phv_out_data_53; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_54 = pipe9_io_pipe_phv_out_data_54; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_55 = pipe9_io_pipe_phv_out_data_55; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_56 = pipe9_io_pipe_phv_out_data_56; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_57 = pipe9_io_pipe_phv_out_data_57; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_58 = pipe9_io_pipe_phv_out_data_58; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_59 = pipe9_io_pipe_phv_out_data_59; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_60 = pipe9_io_pipe_phv_out_data_60; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_61 = pipe9_io_pipe_phv_out_data_61; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_62 = pipe9_io_pipe_phv_out_data_62; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_63 = pipe9_io_pipe_phv_out_data_63; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_64 = pipe9_io_pipe_phv_out_data_64; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_65 = pipe9_io_pipe_phv_out_data_65; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_66 = pipe9_io_pipe_phv_out_data_66; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_67 = pipe9_io_pipe_phv_out_data_67; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_68 = pipe9_io_pipe_phv_out_data_68; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_69 = pipe9_io_pipe_phv_out_data_69; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_70 = pipe9_io_pipe_phv_out_data_70; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_71 = pipe9_io_pipe_phv_out_data_71; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_72 = pipe9_io_pipe_phv_out_data_72; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_73 = pipe9_io_pipe_phv_out_data_73; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_74 = pipe9_io_pipe_phv_out_data_74; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_75 = pipe9_io_pipe_phv_out_data_75; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_76 = pipe9_io_pipe_phv_out_data_76; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_77 = pipe9_io_pipe_phv_out_data_77; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_78 = pipe9_io_pipe_phv_out_data_78; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_79 = pipe9_io_pipe_phv_out_data_79; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_80 = pipe9_io_pipe_phv_out_data_80; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_81 = pipe9_io_pipe_phv_out_data_81; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_82 = pipe9_io_pipe_phv_out_data_82; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_83 = pipe9_io_pipe_phv_out_data_83; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_84 = pipe9_io_pipe_phv_out_data_84; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_85 = pipe9_io_pipe_phv_out_data_85; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_86 = pipe9_io_pipe_phv_out_data_86; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_87 = pipe9_io_pipe_phv_out_data_87; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_88 = pipe9_io_pipe_phv_out_data_88; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_89 = pipe9_io_pipe_phv_out_data_89; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_90 = pipe9_io_pipe_phv_out_data_90; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_91 = pipe9_io_pipe_phv_out_data_91; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_92 = pipe9_io_pipe_phv_out_data_92; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_93 = pipe9_io_pipe_phv_out_data_93; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_94 = pipe9_io_pipe_phv_out_data_94; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_95 = pipe9_io_pipe_phv_out_data_95; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_96 = pipe9_io_pipe_phv_out_data_96; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_97 = pipe9_io_pipe_phv_out_data_97; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_98 = pipe9_io_pipe_phv_out_data_98; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_99 = pipe9_io_pipe_phv_out_data_99; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_100 = pipe9_io_pipe_phv_out_data_100; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_101 = pipe9_io_pipe_phv_out_data_101; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_102 = pipe9_io_pipe_phv_out_data_102; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_103 = pipe9_io_pipe_phv_out_data_103; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_104 = pipe9_io_pipe_phv_out_data_104; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_105 = pipe9_io_pipe_phv_out_data_105; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_106 = pipe9_io_pipe_phv_out_data_106; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_107 = pipe9_io_pipe_phv_out_data_107; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_108 = pipe9_io_pipe_phv_out_data_108; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_109 = pipe9_io_pipe_phv_out_data_109; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_110 = pipe9_io_pipe_phv_out_data_110; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_111 = pipe9_io_pipe_phv_out_data_111; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_112 = pipe9_io_pipe_phv_out_data_112; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_113 = pipe9_io_pipe_phv_out_data_113; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_114 = pipe9_io_pipe_phv_out_data_114; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_115 = pipe9_io_pipe_phv_out_data_115; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_116 = pipe9_io_pipe_phv_out_data_116; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_117 = pipe9_io_pipe_phv_out_data_117; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_118 = pipe9_io_pipe_phv_out_data_118; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_119 = pipe9_io_pipe_phv_out_data_119; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_120 = pipe9_io_pipe_phv_out_data_120; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_121 = pipe9_io_pipe_phv_out_data_121; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_122 = pipe9_io_pipe_phv_out_data_122; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_123 = pipe9_io_pipe_phv_out_data_123; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_124 = pipe9_io_pipe_phv_out_data_124; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_125 = pipe9_io_pipe_phv_out_data_125; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_126 = pipe9_io_pipe_phv_out_data_126; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_127 = pipe9_io_pipe_phv_out_data_127; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_128 = pipe9_io_pipe_phv_out_data_128; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_129 = pipe9_io_pipe_phv_out_data_129; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_130 = pipe9_io_pipe_phv_out_data_130; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_131 = pipe9_io_pipe_phv_out_data_131; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_132 = pipe9_io_pipe_phv_out_data_132; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_133 = pipe9_io_pipe_phv_out_data_133; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_134 = pipe9_io_pipe_phv_out_data_134; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_135 = pipe9_io_pipe_phv_out_data_135; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_136 = pipe9_io_pipe_phv_out_data_136; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_137 = pipe9_io_pipe_phv_out_data_137; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_138 = pipe9_io_pipe_phv_out_data_138; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_139 = pipe9_io_pipe_phv_out_data_139; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_140 = pipe9_io_pipe_phv_out_data_140; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_141 = pipe9_io_pipe_phv_out_data_141; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_142 = pipe9_io_pipe_phv_out_data_142; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_143 = pipe9_io_pipe_phv_out_data_143; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_144 = pipe9_io_pipe_phv_out_data_144; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_145 = pipe9_io_pipe_phv_out_data_145; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_146 = pipe9_io_pipe_phv_out_data_146; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_147 = pipe9_io_pipe_phv_out_data_147; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_148 = pipe9_io_pipe_phv_out_data_148; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_149 = pipe9_io_pipe_phv_out_data_149; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_150 = pipe9_io_pipe_phv_out_data_150; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_151 = pipe9_io_pipe_phv_out_data_151; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_152 = pipe9_io_pipe_phv_out_data_152; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_153 = pipe9_io_pipe_phv_out_data_153; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_154 = pipe9_io_pipe_phv_out_data_154; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_155 = pipe9_io_pipe_phv_out_data_155; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_156 = pipe9_io_pipe_phv_out_data_156; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_157 = pipe9_io_pipe_phv_out_data_157; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_158 = pipe9_io_pipe_phv_out_data_158; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_data_159 = pipe9_io_pipe_phv_out_data_159; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_0 = pipe9_io_pipe_phv_out_header_0; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_1 = pipe9_io_pipe_phv_out_header_1; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_2 = pipe9_io_pipe_phv_out_header_2; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_3 = pipe9_io_pipe_phv_out_header_3; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_4 = pipe9_io_pipe_phv_out_header_4; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_5 = pipe9_io_pipe_phv_out_header_5; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_6 = pipe9_io_pipe_phv_out_header_6; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_7 = pipe9_io_pipe_phv_out_header_7; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_8 = pipe9_io_pipe_phv_out_header_8; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_9 = pipe9_io_pipe_phv_out_header_9; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_10 = pipe9_io_pipe_phv_out_header_10; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_11 = pipe9_io_pipe_phv_out_header_11; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_12 = pipe9_io_pipe_phv_out_header_12; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_13 = pipe9_io_pipe_phv_out_header_13; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_14 = pipe9_io_pipe_phv_out_header_14; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_header_15 = pipe9_io_pipe_phv_out_header_15; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_current_state = pipe9_io_pipe_phv_out_parse_current_state; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_current_offset = pipe9_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_parse_transition_field = pipe9_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_next_processor_id = pipe9_io_pipe_phv_out_next_processor_id; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_next_config_id = pipe9_io_pipe_phv_out_next_config_id; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_is_valid_processor = pipe9_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_valid = pipe9_io_pipe_phv_out_valid; // @[matcher.scala 370:27]
  assign pipe10_io_pipe_phv_in_last = pipe9_io_pipe_phv_out_last; // @[matcher.scala 370:27]
  assign pipe11_clock = clock;
  assign pipe11_io_pipe_phv_in_data_0 = pipe10_io_pipe_phv_out_data_0; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_1 = pipe10_io_pipe_phv_out_data_1; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_2 = pipe10_io_pipe_phv_out_data_2; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_3 = pipe10_io_pipe_phv_out_data_3; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_4 = pipe10_io_pipe_phv_out_data_4; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_5 = pipe10_io_pipe_phv_out_data_5; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_6 = pipe10_io_pipe_phv_out_data_6; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_7 = pipe10_io_pipe_phv_out_data_7; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_8 = pipe10_io_pipe_phv_out_data_8; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_9 = pipe10_io_pipe_phv_out_data_9; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_10 = pipe10_io_pipe_phv_out_data_10; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_11 = pipe10_io_pipe_phv_out_data_11; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_12 = pipe10_io_pipe_phv_out_data_12; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_13 = pipe10_io_pipe_phv_out_data_13; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_14 = pipe10_io_pipe_phv_out_data_14; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_15 = pipe10_io_pipe_phv_out_data_15; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_16 = pipe10_io_pipe_phv_out_data_16; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_17 = pipe10_io_pipe_phv_out_data_17; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_18 = pipe10_io_pipe_phv_out_data_18; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_19 = pipe10_io_pipe_phv_out_data_19; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_20 = pipe10_io_pipe_phv_out_data_20; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_21 = pipe10_io_pipe_phv_out_data_21; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_22 = pipe10_io_pipe_phv_out_data_22; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_23 = pipe10_io_pipe_phv_out_data_23; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_24 = pipe10_io_pipe_phv_out_data_24; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_25 = pipe10_io_pipe_phv_out_data_25; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_26 = pipe10_io_pipe_phv_out_data_26; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_27 = pipe10_io_pipe_phv_out_data_27; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_28 = pipe10_io_pipe_phv_out_data_28; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_29 = pipe10_io_pipe_phv_out_data_29; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_30 = pipe10_io_pipe_phv_out_data_30; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_31 = pipe10_io_pipe_phv_out_data_31; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_32 = pipe10_io_pipe_phv_out_data_32; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_33 = pipe10_io_pipe_phv_out_data_33; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_34 = pipe10_io_pipe_phv_out_data_34; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_35 = pipe10_io_pipe_phv_out_data_35; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_36 = pipe10_io_pipe_phv_out_data_36; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_37 = pipe10_io_pipe_phv_out_data_37; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_38 = pipe10_io_pipe_phv_out_data_38; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_39 = pipe10_io_pipe_phv_out_data_39; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_40 = pipe10_io_pipe_phv_out_data_40; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_41 = pipe10_io_pipe_phv_out_data_41; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_42 = pipe10_io_pipe_phv_out_data_42; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_43 = pipe10_io_pipe_phv_out_data_43; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_44 = pipe10_io_pipe_phv_out_data_44; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_45 = pipe10_io_pipe_phv_out_data_45; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_46 = pipe10_io_pipe_phv_out_data_46; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_47 = pipe10_io_pipe_phv_out_data_47; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_48 = pipe10_io_pipe_phv_out_data_48; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_49 = pipe10_io_pipe_phv_out_data_49; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_50 = pipe10_io_pipe_phv_out_data_50; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_51 = pipe10_io_pipe_phv_out_data_51; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_52 = pipe10_io_pipe_phv_out_data_52; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_53 = pipe10_io_pipe_phv_out_data_53; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_54 = pipe10_io_pipe_phv_out_data_54; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_55 = pipe10_io_pipe_phv_out_data_55; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_56 = pipe10_io_pipe_phv_out_data_56; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_57 = pipe10_io_pipe_phv_out_data_57; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_58 = pipe10_io_pipe_phv_out_data_58; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_59 = pipe10_io_pipe_phv_out_data_59; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_60 = pipe10_io_pipe_phv_out_data_60; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_61 = pipe10_io_pipe_phv_out_data_61; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_62 = pipe10_io_pipe_phv_out_data_62; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_63 = pipe10_io_pipe_phv_out_data_63; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_64 = pipe10_io_pipe_phv_out_data_64; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_65 = pipe10_io_pipe_phv_out_data_65; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_66 = pipe10_io_pipe_phv_out_data_66; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_67 = pipe10_io_pipe_phv_out_data_67; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_68 = pipe10_io_pipe_phv_out_data_68; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_69 = pipe10_io_pipe_phv_out_data_69; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_70 = pipe10_io_pipe_phv_out_data_70; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_71 = pipe10_io_pipe_phv_out_data_71; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_72 = pipe10_io_pipe_phv_out_data_72; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_73 = pipe10_io_pipe_phv_out_data_73; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_74 = pipe10_io_pipe_phv_out_data_74; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_75 = pipe10_io_pipe_phv_out_data_75; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_76 = pipe10_io_pipe_phv_out_data_76; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_77 = pipe10_io_pipe_phv_out_data_77; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_78 = pipe10_io_pipe_phv_out_data_78; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_79 = pipe10_io_pipe_phv_out_data_79; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_80 = pipe10_io_pipe_phv_out_data_80; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_81 = pipe10_io_pipe_phv_out_data_81; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_82 = pipe10_io_pipe_phv_out_data_82; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_83 = pipe10_io_pipe_phv_out_data_83; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_84 = pipe10_io_pipe_phv_out_data_84; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_85 = pipe10_io_pipe_phv_out_data_85; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_86 = pipe10_io_pipe_phv_out_data_86; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_87 = pipe10_io_pipe_phv_out_data_87; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_88 = pipe10_io_pipe_phv_out_data_88; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_89 = pipe10_io_pipe_phv_out_data_89; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_90 = pipe10_io_pipe_phv_out_data_90; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_91 = pipe10_io_pipe_phv_out_data_91; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_92 = pipe10_io_pipe_phv_out_data_92; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_93 = pipe10_io_pipe_phv_out_data_93; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_94 = pipe10_io_pipe_phv_out_data_94; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_95 = pipe10_io_pipe_phv_out_data_95; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_96 = pipe10_io_pipe_phv_out_data_96; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_97 = pipe10_io_pipe_phv_out_data_97; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_98 = pipe10_io_pipe_phv_out_data_98; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_99 = pipe10_io_pipe_phv_out_data_99; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_100 = pipe10_io_pipe_phv_out_data_100; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_101 = pipe10_io_pipe_phv_out_data_101; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_102 = pipe10_io_pipe_phv_out_data_102; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_103 = pipe10_io_pipe_phv_out_data_103; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_104 = pipe10_io_pipe_phv_out_data_104; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_105 = pipe10_io_pipe_phv_out_data_105; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_106 = pipe10_io_pipe_phv_out_data_106; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_107 = pipe10_io_pipe_phv_out_data_107; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_108 = pipe10_io_pipe_phv_out_data_108; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_109 = pipe10_io_pipe_phv_out_data_109; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_110 = pipe10_io_pipe_phv_out_data_110; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_111 = pipe10_io_pipe_phv_out_data_111; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_112 = pipe10_io_pipe_phv_out_data_112; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_113 = pipe10_io_pipe_phv_out_data_113; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_114 = pipe10_io_pipe_phv_out_data_114; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_115 = pipe10_io_pipe_phv_out_data_115; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_116 = pipe10_io_pipe_phv_out_data_116; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_117 = pipe10_io_pipe_phv_out_data_117; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_118 = pipe10_io_pipe_phv_out_data_118; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_119 = pipe10_io_pipe_phv_out_data_119; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_120 = pipe10_io_pipe_phv_out_data_120; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_121 = pipe10_io_pipe_phv_out_data_121; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_122 = pipe10_io_pipe_phv_out_data_122; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_123 = pipe10_io_pipe_phv_out_data_123; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_124 = pipe10_io_pipe_phv_out_data_124; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_125 = pipe10_io_pipe_phv_out_data_125; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_126 = pipe10_io_pipe_phv_out_data_126; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_127 = pipe10_io_pipe_phv_out_data_127; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_128 = pipe10_io_pipe_phv_out_data_128; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_129 = pipe10_io_pipe_phv_out_data_129; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_130 = pipe10_io_pipe_phv_out_data_130; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_131 = pipe10_io_pipe_phv_out_data_131; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_132 = pipe10_io_pipe_phv_out_data_132; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_133 = pipe10_io_pipe_phv_out_data_133; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_134 = pipe10_io_pipe_phv_out_data_134; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_135 = pipe10_io_pipe_phv_out_data_135; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_136 = pipe10_io_pipe_phv_out_data_136; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_137 = pipe10_io_pipe_phv_out_data_137; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_138 = pipe10_io_pipe_phv_out_data_138; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_139 = pipe10_io_pipe_phv_out_data_139; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_140 = pipe10_io_pipe_phv_out_data_140; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_141 = pipe10_io_pipe_phv_out_data_141; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_142 = pipe10_io_pipe_phv_out_data_142; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_143 = pipe10_io_pipe_phv_out_data_143; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_144 = pipe10_io_pipe_phv_out_data_144; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_145 = pipe10_io_pipe_phv_out_data_145; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_146 = pipe10_io_pipe_phv_out_data_146; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_147 = pipe10_io_pipe_phv_out_data_147; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_148 = pipe10_io_pipe_phv_out_data_148; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_149 = pipe10_io_pipe_phv_out_data_149; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_150 = pipe10_io_pipe_phv_out_data_150; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_151 = pipe10_io_pipe_phv_out_data_151; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_152 = pipe10_io_pipe_phv_out_data_152; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_153 = pipe10_io_pipe_phv_out_data_153; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_154 = pipe10_io_pipe_phv_out_data_154; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_155 = pipe10_io_pipe_phv_out_data_155; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_156 = pipe10_io_pipe_phv_out_data_156; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_157 = pipe10_io_pipe_phv_out_data_157; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_158 = pipe10_io_pipe_phv_out_data_158; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_data_159 = pipe10_io_pipe_phv_out_data_159; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_0 = pipe10_io_pipe_phv_out_header_0; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_1 = pipe10_io_pipe_phv_out_header_1; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_2 = pipe10_io_pipe_phv_out_header_2; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_3 = pipe10_io_pipe_phv_out_header_3; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_4 = pipe10_io_pipe_phv_out_header_4; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_5 = pipe10_io_pipe_phv_out_header_5; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_6 = pipe10_io_pipe_phv_out_header_6; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_7 = pipe10_io_pipe_phv_out_header_7; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_8 = pipe10_io_pipe_phv_out_header_8; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_9 = pipe10_io_pipe_phv_out_header_9; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_10 = pipe10_io_pipe_phv_out_header_10; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_11 = pipe10_io_pipe_phv_out_header_11; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_12 = pipe10_io_pipe_phv_out_header_12; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_13 = pipe10_io_pipe_phv_out_header_13; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_14 = pipe10_io_pipe_phv_out_header_14; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_header_15 = pipe10_io_pipe_phv_out_header_15; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_current_state = pipe10_io_pipe_phv_out_parse_current_state; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_current_offset = pipe10_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_parse_transition_field = pipe10_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_next_processor_id = pipe10_io_pipe_phv_out_next_processor_id; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_next_config_id = pipe10_io_pipe_phv_out_next_config_id; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_is_valid_processor = pipe10_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_valid = pipe10_io_pipe_phv_out_valid; // @[matcher.scala 377:27]
  assign pipe11_io_pipe_phv_in_last = pipe10_io_pipe_phv_out_last; // @[matcher.scala 377:27]
  assign pipe12_clock = clock;
  assign pipe12_io_pipe_phv_in_data_0 = pipe11_io_pipe_phv_out_data_0; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_1 = pipe11_io_pipe_phv_out_data_1; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_2 = pipe11_io_pipe_phv_out_data_2; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_3 = pipe11_io_pipe_phv_out_data_3; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_4 = pipe11_io_pipe_phv_out_data_4; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_5 = pipe11_io_pipe_phv_out_data_5; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_6 = pipe11_io_pipe_phv_out_data_6; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_7 = pipe11_io_pipe_phv_out_data_7; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_8 = pipe11_io_pipe_phv_out_data_8; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_9 = pipe11_io_pipe_phv_out_data_9; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_10 = pipe11_io_pipe_phv_out_data_10; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_11 = pipe11_io_pipe_phv_out_data_11; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_12 = pipe11_io_pipe_phv_out_data_12; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_13 = pipe11_io_pipe_phv_out_data_13; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_14 = pipe11_io_pipe_phv_out_data_14; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_15 = pipe11_io_pipe_phv_out_data_15; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_16 = pipe11_io_pipe_phv_out_data_16; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_17 = pipe11_io_pipe_phv_out_data_17; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_18 = pipe11_io_pipe_phv_out_data_18; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_19 = pipe11_io_pipe_phv_out_data_19; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_20 = pipe11_io_pipe_phv_out_data_20; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_21 = pipe11_io_pipe_phv_out_data_21; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_22 = pipe11_io_pipe_phv_out_data_22; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_23 = pipe11_io_pipe_phv_out_data_23; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_24 = pipe11_io_pipe_phv_out_data_24; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_25 = pipe11_io_pipe_phv_out_data_25; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_26 = pipe11_io_pipe_phv_out_data_26; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_27 = pipe11_io_pipe_phv_out_data_27; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_28 = pipe11_io_pipe_phv_out_data_28; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_29 = pipe11_io_pipe_phv_out_data_29; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_30 = pipe11_io_pipe_phv_out_data_30; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_31 = pipe11_io_pipe_phv_out_data_31; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_32 = pipe11_io_pipe_phv_out_data_32; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_33 = pipe11_io_pipe_phv_out_data_33; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_34 = pipe11_io_pipe_phv_out_data_34; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_35 = pipe11_io_pipe_phv_out_data_35; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_36 = pipe11_io_pipe_phv_out_data_36; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_37 = pipe11_io_pipe_phv_out_data_37; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_38 = pipe11_io_pipe_phv_out_data_38; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_39 = pipe11_io_pipe_phv_out_data_39; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_40 = pipe11_io_pipe_phv_out_data_40; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_41 = pipe11_io_pipe_phv_out_data_41; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_42 = pipe11_io_pipe_phv_out_data_42; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_43 = pipe11_io_pipe_phv_out_data_43; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_44 = pipe11_io_pipe_phv_out_data_44; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_45 = pipe11_io_pipe_phv_out_data_45; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_46 = pipe11_io_pipe_phv_out_data_46; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_47 = pipe11_io_pipe_phv_out_data_47; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_48 = pipe11_io_pipe_phv_out_data_48; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_49 = pipe11_io_pipe_phv_out_data_49; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_50 = pipe11_io_pipe_phv_out_data_50; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_51 = pipe11_io_pipe_phv_out_data_51; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_52 = pipe11_io_pipe_phv_out_data_52; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_53 = pipe11_io_pipe_phv_out_data_53; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_54 = pipe11_io_pipe_phv_out_data_54; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_55 = pipe11_io_pipe_phv_out_data_55; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_56 = pipe11_io_pipe_phv_out_data_56; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_57 = pipe11_io_pipe_phv_out_data_57; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_58 = pipe11_io_pipe_phv_out_data_58; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_59 = pipe11_io_pipe_phv_out_data_59; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_60 = pipe11_io_pipe_phv_out_data_60; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_61 = pipe11_io_pipe_phv_out_data_61; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_62 = pipe11_io_pipe_phv_out_data_62; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_63 = pipe11_io_pipe_phv_out_data_63; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_64 = pipe11_io_pipe_phv_out_data_64; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_65 = pipe11_io_pipe_phv_out_data_65; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_66 = pipe11_io_pipe_phv_out_data_66; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_67 = pipe11_io_pipe_phv_out_data_67; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_68 = pipe11_io_pipe_phv_out_data_68; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_69 = pipe11_io_pipe_phv_out_data_69; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_70 = pipe11_io_pipe_phv_out_data_70; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_71 = pipe11_io_pipe_phv_out_data_71; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_72 = pipe11_io_pipe_phv_out_data_72; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_73 = pipe11_io_pipe_phv_out_data_73; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_74 = pipe11_io_pipe_phv_out_data_74; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_75 = pipe11_io_pipe_phv_out_data_75; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_76 = pipe11_io_pipe_phv_out_data_76; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_77 = pipe11_io_pipe_phv_out_data_77; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_78 = pipe11_io_pipe_phv_out_data_78; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_79 = pipe11_io_pipe_phv_out_data_79; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_80 = pipe11_io_pipe_phv_out_data_80; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_81 = pipe11_io_pipe_phv_out_data_81; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_82 = pipe11_io_pipe_phv_out_data_82; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_83 = pipe11_io_pipe_phv_out_data_83; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_84 = pipe11_io_pipe_phv_out_data_84; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_85 = pipe11_io_pipe_phv_out_data_85; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_86 = pipe11_io_pipe_phv_out_data_86; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_87 = pipe11_io_pipe_phv_out_data_87; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_88 = pipe11_io_pipe_phv_out_data_88; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_89 = pipe11_io_pipe_phv_out_data_89; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_90 = pipe11_io_pipe_phv_out_data_90; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_91 = pipe11_io_pipe_phv_out_data_91; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_92 = pipe11_io_pipe_phv_out_data_92; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_93 = pipe11_io_pipe_phv_out_data_93; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_94 = pipe11_io_pipe_phv_out_data_94; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_95 = pipe11_io_pipe_phv_out_data_95; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_96 = pipe11_io_pipe_phv_out_data_96; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_97 = pipe11_io_pipe_phv_out_data_97; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_98 = pipe11_io_pipe_phv_out_data_98; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_99 = pipe11_io_pipe_phv_out_data_99; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_100 = pipe11_io_pipe_phv_out_data_100; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_101 = pipe11_io_pipe_phv_out_data_101; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_102 = pipe11_io_pipe_phv_out_data_102; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_103 = pipe11_io_pipe_phv_out_data_103; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_104 = pipe11_io_pipe_phv_out_data_104; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_105 = pipe11_io_pipe_phv_out_data_105; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_106 = pipe11_io_pipe_phv_out_data_106; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_107 = pipe11_io_pipe_phv_out_data_107; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_108 = pipe11_io_pipe_phv_out_data_108; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_109 = pipe11_io_pipe_phv_out_data_109; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_110 = pipe11_io_pipe_phv_out_data_110; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_111 = pipe11_io_pipe_phv_out_data_111; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_112 = pipe11_io_pipe_phv_out_data_112; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_113 = pipe11_io_pipe_phv_out_data_113; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_114 = pipe11_io_pipe_phv_out_data_114; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_115 = pipe11_io_pipe_phv_out_data_115; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_116 = pipe11_io_pipe_phv_out_data_116; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_117 = pipe11_io_pipe_phv_out_data_117; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_118 = pipe11_io_pipe_phv_out_data_118; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_119 = pipe11_io_pipe_phv_out_data_119; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_120 = pipe11_io_pipe_phv_out_data_120; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_121 = pipe11_io_pipe_phv_out_data_121; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_122 = pipe11_io_pipe_phv_out_data_122; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_123 = pipe11_io_pipe_phv_out_data_123; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_124 = pipe11_io_pipe_phv_out_data_124; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_125 = pipe11_io_pipe_phv_out_data_125; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_126 = pipe11_io_pipe_phv_out_data_126; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_127 = pipe11_io_pipe_phv_out_data_127; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_128 = pipe11_io_pipe_phv_out_data_128; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_129 = pipe11_io_pipe_phv_out_data_129; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_130 = pipe11_io_pipe_phv_out_data_130; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_131 = pipe11_io_pipe_phv_out_data_131; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_132 = pipe11_io_pipe_phv_out_data_132; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_133 = pipe11_io_pipe_phv_out_data_133; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_134 = pipe11_io_pipe_phv_out_data_134; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_135 = pipe11_io_pipe_phv_out_data_135; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_136 = pipe11_io_pipe_phv_out_data_136; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_137 = pipe11_io_pipe_phv_out_data_137; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_138 = pipe11_io_pipe_phv_out_data_138; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_139 = pipe11_io_pipe_phv_out_data_139; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_140 = pipe11_io_pipe_phv_out_data_140; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_141 = pipe11_io_pipe_phv_out_data_141; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_142 = pipe11_io_pipe_phv_out_data_142; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_143 = pipe11_io_pipe_phv_out_data_143; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_144 = pipe11_io_pipe_phv_out_data_144; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_145 = pipe11_io_pipe_phv_out_data_145; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_146 = pipe11_io_pipe_phv_out_data_146; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_147 = pipe11_io_pipe_phv_out_data_147; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_148 = pipe11_io_pipe_phv_out_data_148; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_149 = pipe11_io_pipe_phv_out_data_149; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_150 = pipe11_io_pipe_phv_out_data_150; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_151 = pipe11_io_pipe_phv_out_data_151; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_152 = pipe11_io_pipe_phv_out_data_152; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_153 = pipe11_io_pipe_phv_out_data_153; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_154 = pipe11_io_pipe_phv_out_data_154; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_155 = pipe11_io_pipe_phv_out_data_155; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_156 = pipe11_io_pipe_phv_out_data_156; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_157 = pipe11_io_pipe_phv_out_data_157; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_158 = pipe11_io_pipe_phv_out_data_158; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_data_159 = pipe11_io_pipe_phv_out_data_159; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_0 = pipe11_io_pipe_phv_out_header_0; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_1 = pipe11_io_pipe_phv_out_header_1; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_2 = pipe11_io_pipe_phv_out_header_2; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_3 = pipe11_io_pipe_phv_out_header_3; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_4 = pipe11_io_pipe_phv_out_header_4; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_5 = pipe11_io_pipe_phv_out_header_5; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_6 = pipe11_io_pipe_phv_out_header_6; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_7 = pipe11_io_pipe_phv_out_header_7; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_8 = pipe11_io_pipe_phv_out_header_8; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_9 = pipe11_io_pipe_phv_out_header_9; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_10 = pipe11_io_pipe_phv_out_header_10; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_11 = pipe11_io_pipe_phv_out_header_11; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_12 = pipe11_io_pipe_phv_out_header_12; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_13 = pipe11_io_pipe_phv_out_header_13; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_14 = pipe11_io_pipe_phv_out_header_14; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_header_15 = pipe11_io_pipe_phv_out_header_15; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_current_state = pipe11_io_pipe_phv_out_parse_current_state; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_current_offset = pipe11_io_pipe_phv_out_parse_current_offset; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_parse_transition_field = pipe11_io_pipe_phv_out_parse_transition_field; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_next_processor_id = pipe11_io_pipe_phv_out_next_processor_id; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_next_config_id = pipe11_io_pipe_phv_out_next_config_id; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_is_valid_processor = pipe11_io_pipe_phv_out_is_valid_processor; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_valid = pipe11_io_pipe_phv_out_valid; // @[matcher.scala 383:27]
  assign pipe12_io_pipe_phv_in_last = pipe11_io_pipe_phv_out_last; // @[matcher.scala 383:27]
endmodule
