module PrimitiveGetSource(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  input  [7:0]  io_offset_in_0,
  input  [7:0]  io_offset_in_1,
  input  [7:0]  io_offset_in_2,
  input  [7:0]  io_offset_in_3,
  input  [7:0]  io_length_in_0,
  input  [7:0]  io_length_in_1,
  input  [7:0]  io_length_in_2,
  input  [7:0]  io_length_in_3,
  output [31:0] io_vliw_out_0,
  output [31:0] io_vliw_out_1,
  output [31:0] io_vliw_out_2,
  output [31:0] io_vliw_out_3,
  output [31:0] io_field_out_0,
  output [31:0] io_field_out_1,
  output [31:0] io_field_out_2,
  output [31:0] io_field_out_3,
  output [3:0]  io_mask_out_0,
  output [3:0]  io_mask_out_1,
  output [3:0]  io_mask_out_2,
  output [3:0]  io_mask_out_3,
  output [1:0]  io_bias_out_0,
  output [1:0]  io_bias_out_1,
  output [1:0]  io_bias_out_2,
  output [1:0]  io_bias_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor.scala 151:22]
  reg [7:0] phv_data_1; // @[executor.scala 151:22]
  reg [7:0] phv_data_2; // @[executor.scala 151:22]
  reg [7:0] phv_data_3; // @[executor.scala 151:22]
  reg [7:0] phv_data_4; // @[executor.scala 151:22]
  reg [7:0] phv_data_5; // @[executor.scala 151:22]
  reg [7:0] phv_data_6; // @[executor.scala 151:22]
  reg [7:0] phv_data_7; // @[executor.scala 151:22]
  reg [7:0] phv_data_8; // @[executor.scala 151:22]
  reg [7:0] phv_data_9; // @[executor.scala 151:22]
  reg [7:0] phv_data_10; // @[executor.scala 151:22]
  reg [7:0] phv_data_11; // @[executor.scala 151:22]
  reg [7:0] phv_data_12; // @[executor.scala 151:22]
  reg [7:0] phv_data_13; // @[executor.scala 151:22]
  reg [7:0] phv_data_14; // @[executor.scala 151:22]
  reg [7:0] phv_data_15; // @[executor.scala 151:22]
  reg [7:0] phv_data_16; // @[executor.scala 151:22]
  reg [7:0] phv_data_17; // @[executor.scala 151:22]
  reg [7:0] phv_data_18; // @[executor.scala 151:22]
  reg [7:0] phv_data_19; // @[executor.scala 151:22]
  reg [7:0] phv_data_20; // @[executor.scala 151:22]
  reg [7:0] phv_data_21; // @[executor.scala 151:22]
  reg [7:0] phv_data_22; // @[executor.scala 151:22]
  reg [7:0] phv_data_23; // @[executor.scala 151:22]
  reg [7:0] phv_data_24; // @[executor.scala 151:22]
  reg [7:0] phv_data_25; // @[executor.scala 151:22]
  reg [7:0] phv_data_26; // @[executor.scala 151:22]
  reg [7:0] phv_data_27; // @[executor.scala 151:22]
  reg [7:0] phv_data_28; // @[executor.scala 151:22]
  reg [7:0] phv_data_29; // @[executor.scala 151:22]
  reg [7:0] phv_data_30; // @[executor.scala 151:22]
  reg [7:0] phv_data_31; // @[executor.scala 151:22]
  reg [7:0] phv_data_32; // @[executor.scala 151:22]
  reg [7:0] phv_data_33; // @[executor.scala 151:22]
  reg [7:0] phv_data_34; // @[executor.scala 151:22]
  reg [7:0] phv_data_35; // @[executor.scala 151:22]
  reg [7:0] phv_data_36; // @[executor.scala 151:22]
  reg [7:0] phv_data_37; // @[executor.scala 151:22]
  reg [7:0] phv_data_38; // @[executor.scala 151:22]
  reg [7:0] phv_data_39; // @[executor.scala 151:22]
  reg [7:0] phv_data_40; // @[executor.scala 151:22]
  reg [7:0] phv_data_41; // @[executor.scala 151:22]
  reg [7:0] phv_data_42; // @[executor.scala 151:22]
  reg [7:0] phv_data_43; // @[executor.scala 151:22]
  reg [7:0] phv_data_44; // @[executor.scala 151:22]
  reg [7:0] phv_data_45; // @[executor.scala 151:22]
  reg [7:0] phv_data_46; // @[executor.scala 151:22]
  reg [7:0] phv_data_47; // @[executor.scala 151:22]
  reg [7:0] phv_data_48; // @[executor.scala 151:22]
  reg [7:0] phv_data_49; // @[executor.scala 151:22]
  reg [7:0] phv_data_50; // @[executor.scala 151:22]
  reg [7:0] phv_data_51; // @[executor.scala 151:22]
  reg [7:0] phv_data_52; // @[executor.scala 151:22]
  reg [7:0] phv_data_53; // @[executor.scala 151:22]
  reg [7:0] phv_data_54; // @[executor.scala 151:22]
  reg [7:0] phv_data_55; // @[executor.scala 151:22]
  reg [7:0] phv_data_56; // @[executor.scala 151:22]
  reg [7:0] phv_data_57; // @[executor.scala 151:22]
  reg [7:0] phv_data_58; // @[executor.scala 151:22]
  reg [7:0] phv_data_59; // @[executor.scala 151:22]
  reg [7:0] phv_data_60; // @[executor.scala 151:22]
  reg [7:0] phv_data_61; // @[executor.scala 151:22]
  reg [7:0] phv_data_62; // @[executor.scala 151:22]
  reg [7:0] phv_data_63; // @[executor.scala 151:22]
  reg [7:0] phv_data_64; // @[executor.scala 151:22]
  reg [7:0] phv_data_65; // @[executor.scala 151:22]
  reg [7:0] phv_data_66; // @[executor.scala 151:22]
  reg [7:0] phv_data_67; // @[executor.scala 151:22]
  reg [7:0] phv_data_68; // @[executor.scala 151:22]
  reg [7:0] phv_data_69; // @[executor.scala 151:22]
  reg [7:0] phv_data_70; // @[executor.scala 151:22]
  reg [7:0] phv_data_71; // @[executor.scala 151:22]
  reg [7:0] phv_data_72; // @[executor.scala 151:22]
  reg [7:0] phv_data_73; // @[executor.scala 151:22]
  reg [7:0] phv_data_74; // @[executor.scala 151:22]
  reg [7:0] phv_data_75; // @[executor.scala 151:22]
  reg [7:0] phv_data_76; // @[executor.scala 151:22]
  reg [7:0] phv_data_77; // @[executor.scala 151:22]
  reg [7:0] phv_data_78; // @[executor.scala 151:22]
  reg [7:0] phv_data_79; // @[executor.scala 151:22]
  reg [7:0] phv_data_80; // @[executor.scala 151:22]
  reg [7:0] phv_data_81; // @[executor.scala 151:22]
  reg [7:0] phv_data_82; // @[executor.scala 151:22]
  reg [7:0] phv_data_83; // @[executor.scala 151:22]
  reg [7:0] phv_data_84; // @[executor.scala 151:22]
  reg [7:0] phv_data_85; // @[executor.scala 151:22]
  reg [7:0] phv_data_86; // @[executor.scala 151:22]
  reg [7:0] phv_data_87; // @[executor.scala 151:22]
  reg [7:0] phv_data_88; // @[executor.scala 151:22]
  reg [7:0] phv_data_89; // @[executor.scala 151:22]
  reg [7:0] phv_data_90; // @[executor.scala 151:22]
  reg [7:0] phv_data_91; // @[executor.scala 151:22]
  reg [7:0] phv_data_92; // @[executor.scala 151:22]
  reg [7:0] phv_data_93; // @[executor.scala 151:22]
  reg [7:0] phv_data_94; // @[executor.scala 151:22]
  reg [7:0] phv_data_95; // @[executor.scala 151:22]
  reg [7:0] phv_data_96; // @[executor.scala 151:22]
  reg [7:0] phv_data_97; // @[executor.scala 151:22]
  reg [7:0] phv_data_98; // @[executor.scala 151:22]
  reg [7:0] phv_data_99; // @[executor.scala 151:22]
  reg [7:0] phv_data_100; // @[executor.scala 151:22]
  reg [7:0] phv_data_101; // @[executor.scala 151:22]
  reg [7:0] phv_data_102; // @[executor.scala 151:22]
  reg [7:0] phv_data_103; // @[executor.scala 151:22]
  reg [7:0] phv_data_104; // @[executor.scala 151:22]
  reg [7:0] phv_data_105; // @[executor.scala 151:22]
  reg [7:0] phv_data_106; // @[executor.scala 151:22]
  reg [7:0] phv_data_107; // @[executor.scala 151:22]
  reg [7:0] phv_data_108; // @[executor.scala 151:22]
  reg [7:0] phv_data_109; // @[executor.scala 151:22]
  reg [7:0] phv_data_110; // @[executor.scala 151:22]
  reg [7:0] phv_data_111; // @[executor.scala 151:22]
  reg [7:0] phv_data_112; // @[executor.scala 151:22]
  reg [7:0] phv_data_113; // @[executor.scala 151:22]
  reg [7:0] phv_data_114; // @[executor.scala 151:22]
  reg [7:0] phv_data_115; // @[executor.scala 151:22]
  reg [7:0] phv_data_116; // @[executor.scala 151:22]
  reg [7:0] phv_data_117; // @[executor.scala 151:22]
  reg [7:0] phv_data_118; // @[executor.scala 151:22]
  reg [7:0] phv_data_119; // @[executor.scala 151:22]
  reg [7:0] phv_data_120; // @[executor.scala 151:22]
  reg [7:0] phv_data_121; // @[executor.scala 151:22]
  reg [7:0] phv_data_122; // @[executor.scala 151:22]
  reg [7:0] phv_data_123; // @[executor.scala 151:22]
  reg [7:0] phv_data_124; // @[executor.scala 151:22]
  reg [7:0] phv_data_125; // @[executor.scala 151:22]
  reg [7:0] phv_data_126; // @[executor.scala 151:22]
  reg [7:0] phv_data_127; // @[executor.scala 151:22]
  reg [7:0] phv_data_128; // @[executor.scala 151:22]
  reg [7:0] phv_data_129; // @[executor.scala 151:22]
  reg [7:0] phv_data_130; // @[executor.scala 151:22]
  reg [7:0] phv_data_131; // @[executor.scala 151:22]
  reg [7:0] phv_data_132; // @[executor.scala 151:22]
  reg [7:0] phv_data_133; // @[executor.scala 151:22]
  reg [7:0] phv_data_134; // @[executor.scala 151:22]
  reg [7:0] phv_data_135; // @[executor.scala 151:22]
  reg [7:0] phv_data_136; // @[executor.scala 151:22]
  reg [7:0] phv_data_137; // @[executor.scala 151:22]
  reg [7:0] phv_data_138; // @[executor.scala 151:22]
  reg [7:0] phv_data_139; // @[executor.scala 151:22]
  reg [7:0] phv_data_140; // @[executor.scala 151:22]
  reg [7:0] phv_data_141; // @[executor.scala 151:22]
  reg [7:0] phv_data_142; // @[executor.scala 151:22]
  reg [7:0] phv_data_143; // @[executor.scala 151:22]
  reg [7:0] phv_data_144; // @[executor.scala 151:22]
  reg [7:0] phv_data_145; // @[executor.scala 151:22]
  reg [7:0] phv_data_146; // @[executor.scala 151:22]
  reg [7:0] phv_data_147; // @[executor.scala 151:22]
  reg [7:0] phv_data_148; // @[executor.scala 151:22]
  reg [7:0] phv_data_149; // @[executor.scala 151:22]
  reg [7:0] phv_data_150; // @[executor.scala 151:22]
  reg [7:0] phv_data_151; // @[executor.scala 151:22]
  reg [7:0] phv_data_152; // @[executor.scala 151:22]
  reg [7:0] phv_data_153; // @[executor.scala 151:22]
  reg [7:0] phv_data_154; // @[executor.scala 151:22]
  reg [7:0] phv_data_155; // @[executor.scala 151:22]
  reg [7:0] phv_data_156; // @[executor.scala 151:22]
  reg [7:0] phv_data_157; // @[executor.scala 151:22]
  reg [7:0] phv_data_158; // @[executor.scala 151:22]
  reg [7:0] phv_data_159; // @[executor.scala 151:22]
  reg [7:0] phv_data_160; // @[executor.scala 151:22]
  reg [7:0] phv_data_161; // @[executor.scala 151:22]
  reg [7:0] phv_data_162; // @[executor.scala 151:22]
  reg [7:0] phv_data_163; // @[executor.scala 151:22]
  reg [7:0] phv_data_164; // @[executor.scala 151:22]
  reg [7:0] phv_data_165; // @[executor.scala 151:22]
  reg [7:0] phv_data_166; // @[executor.scala 151:22]
  reg [7:0] phv_data_167; // @[executor.scala 151:22]
  reg [7:0] phv_data_168; // @[executor.scala 151:22]
  reg [7:0] phv_data_169; // @[executor.scala 151:22]
  reg [7:0] phv_data_170; // @[executor.scala 151:22]
  reg [7:0] phv_data_171; // @[executor.scala 151:22]
  reg [7:0] phv_data_172; // @[executor.scala 151:22]
  reg [7:0] phv_data_173; // @[executor.scala 151:22]
  reg [7:0] phv_data_174; // @[executor.scala 151:22]
  reg [7:0] phv_data_175; // @[executor.scala 151:22]
  reg [7:0] phv_data_176; // @[executor.scala 151:22]
  reg [7:0] phv_data_177; // @[executor.scala 151:22]
  reg [7:0] phv_data_178; // @[executor.scala 151:22]
  reg [7:0] phv_data_179; // @[executor.scala 151:22]
  reg [7:0] phv_data_180; // @[executor.scala 151:22]
  reg [7:0] phv_data_181; // @[executor.scala 151:22]
  reg [7:0] phv_data_182; // @[executor.scala 151:22]
  reg [7:0] phv_data_183; // @[executor.scala 151:22]
  reg [7:0] phv_data_184; // @[executor.scala 151:22]
  reg [7:0] phv_data_185; // @[executor.scala 151:22]
  reg [7:0] phv_data_186; // @[executor.scala 151:22]
  reg [7:0] phv_data_187; // @[executor.scala 151:22]
  reg [7:0] phv_data_188; // @[executor.scala 151:22]
  reg [7:0] phv_data_189; // @[executor.scala 151:22]
  reg [7:0] phv_data_190; // @[executor.scala 151:22]
  reg [7:0] phv_data_191; // @[executor.scala 151:22]
  reg [7:0] phv_data_192; // @[executor.scala 151:22]
  reg [7:0] phv_data_193; // @[executor.scala 151:22]
  reg [7:0] phv_data_194; // @[executor.scala 151:22]
  reg [7:0] phv_data_195; // @[executor.scala 151:22]
  reg [7:0] phv_data_196; // @[executor.scala 151:22]
  reg [7:0] phv_data_197; // @[executor.scala 151:22]
  reg [7:0] phv_data_198; // @[executor.scala 151:22]
  reg [7:0] phv_data_199; // @[executor.scala 151:22]
  reg [7:0] phv_data_200; // @[executor.scala 151:22]
  reg [7:0] phv_data_201; // @[executor.scala 151:22]
  reg [7:0] phv_data_202; // @[executor.scala 151:22]
  reg [7:0] phv_data_203; // @[executor.scala 151:22]
  reg [7:0] phv_data_204; // @[executor.scala 151:22]
  reg [7:0] phv_data_205; // @[executor.scala 151:22]
  reg [7:0] phv_data_206; // @[executor.scala 151:22]
  reg [7:0] phv_data_207; // @[executor.scala 151:22]
  reg [7:0] phv_data_208; // @[executor.scala 151:22]
  reg [7:0] phv_data_209; // @[executor.scala 151:22]
  reg [7:0] phv_data_210; // @[executor.scala 151:22]
  reg [7:0] phv_data_211; // @[executor.scala 151:22]
  reg [7:0] phv_data_212; // @[executor.scala 151:22]
  reg [7:0] phv_data_213; // @[executor.scala 151:22]
  reg [7:0] phv_data_214; // @[executor.scala 151:22]
  reg [7:0] phv_data_215; // @[executor.scala 151:22]
  reg [7:0] phv_data_216; // @[executor.scala 151:22]
  reg [7:0] phv_data_217; // @[executor.scala 151:22]
  reg [7:0] phv_data_218; // @[executor.scala 151:22]
  reg [7:0] phv_data_219; // @[executor.scala 151:22]
  reg [7:0] phv_data_220; // @[executor.scala 151:22]
  reg [7:0] phv_data_221; // @[executor.scala 151:22]
  reg [7:0] phv_data_222; // @[executor.scala 151:22]
  reg [7:0] phv_data_223; // @[executor.scala 151:22]
  reg [7:0] phv_data_224; // @[executor.scala 151:22]
  reg [7:0] phv_data_225; // @[executor.scala 151:22]
  reg [7:0] phv_data_226; // @[executor.scala 151:22]
  reg [7:0] phv_data_227; // @[executor.scala 151:22]
  reg [7:0] phv_data_228; // @[executor.scala 151:22]
  reg [7:0] phv_data_229; // @[executor.scala 151:22]
  reg [7:0] phv_data_230; // @[executor.scala 151:22]
  reg [7:0] phv_data_231; // @[executor.scala 151:22]
  reg [7:0] phv_data_232; // @[executor.scala 151:22]
  reg [7:0] phv_data_233; // @[executor.scala 151:22]
  reg [7:0] phv_data_234; // @[executor.scala 151:22]
  reg [7:0] phv_data_235; // @[executor.scala 151:22]
  reg [7:0] phv_data_236; // @[executor.scala 151:22]
  reg [7:0] phv_data_237; // @[executor.scala 151:22]
  reg [7:0] phv_data_238; // @[executor.scala 151:22]
  reg [7:0] phv_data_239; // @[executor.scala 151:22]
  reg [7:0] phv_data_240; // @[executor.scala 151:22]
  reg [7:0] phv_data_241; // @[executor.scala 151:22]
  reg [7:0] phv_data_242; // @[executor.scala 151:22]
  reg [7:0] phv_data_243; // @[executor.scala 151:22]
  reg [7:0] phv_data_244; // @[executor.scala 151:22]
  reg [7:0] phv_data_245; // @[executor.scala 151:22]
  reg [7:0] phv_data_246; // @[executor.scala 151:22]
  reg [7:0] phv_data_247; // @[executor.scala 151:22]
  reg [7:0] phv_data_248; // @[executor.scala 151:22]
  reg [7:0] phv_data_249; // @[executor.scala 151:22]
  reg [7:0] phv_data_250; // @[executor.scala 151:22]
  reg [7:0] phv_data_251; // @[executor.scala 151:22]
  reg [7:0] phv_data_252; // @[executor.scala 151:22]
  reg [7:0] phv_data_253; // @[executor.scala 151:22]
  reg [7:0] phv_data_254; // @[executor.scala 151:22]
  reg [7:0] phv_data_255; // @[executor.scala 151:22]
  reg [7:0] phv_data_256; // @[executor.scala 151:22]
  reg [7:0] phv_data_257; // @[executor.scala 151:22]
  reg [7:0] phv_data_258; // @[executor.scala 151:22]
  reg [7:0] phv_data_259; // @[executor.scala 151:22]
  reg [7:0] phv_data_260; // @[executor.scala 151:22]
  reg [7:0] phv_data_261; // @[executor.scala 151:22]
  reg [7:0] phv_data_262; // @[executor.scala 151:22]
  reg [7:0] phv_data_263; // @[executor.scala 151:22]
  reg [7:0] phv_data_264; // @[executor.scala 151:22]
  reg [7:0] phv_data_265; // @[executor.scala 151:22]
  reg [7:0] phv_data_266; // @[executor.scala 151:22]
  reg [7:0] phv_data_267; // @[executor.scala 151:22]
  reg [7:0] phv_data_268; // @[executor.scala 151:22]
  reg [7:0] phv_data_269; // @[executor.scala 151:22]
  reg [7:0] phv_data_270; // @[executor.scala 151:22]
  reg [7:0] phv_data_271; // @[executor.scala 151:22]
  reg [7:0] phv_data_272; // @[executor.scala 151:22]
  reg [7:0] phv_data_273; // @[executor.scala 151:22]
  reg [7:0] phv_data_274; // @[executor.scala 151:22]
  reg [7:0] phv_data_275; // @[executor.scala 151:22]
  reg [7:0] phv_data_276; // @[executor.scala 151:22]
  reg [7:0] phv_data_277; // @[executor.scala 151:22]
  reg [7:0] phv_data_278; // @[executor.scala 151:22]
  reg [7:0] phv_data_279; // @[executor.scala 151:22]
  reg [7:0] phv_data_280; // @[executor.scala 151:22]
  reg [7:0] phv_data_281; // @[executor.scala 151:22]
  reg [7:0] phv_data_282; // @[executor.scala 151:22]
  reg [7:0] phv_data_283; // @[executor.scala 151:22]
  reg [7:0] phv_data_284; // @[executor.scala 151:22]
  reg [7:0] phv_data_285; // @[executor.scala 151:22]
  reg [7:0] phv_data_286; // @[executor.scala 151:22]
  reg [7:0] phv_data_287; // @[executor.scala 151:22]
  reg [7:0] phv_data_288; // @[executor.scala 151:22]
  reg [7:0] phv_data_289; // @[executor.scala 151:22]
  reg [7:0] phv_data_290; // @[executor.scala 151:22]
  reg [7:0] phv_data_291; // @[executor.scala 151:22]
  reg [7:0] phv_data_292; // @[executor.scala 151:22]
  reg [7:0] phv_data_293; // @[executor.scala 151:22]
  reg [7:0] phv_data_294; // @[executor.scala 151:22]
  reg [7:0] phv_data_295; // @[executor.scala 151:22]
  reg [7:0] phv_data_296; // @[executor.scala 151:22]
  reg [7:0] phv_data_297; // @[executor.scala 151:22]
  reg [7:0] phv_data_298; // @[executor.scala 151:22]
  reg [7:0] phv_data_299; // @[executor.scala 151:22]
  reg [7:0] phv_data_300; // @[executor.scala 151:22]
  reg [7:0] phv_data_301; // @[executor.scala 151:22]
  reg [7:0] phv_data_302; // @[executor.scala 151:22]
  reg [7:0] phv_data_303; // @[executor.scala 151:22]
  reg [7:0] phv_data_304; // @[executor.scala 151:22]
  reg [7:0] phv_data_305; // @[executor.scala 151:22]
  reg [7:0] phv_data_306; // @[executor.scala 151:22]
  reg [7:0] phv_data_307; // @[executor.scala 151:22]
  reg [7:0] phv_data_308; // @[executor.scala 151:22]
  reg [7:0] phv_data_309; // @[executor.scala 151:22]
  reg [7:0] phv_data_310; // @[executor.scala 151:22]
  reg [7:0] phv_data_311; // @[executor.scala 151:22]
  reg [7:0] phv_data_312; // @[executor.scala 151:22]
  reg [7:0] phv_data_313; // @[executor.scala 151:22]
  reg [7:0] phv_data_314; // @[executor.scala 151:22]
  reg [7:0] phv_data_315; // @[executor.scala 151:22]
  reg [7:0] phv_data_316; // @[executor.scala 151:22]
  reg [7:0] phv_data_317; // @[executor.scala 151:22]
  reg [7:0] phv_data_318; // @[executor.scala 151:22]
  reg [7:0] phv_data_319; // @[executor.scala 151:22]
  reg [7:0] phv_data_320; // @[executor.scala 151:22]
  reg [7:0] phv_data_321; // @[executor.scala 151:22]
  reg [7:0] phv_data_322; // @[executor.scala 151:22]
  reg [7:0] phv_data_323; // @[executor.scala 151:22]
  reg [7:0] phv_data_324; // @[executor.scala 151:22]
  reg [7:0] phv_data_325; // @[executor.scala 151:22]
  reg [7:0] phv_data_326; // @[executor.scala 151:22]
  reg [7:0] phv_data_327; // @[executor.scala 151:22]
  reg [7:0] phv_data_328; // @[executor.scala 151:22]
  reg [7:0] phv_data_329; // @[executor.scala 151:22]
  reg [7:0] phv_data_330; // @[executor.scala 151:22]
  reg [7:0] phv_data_331; // @[executor.scala 151:22]
  reg [7:0] phv_data_332; // @[executor.scala 151:22]
  reg [7:0] phv_data_333; // @[executor.scala 151:22]
  reg [7:0] phv_data_334; // @[executor.scala 151:22]
  reg [7:0] phv_data_335; // @[executor.scala 151:22]
  reg [7:0] phv_data_336; // @[executor.scala 151:22]
  reg [7:0] phv_data_337; // @[executor.scala 151:22]
  reg [7:0] phv_data_338; // @[executor.scala 151:22]
  reg [7:0] phv_data_339; // @[executor.scala 151:22]
  reg [7:0] phv_data_340; // @[executor.scala 151:22]
  reg [7:0] phv_data_341; // @[executor.scala 151:22]
  reg [7:0] phv_data_342; // @[executor.scala 151:22]
  reg [7:0] phv_data_343; // @[executor.scala 151:22]
  reg [7:0] phv_data_344; // @[executor.scala 151:22]
  reg [7:0] phv_data_345; // @[executor.scala 151:22]
  reg [7:0] phv_data_346; // @[executor.scala 151:22]
  reg [7:0] phv_data_347; // @[executor.scala 151:22]
  reg [7:0] phv_data_348; // @[executor.scala 151:22]
  reg [7:0] phv_data_349; // @[executor.scala 151:22]
  reg [7:0] phv_data_350; // @[executor.scala 151:22]
  reg [7:0] phv_data_351; // @[executor.scala 151:22]
  reg [7:0] phv_data_352; // @[executor.scala 151:22]
  reg [7:0] phv_data_353; // @[executor.scala 151:22]
  reg [7:0] phv_data_354; // @[executor.scala 151:22]
  reg [7:0] phv_data_355; // @[executor.scala 151:22]
  reg [7:0] phv_data_356; // @[executor.scala 151:22]
  reg [7:0] phv_data_357; // @[executor.scala 151:22]
  reg [7:0] phv_data_358; // @[executor.scala 151:22]
  reg [7:0] phv_data_359; // @[executor.scala 151:22]
  reg [7:0] phv_data_360; // @[executor.scala 151:22]
  reg [7:0] phv_data_361; // @[executor.scala 151:22]
  reg [7:0] phv_data_362; // @[executor.scala 151:22]
  reg [7:0] phv_data_363; // @[executor.scala 151:22]
  reg [7:0] phv_data_364; // @[executor.scala 151:22]
  reg [7:0] phv_data_365; // @[executor.scala 151:22]
  reg [7:0] phv_data_366; // @[executor.scala 151:22]
  reg [7:0] phv_data_367; // @[executor.scala 151:22]
  reg [7:0] phv_data_368; // @[executor.scala 151:22]
  reg [7:0] phv_data_369; // @[executor.scala 151:22]
  reg [7:0] phv_data_370; // @[executor.scala 151:22]
  reg [7:0] phv_data_371; // @[executor.scala 151:22]
  reg [7:0] phv_data_372; // @[executor.scala 151:22]
  reg [7:0] phv_data_373; // @[executor.scala 151:22]
  reg [7:0] phv_data_374; // @[executor.scala 151:22]
  reg [7:0] phv_data_375; // @[executor.scala 151:22]
  reg [7:0] phv_data_376; // @[executor.scala 151:22]
  reg [7:0] phv_data_377; // @[executor.scala 151:22]
  reg [7:0] phv_data_378; // @[executor.scala 151:22]
  reg [7:0] phv_data_379; // @[executor.scala 151:22]
  reg [7:0] phv_data_380; // @[executor.scala 151:22]
  reg [7:0] phv_data_381; // @[executor.scala 151:22]
  reg [7:0] phv_data_382; // @[executor.scala 151:22]
  reg [7:0] phv_data_383; // @[executor.scala 151:22]
  reg [7:0] phv_data_384; // @[executor.scala 151:22]
  reg [7:0] phv_data_385; // @[executor.scala 151:22]
  reg [7:0] phv_data_386; // @[executor.scala 151:22]
  reg [7:0] phv_data_387; // @[executor.scala 151:22]
  reg [7:0] phv_data_388; // @[executor.scala 151:22]
  reg [7:0] phv_data_389; // @[executor.scala 151:22]
  reg [7:0] phv_data_390; // @[executor.scala 151:22]
  reg [7:0] phv_data_391; // @[executor.scala 151:22]
  reg [7:0] phv_data_392; // @[executor.scala 151:22]
  reg [7:0] phv_data_393; // @[executor.scala 151:22]
  reg [7:0] phv_data_394; // @[executor.scala 151:22]
  reg [7:0] phv_data_395; // @[executor.scala 151:22]
  reg [7:0] phv_data_396; // @[executor.scala 151:22]
  reg [7:0] phv_data_397; // @[executor.scala 151:22]
  reg [7:0] phv_data_398; // @[executor.scala 151:22]
  reg [7:0] phv_data_399; // @[executor.scala 151:22]
  reg [7:0] phv_data_400; // @[executor.scala 151:22]
  reg [7:0] phv_data_401; // @[executor.scala 151:22]
  reg [7:0] phv_data_402; // @[executor.scala 151:22]
  reg [7:0] phv_data_403; // @[executor.scala 151:22]
  reg [7:0] phv_data_404; // @[executor.scala 151:22]
  reg [7:0] phv_data_405; // @[executor.scala 151:22]
  reg [7:0] phv_data_406; // @[executor.scala 151:22]
  reg [7:0] phv_data_407; // @[executor.scala 151:22]
  reg [7:0] phv_data_408; // @[executor.scala 151:22]
  reg [7:0] phv_data_409; // @[executor.scala 151:22]
  reg [7:0] phv_data_410; // @[executor.scala 151:22]
  reg [7:0] phv_data_411; // @[executor.scala 151:22]
  reg [7:0] phv_data_412; // @[executor.scala 151:22]
  reg [7:0] phv_data_413; // @[executor.scala 151:22]
  reg [7:0] phv_data_414; // @[executor.scala 151:22]
  reg [7:0] phv_data_415; // @[executor.scala 151:22]
  reg [7:0] phv_data_416; // @[executor.scala 151:22]
  reg [7:0] phv_data_417; // @[executor.scala 151:22]
  reg [7:0] phv_data_418; // @[executor.scala 151:22]
  reg [7:0] phv_data_419; // @[executor.scala 151:22]
  reg [7:0] phv_data_420; // @[executor.scala 151:22]
  reg [7:0] phv_data_421; // @[executor.scala 151:22]
  reg [7:0] phv_data_422; // @[executor.scala 151:22]
  reg [7:0] phv_data_423; // @[executor.scala 151:22]
  reg [7:0] phv_data_424; // @[executor.scala 151:22]
  reg [7:0] phv_data_425; // @[executor.scala 151:22]
  reg [7:0] phv_data_426; // @[executor.scala 151:22]
  reg [7:0] phv_data_427; // @[executor.scala 151:22]
  reg [7:0] phv_data_428; // @[executor.scala 151:22]
  reg [7:0] phv_data_429; // @[executor.scala 151:22]
  reg [7:0] phv_data_430; // @[executor.scala 151:22]
  reg [7:0] phv_data_431; // @[executor.scala 151:22]
  reg [7:0] phv_data_432; // @[executor.scala 151:22]
  reg [7:0] phv_data_433; // @[executor.scala 151:22]
  reg [7:0] phv_data_434; // @[executor.scala 151:22]
  reg [7:0] phv_data_435; // @[executor.scala 151:22]
  reg [7:0] phv_data_436; // @[executor.scala 151:22]
  reg [7:0] phv_data_437; // @[executor.scala 151:22]
  reg [7:0] phv_data_438; // @[executor.scala 151:22]
  reg [7:0] phv_data_439; // @[executor.scala 151:22]
  reg [7:0] phv_data_440; // @[executor.scala 151:22]
  reg [7:0] phv_data_441; // @[executor.scala 151:22]
  reg [7:0] phv_data_442; // @[executor.scala 151:22]
  reg [7:0] phv_data_443; // @[executor.scala 151:22]
  reg [7:0] phv_data_444; // @[executor.scala 151:22]
  reg [7:0] phv_data_445; // @[executor.scala 151:22]
  reg [7:0] phv_data_446; // @[executor.scala 151:22]
  reg [7:0] phv_data_447; // @[executor.scala 151:22]
  reg [7:0] phv_data_448; // @[executor.scala 151:22]
  reg [7:0] phv_data_449; // @[executor.scala 151:22]
  reg [7:0] phv_data_450; // @[executor.scala 151:22]
  reg [7:0] phv_data_451; // @[executor.scala 151:22]
  reg [7:0] phv_data_452; // @[executor.scala 151:22]
  reg [7:0] phv_data_453; // @[executor.scala 151:22]
  reg [7:0] phv_data_454; // @[executor.scala 151:22]
  reg [7:0] phv_data_455; // @[executor.scala 151:22]
  reg [7:0] phv_data_456; // @[executor.scala 151:22]
  reg [7:0] phv_data_457; // @[executor.scala 151:22]
  reg [7:0] phv_data_458; // @[executor.scala 151:22]
  reg [7:0] phv_data_459; // @[executor.scala 151:22]
  reg [7:0] phv_data_460; // @[executor.scala 151:22]
  reg [7:0] phv_data_461; // @[executor.scala 151:22]
  reg [7:0] phv_data_462; // @[executor.scala 151:22]
  reg [7:0] phv_data_463; // @[executor.scala 151:22]
  reg [7:0] phv_data_464; // @[executor.scala 151:22]
  reg [7:0] phv_data_465; // @[executor.scala 151:22]
  reg [7:0] phv_data_466; // @[executor.scala 151:22]
  reg [7:0] phv_data_467; // @[executor.scala 151:22]
  reg [7:0] phv_data_468; // @[executor.scala 151:22]
  reg [7:0] phv_data_469; // @[executor.scala 151:22]
  reg [7:0] phv_data_470; // @[executor.scala 151:22]
  reg [7:0] phv_data_471; // @[executor.scala 151:22]
  reg [7:0] phv_data_472; // @[executor.scala 151:22]
  reg [7:0] phv_data_473; // @[executor.scala 151:22]
  reg [7:0] phv_data_474; // @[executor.scala 151:22]
  reg [7:0] phv_data_475; // @[executor.scala 151:22]
  reg [7:0] phv_data_476; // @[executor.scala 151:22]
  reg [7:0] phv_data_477; // @[executor.scala 151:22]
  reg [7:0] phv_data_478; // @[executor.scala 151:22]
  reg [7:0] phv_data_479; // @[executor.scala 151:22]
  reg [7:0] phv_data_480; // @[executor.scala 151:22]
  reg [7:0] phv_data_481; // @[executor.scala 151:22]
  reg [7:0] phv_data_482; // @[executor.scala 151:22]
  reg [7:0] phv_data_483; // @[executor.scala 151:22]
  reg [7:0] phv_data_484; // @[executor.scala 151:22]
  reg [7:0] phv_data_485; // @[executor.scala 151:22]
  reg [7:0] phv_data_486; // @[executor.scala 151:22]
  reg [7:0] phv_data_487; // @[executor.scala 151:22]
  reg [7:0] phv_data_488; // @[executor.scala 151:22]
  reg [7:0] phv_data_489; // @[executor.scala 151:22]
  reg [7:0] phv_data_490; // @[executor.scala 151:22]
  reg [7:0] phv_data_491; // @[executor.scala 151:22]
  reg [7:0] phv_data_492; // @[executor.scala 151:22]
  reg [7:0] phv_data_493; // @[executor.scala 151:22]
  reg [7:0] phv_data_494; // @[executor.scala 151:22]
  reg [7:0] phv_data_495; // @[executor.scala 151:22]
  reg [7:0] phv_data_496; // @[executor.scala 151:22]
  reg [7:0] phv_data_497; // @[executor.scala 151:22]
  reg [7:0] phv_data_498; // @[executor.scala 151:22]
  reg [7:0] phv_data_499; // @[executor.scala 151:22]
  reg [7:0] phv_data_500; // @[executor.scala 151:22]
  reg [7:0] phv_data_501; // @[executor.scala 151:22]
  reg [7:0] phv_data_502; // @[executor.scala 151:22]
  reg [7:0] phv_data_503; // @[executor.scala 151:22]
  reg [7:0] phv_data_504; // @[executor.scala 151:22]
  reg [7:0] phv_data_505; // @[executor.scala 151:22]
  reg [7:0] phv_data_506; // @[executor.scala 151:22]
  reg [7:0] phv_data_507; // @[executor.scala 151:22]
  reg [7:0] phv_data_508; // @[executor.scala 151:22]
  reg [7:0] phv_data_509; // @[executor.scala 151:22]
  reg [7:0] phv_data_510; // @[executor.scala 151:22]
  reg [7:0] phv_data_511; // @[executor.scala 151:22]
  reg [15:0] phv_header_0; // @[executor.scala 151:22]
  reg [15:0] phv_header_1; // @[executor.scala 151:22]
  reg [15:0] phv_header_2; // @[executor.scala 151:22]
  reg [15:0] phv_header_3; // @[executor.scala 151:22]
  reg [15:0] phv_header_4; // @[executor.scala 151:22]
  reg [15:0] phv_header_5; // @[executor.scala 151:22]
  reg [15:0] phv_header_6; // @[executor.scala 151:22]
  reg [15:0] phv_header_7; // @[executor.scala 151:22]
  reg [15:0] phv_header_8; // @[executor.scala 151:22]
  reg [15:0] phv_header_9; // @[executor.scala 151:22]
  reg [15:0] phv_header_10; // @[executor.scala 151:22]
  reg [15:0] phv_header_11; // @[executor.scala 151:22]
  reg [15:0] phv_header_12; // @[executor.scala 151:22]
  reg [15:0] phv_header_13; // @[executor.scala 151:22]
  reg [15:0] phv_header_14; // @[executor.scala 151:22]
  reg [15:0] phv_header_15; // @[executor.scala 151:22]
  reg [7:0] phv_parse_current_state; // @[executor.scala 151:22]
  reg [7:0] phv_parse_current_offset; // @[executor.scala 151:22]
  reg [15:0] phv_parse_transition_field; // @[executor.scala 151:22]
  reg [3:0] phv_next_processor_id; // @[executor.scala 151:22]
  reg  phv_next_config_id; // @[executor.scala 151:22]
  reg  phv_is_valid_processor; // @[executor.scala 151:22]
  reg [7:0] args_0; // @[executor.scala 155:23]
  reg [7:0] args_1; // @[executor.scala 155:23]
  reg [7:0] args_2; // @[executor.scala 155:23]
  reg [7:0] args_3; // @[executor.scala 155:23]
  reg [7:0] args_4; // @[executor.scala 155:23]
  reg [7:0] args_5; // @[executor.scala 155:23]
  reg [7:0] args_6; // @[executor.scala 155:23]
  reg [31:0] vliw_0; // @[executor.scala 158:23]
  reg [31:0] vliw_1; // @[executor.scala 158:23]
  reg [31:0] vliw_2; // @[executor.scala 158:23]
  reg [31:0] vliw_3; // @[executor.scala 158:23]
  reg [7:0] offset_0; // @[executor.scala 162:25]
  reg [7:0] offset_1; // @[executor.scala 162:25]
  reg [7:0] offset_2; // @[executor.scala 162:25]
  reg [7:0] offset_3; // @[executor.scala 162:25]
  reg [7:0] length_0; // @[executor.scala 163:25]
  reg [7:0] length_1; // @[executor.scala 163:25]
  reg [7:0] length_2; // @[executor.scala 163:25]
  reg [7:0] length_3; // @[executor.scala 163:25]
  wire [3:0] opcode = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_0_lo = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire  from_header = length_0 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi = offset_0[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_1 = offset_0 + length_0; // @[executor.scala 193:46]
  wire [1:0] ending = _ending_T_1[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_9120 = {{2'd0}, ending}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_1 = 4'h4 - _GEN_9120; // @[executor.scala 194:45]
  wire [1:0] bias = _bias_T_1[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset = {total_offset_hi,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1 = 8'h1 == total_offset ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2 = 8'h2 == total_offset ? phv_data_2 : _GEN_1; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3 = 8'h3 == total_offset ? phv_data_3 : _GEN_2; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4 = 8'h4 == total_offset ? phv_data_4 : _GEN_3; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5 = 8'h5 == total_offset ? phv_data_5 : _GEN_4; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6 = 8'h6 == total_offset ? phv_data_6 : _GEN_5; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7 = 8'h7 == total_offset ? phv_data_7 : _GEN_6; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8 = 8'h8 == total_offset ? phv_data_8 : _GEN_7; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_9 = 8'h9 == total_offset ? phv_data_9 : _GEN_8; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_10 = 8'ha == total_offset ? phv_data_10 : _GEN_9; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_11 = 8'hb == total_offset ? phv_data_11 : _GEN_10; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_12 = 8'hc == total_offset ? phv_data_12 : _GEN_11; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_13 = 8'hd == total_offset ? phv_data_13 : _GEN_12; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_14 = 8'he == total_offset ? phv_data_14 : _GEN_13; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_15 = 8'hf == total_offset ? phv_data_15 : _GEN_14; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_16 = 8'h10 == total_offset ? phv_data_16 : _GEN_15; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_17 = 8'h11 == total_offset ? phv_data_17 : _GEN_16; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_18 = 8'h12 == total_offset ? phv_data_18 : _GEN_17; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_19 = 8'h13 == total_offset ? phv_data_19 : _GEN_18; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_20 = 8'h14 == total_offset ? phv_data_20 : _GEN_19; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_21 = 8'h15 == total_offset ? phv_data_21 : _GEN_20; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_22 = 8'h16 == total_offset ? phv_data_22 : _GEN_21; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_23 = 8'h17 == total_offset ? phv_data_23 : _GEN_22; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_24 = 8'h18 == total_offset ? phv_data_24 : _GEN_23; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_25 = 8'h19 == total_offset ? phv_data_25 : _GEN_24; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_26 = 8'h1a == total_offset ? phv_data_26 : _GEN_25; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_27 = 8'h1b == total_offset ? phv_data_27 : _GEN_26; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_28 = 8'h1c == total_offset ? phv_data_28 : _GEN_27; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_29 = 8'h1d == total_offset ? phv_data_29 : _GEN_28; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_30 = 8'h1e == total_offset ? phv_data_30 : _GEN_29; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_31 = 8'h1f == total_offset ? phv_data_31 : _GEN_30; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_32 = 8'h20 == total_offset ? phv_data_32 : _GEN_31; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_33 = 8'h21 == total_offset ? phv_data_33 : _GEN_32; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_34 = 8'h22 == total_offset ? phv_data_34 : _GEN_33; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_35 = 8'h23 == total_offset ? phv_data_35 : _GEN_34; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_36 = 8'h24 == total_offset ? phv_data_36 : _GEN_35; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_37 = 8'h25 == total_offset ? phv_data_37 : _GEN_36; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_38 = 8'h26 == total_offset ? phv_data_38 : _GEN_37; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_39 = 8'h27 == total_offset ? phv_data_39 : _GEN_38; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_40 = 8'h28 == total_offset ? phv_data_40 : _GEN_39; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_41 = 8'h29 == total_offset ? phv_data_41 : _GEN_40; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_42 = 8'h2a == total_offset ? phv_data_42 : _GEN_41; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_43 = 8'h2b == total_offset ? phv_data_43 : _GEN_42; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_44 = 8'h2c == total_offset ? phv_data_44 : _GEN_43; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_45 = 8'h2d == total_offset ? phv_data_45 : _GEN_44; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_46 = 8'h2e == total_offset ? phv_data_46 : _GEN_45; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_47 = 8'h2f == total_offset ? phv_data_47 : _GEN_46; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_48 = 8'h30 == total_offset ? phv_data_48 : _GEN_47; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_49 = 8'h31 == total_offset ? phv_data_49 : _GEN_48; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_50 = 8'h32 == total_offset ? phv_data_50 : _GEN_49; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_51 = 8'h33 == total_offset ? phv_data_51 : _GEN_50; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_52 = 8'h34 == total_offset ? phv_data_52 : _GEN_51; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_53 = 8'h35 == total_offset ? phv_data_53 : _GEN_52; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_54 = 8'h36 == total_offset ? phv_data_54 : _GEN_53; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_55 = 8'h37 == total_offset ? phv_data_55 : _GEN_54; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_56 = 8'h38 == total_offset ? phv_data_56 : _GEN_55; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_57 = 8'h39 == total_offset ? phv_data_57 : _GEN_56; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_58 = 8'h3a == total_offset ? phv_data_58 : _GEN_57; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_59 = 8'h3b == total_offset ? phv_data_59 : _GEN_58; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_60 = 8'h3c == total_offset ? phv_data_60 : _GEN_59; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_61 = 8'h3d == total_offset ? phv_data_61 : _GEN_60; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_62 = 8'h3e == total_offset ? phv_data_62 : _GEN_61; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_63 = 8'h3f == total_offset ? phv_data_63 : _GEN_62; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_64 = 8'h40 == total_offset ? phv_data_64 : _GEN_63; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_65 = 8'h41 == total_offset ? phv_data_65 : _GEN_64; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_66 = 8'h42 == total_offset ? phv_data_66 : _GEN_65; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_67 = 8'h43 == total_offset ? phv_data_67 : _GEN_66; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_68 = 8'h44 == total_offset ? phv_data_68 : _GEN_67; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_69 = 8'h45 == total_offset ? phv_data_69 : _GEN_68; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_70 = 8'h46 == total_offset ? phv_data_70 : _GEN_69; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_71 = 8'h47 == total_offset ? phv_data_71 : _GEN_70; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_72 = 8'h48 == total_offset ? phv_data_72 : _GEN_71; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_73 = 8'h49 == total_offset ? phv_data_73 : _GEN_72; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_74 = 8'h4a == total_offset ? phv_data_74 : _GEN_73; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_75 = 8'h4b == total_offset ? phv_data_75 : _GEN_74; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_76 = 8'h4c == total_offset ? phv_data_76 : _GEN_75; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_77 = 8'h4d == total_offset ? phv_data_77 : _GEN_76; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_78 = 8'h4e == total_offset ? phv_data_78 : _GEN_77; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_79 = 8'h4f == total_offset ? phv_data_79 : _GEN_78; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_80 = 8'h50 == total_offset ? phv_data_80 : _GEN_79; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_81 = 8'h51 == total_offset ? phv_data_81 : _GEN_80; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_82 = 8'h52 == total_offset ? phv_data_82 : _GEN_81; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_83 = 8'h53 == total_offset ? phv_data_83 : _GEN_82; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_84 = 8'h54 == total_offset ? phv_data_84 : _GEN_83; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_85 = 8'h55 == total_offset ? phv_data_85 : _GEN_84; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_86 = 8'h56 == total_offset ? phv_data_86 : _GEN_85; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_87 = 8'h57 == total_offset ? phv_data_87 : _GEN_86; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_88 = 8'h58 == total_offset ? phv_data_88 : _GEN_87; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_89 = 8'h59 == total_offset ? phv_data_89 : _GEN_88; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_90 = 8'h5a == total_offset ? phv_data_90 : _GEN_89; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_91 = 8'h5b == total_offset ? phv_data_91 : _GEN_90; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_92 = 8'h5c == total_offset ? phv_data_92 : _GEN_91; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_93 = 8'h5d == total_offset ? phv_data_93 : _GEN_92; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_94 = 8'h5e == total_offset ? phv_data_94 : _GEN_93; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_95 = 8'h5f == total_offset ? phv_data_95 : _GEN_94; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_96 = 8'h60 == total_offset ? phv_data_96 : _GEN_95; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_97 = 8'h61 == total_offset ? phv_data_97 : _GEN_96; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_98 = 8'h62 == total_offset ? phv_data_98 : _GEN_97; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_99 = 8'h63 == total_offset ? phv_data_99 : _GEN_98; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_100 = 8'h64 == total_offset ? phv_data_100 : _GEN_99; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_101 = 8'h65 == total_offset ? phv_data_101 : _GEN_100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_102 = 8'h66 == total_offset ? phv_data_102 : _GEN_101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_103 = 8'h67 == total_offset ? phv_data_103 : _GEN_102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_104 = 8'h68 == total_offset ? phv_data_104 : _GEN_103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_105 = 8'h69 == total_offset ? phv_data_105 : _GEN_104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_106 = 8'h6a == total_offset ? phv_data_106 : _GEN_105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_107 = 8'h6b == total_offset ? phv_data_107 : _GEN_106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_108 = 8'h6c == total_offset ? phv_data_108 : _GEN_107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_109 = 8'h6d == total_offset ? phv_data_109 : _GEN_108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_110 = 8'h6e == total_offset ? phv_data_110 : _GEN_109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_111 = 8'h6f == total_offset ? phv_data_111 : _GEN_110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_112 = 8'h70 == total_offset ? phv_data_112 : _GEN_111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_113 = 8'h71 == total_offset ? phv_data_113 : _GEN_112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_114 = 8'h72 == total_offset ? phv_data_114 : _GEN_113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_115 = 8'h73 == total_offset ? phv_data_115 : _GEN_114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_116 = 8'h74 == total_offset ? phv_data_116 : _GEN_115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_117 = 8'h75 == total_offset ? phv_data_117 : _GEN_116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_118 = 8'h76 == total_offset ? phv_data_118 : _GEN_117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_119 = 8'h77 == total_offset ? phv_data_119 : _GEN_118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_120 = 8'h78 == total_offset ? phv_data_120 : _GEN_119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_121 = 8'h79 == total_offset ? phv_data_121 : _GEN_120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_122 = 8'h7a == total_offset ? phv_data_122 : _GEN_121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_123 = 8'h7b == total_offset ? phv_data_123 : _GEN_122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_124 = 8'h7c == total_offset ? phv_data_124 : _GEN_123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_125 = 8'h7d == total_offset ? phv_data_125 : _GEN_124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_126 = 8'h7e == total_offset ? phv_data_126 : _GEN_125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_127 = 8'h7f == total_offset ? phv_data_127 : _GEN_126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_128 = 8'h80 == total_offset ? phv_data_128 : _GEN_127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_129 = 8'h81 == total_offset ? phv_data_129 : _GEN_128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_130 = 8'h82 == total_offset ? phv_data_130 : _GEN_129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_131 = 8'h83 == total_offset ? phv_data_131 : _GEN_130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_132 = 8'h84 == total_offset ? phv_data_132 : _GEN_131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_133 = 8'h85 == total_offset ? phv_data_133 : _GEN_132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_134 = 8'h86 == total_offset ? phv_data_134 : _GEN_133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_135 = 8'h87 == total_offset ? phv_data_135 : _GEN_134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_136 = 8'h88 == total_offset ? phv_data_136 : _GEN_135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_137 = 8'h89 == total_offset ? phv_data_137 : _GEN_136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_138 = 8'h8a == total_offset ? phv_data_138 : _GEN_137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_139 = 8'h8b == total_offset ? phv_data_139 : _GEN_138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_140 = 8'h8c == total_offset ? phv_data_140 : _GEN_139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_141 = 8'h8d == total_offset ? phv_data_141 : _GEN_140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_142 = 8'h8e == total_offset ? phv_data_142 : _GEN_141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_143 = 8'h8f == total_offset ? phv_data_143 : _GEN_142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_144 = 8'h90 == total_offset ? phv_data_144 : _GEN_143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_145 = 8'h91 == total_offset ? phv_data_145 : _GEN_144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_146 = 8'h92 == total_offset ? phv_data_146 : _GEN_145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_147 = 8'h93 == total_offset ? phv_data_147 : _GEN_146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_148 = 8'h94 == total_offset ? phv_data_148 : _GEN_147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_149 = 8'h95 == total_offset ? phv_data_149 : _GEN_148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_150 = 8'h96 == total_offset ? phv_data_150 : _GEN_149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_151 = 8'h97 == total_offset ? phv_data_151 : _GEN_150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_152 = 8'h98 == total_offset ? phv_data_152 : _GEN_151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_153 = 8'h99 == total_offset ? phv_data_153 : _GEN_152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_154 = 8'h9a == total_offset ? phv_data_154 : _GEN_153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_155 = 8'h9b == total_offset ? phv_data_155 : _GEN_154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_156 = 8'h9c == total_offset ? phv_data_156 : _GEN_155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_157 = 8'h9d == total_offset ? phv_data_157 : _GEN_156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_158 = 8'h9e == total_offset ? phv_data_158 : _GEN_157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_159 = 8'h9f == total_offset ? phv_data_159 : _GEN_158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_160 = 8'ha0 == total_offset ? phv_data_160 : _GEN_159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_161 = 8'ha1 == total_offset ? phv_data_161 : _GEN_160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_162 = 8'ha2 == total_offset ? phv_data_162 : _GEN_161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_163 = 8'ha3 == total_offset ? phv_data_163 : _GEN_162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_164 = 8'ha4 == total_offset ? phv_data_164 : _GEN_163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_165 = 8'ha5 == total_offset ? phv_data_165 : _GEN_164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_166 = 8'ha6 == total_offset ? phv_data_166 : _GEN_165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_167 = 8'ha7 == total_offset ? phv_data_167 : _GEN_166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_168 = 8'ha8 == total_offset ? phv_data_168 : _GEN_167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_169 = 8'ha9 == total_offset ? phv_data_169 : _GEN_168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_170 = 8'haa == total_offset ? phv_data_170 : _GEN_169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_171 = 8'hab == total_offset ? phv_data_171 : _GEN_170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_172 = 8'hac == total_offset ? phv_data_172 : _GEN_171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_173 = 8'had == total_offset ? phv_data_173 : _GEN_172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_174 = 8'hae == total_offset ? phv_data_174 : _GEN_173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_175 = 8'haf == total_offset ? phv_data_175 : _GEN_174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_176 = 8'hb0 == total_offset ? phv_data_176 : _GEN_175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_177 = 8'hb1 == total_offset ? phv_data_177 : _GEN_176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_178 = 8'hb2 == total_offset ? phv_data_178 : _GEN_177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_179 = 8'hb3 == total_offset ? phv_data_179 : _GEN_178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_180 = 8'hb4 == total_offset ? phv_data_180 : _GEN_179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_181 = 8'hb5 == total_offset ? phv_data_181 : _GEN_180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_182 = 8'hb6 == total_offset ? phv_data_182 : _GEN_181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_183 = 8'hb7 == total_offset ? phv_data_183 : _GEN_182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_184 = 8'hb8 == total_offset ? phv_data_184 : _GEN_183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_185 = 8'hb9 == total_offset ? phv_data_185 : _GEN_184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_186 = 8'hba == total_offset ? phv_data_186 : _GEN_185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_187 = 8'hbb == total_offset ? phv_data_187 : _GEN_186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_188 = 8'hbc == total_offset ? phv_data_188 : _GEN_187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_189 = 8'hbd == total_offset ? phv_data_189 : _GEN_188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_190 = 8'hbe == total_offset ? phv_data_190 : _GEN_189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_191 = 8'hbf == total_offset ? phv_data_191 : _GEN_190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_192 = 8'hc0 == total_offset ? phv_data_192 : _GEN_191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_193 = 8'hc1 == total_offset ? phv_data_193 : _GEN_192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_194 = 8'hc2 == total_offset ? phv_data_194 : _GEN_193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_195 = 8'hc3 == total_offset ? phv_data_195 : _GEN_194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_196 = 8'hc4 == total_offset ? phv_data_196 : _GEN_195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_197 = 8'hc5 == total_offset ? phv_data_197 : _GEN_196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_198 = 8'hc6 == total_offset ? phv_data_198 : _GEN_197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_199 = 8'hc7 == total_offset ? phv_data_199 : _GEN_198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_200 = 8'hc8 == total_offset ? phv_data_200 : _GEN_199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_201 = 8'hc9 == total_offset ? phv_data_201 : _GEN_200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_202 = 8'hca == total_offset ? phv_data_202 : _GEN_201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_203 = 8'hcb == total_offset ? phv_data_203 : _GEN_202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_204 = 8'hcc == total_offset ? phv_data_204 : _GEN_203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_205 = 8'hcd == total_offset ? phv_data_205 : _GEN_204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_206 = 8'hce == total_offset ? phv_data_206 : _GEN_205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_207 = 8'hcf == total_offset ? phv_data_207 : _GEN_206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_208 = 8'hd0 == total_offset ? phv_data_208 : _GEN_207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_209 = 8'hd1 == total_offset ? phv_data_209 : _GEN_208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_210 = 8'hd2 == total_offset ? phv_data_210 : _GEN_209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_211 = 8'hd3 == total_offset ? phv_data_211 : _GEN_210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_212 = 8'hd4 == total_offset ? phv_data_212 : _GEN_211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_213 = 8'hd5 == total_offset ? phv_data_213 : _GEN_212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_214 = 8'hd6 == total_offset ? phv_data_214 : _GEN_213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_215 = 8'hd7 == total_offset ? phv_data_215 : _GEN_214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_216 = 8'hd8 == total_offset ? phv_data_216 : _GEN_215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_217 = 8'hd9 == total_offset ? phv_data_217 : _GEN_216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_218 = 8'hda == total_offset ? phv_data_218 : _GEN_217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_219 = 8'hdb == total_offset ? phv_data_219 : _GEN_218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_220 = 8'hdc == total_offset ? phv_data_220 : _GEN_219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_221 = 8'hdd == total_offset ? phv_data_221 : _GEN_220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_222 = 8'hde == total_offset ? phv_data_222 : _GEN_221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_223 = 8'hdf == total_offset ? phv_data_223 : _GEN_222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_224 = 8'he0 == total_offset ? phv_data_224 : _GEN_223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_225 = 8'he1 == total_offset ? phv_data_225 : _GEN_224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_226 = 8'he2 == total_offset ? phv_data_226 : _GEN_225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_227 = 8'he3 == total_offset ? phv_data_227 : _GEN_226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_228 = 8'he4 == total_offset ? phv_data_228 : _GEN_227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_229 = 8'he5 == total_offset ? phv_data_229 : _GEN_228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_230 = 8'he6 == total_offset ? phv_data_230 : _GEN_229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_231 = 8'he7 == total_offset ? phv_data_231 : _GEN_230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_232 = 8'he8 == total_offset ? phv_data_232 : _GEN_231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_233 = 8'he9 == total_offset ? phv_data_233 : _GEN_232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_234 = 8'hea == total_offset ? phv_data_234 : _GEN_233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_235 = 8'heb == total_offset ? phv_data_235 : _GEN_234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_236 = 8'hec == total_offset ? phv_data_236 : _GEN_235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_237 = 8'hed == total_offset ? phv_data_237 : _GEN_236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_238 = 8'hee == total_offset ? phv_data_238 : _GEN_237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_239 = 8'hef == total_offset ? phv_data_239 : _GEN_238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_240 = 8'hf0 == total_offset ? phv_data_240 : _GEN_239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_241 = 8'hf1 == total_offset ? phv_data_241 : _GEN_240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_242 = 8'hf2 == total_offset ? phv_data_242 : _GEN_241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_243 = 8'hf3 == total_offset ? phv_data_243 : _GEN_242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_244 = 8'hf4 == total_offset ? phv_data_244 : _GEN_243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_245 = 8'hf5 == total_offset ? phv_data_245 : _GEN_244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_246 = 8'hf6 == total_offset ? phv_data_246 : _GEN_245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_247 = 8'hf7 == total_offset ? phv_data_247 : _GEN_246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_248 = 8'hf8 == total_offset ? phv_data_248 : _GEN_247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_249 = 8'hf9 == total_offset ? phv_data_249 : _GEN_248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_250 = 8'hfa == total_offset ? phv_data_250 : _GEN_249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_251 = 8'hfb == total_offset ? phv_data_251 : _GEN_250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_252 = 8'hfc == total_offset ? phv_data_252 : _GEN_251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_253 = 8'hfd == total_offset ? phv_data_253 : _GEN_252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_254 = 8'hfe == total_offset ? phv_data_254 : _GEN_253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_255 = 8'hff == total_offset ? phv_data_255 : _GEN_254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_9121 = {{1'd0}, total_offset}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_256 = 9'h100 == _GEN_9121 ? phv_data_256 : _GEN_255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_257 = 9'h101 == _GEN_9121 ? phv_data_257 : _GEN_256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_258 = 9'h102 == _GEN_9121 ? phv_data_258 : _GEN_257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_259 = 9'h103 == _GEN_9121 ? phv_data_259 : _GEN_258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_260 = 9'h104 == _GEN_9121 ? phv_data_260 : _GEN_259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_261 = 9'h105 == _GEN_9121 ? phv_data_261 : _GEN_260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_262 = 9'h106 == _GEN_9121 ? phv_data_262 : _GEN_261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_263 = 9'h107 == _GEN_9121 ? phv_data_263 : _GEN_262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_264 = 9'h108 == _GEN_9121 ? phv_data_264 : _GEN_263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_265 = 9'h109 == _GEN_9121 ? phv_data_265 : _GEN_264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_266 = 9'h10a == _GEN_9121 ? phv_data_266 : _GEN_265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_267 = 9'h10b == _GEN_9121 ? phv_data_267 : _GEN_266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_268 = 9'h10c == _GEN_9121 ? phv_data_268 : _GEN_267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_269 = 9'h10d == _GEN_9121 ? phv_data_269 : _GEN_268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_270 = 9'h10e == _GEN_9121 ? phv_data_270 : _GEN_269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_271 = 9'h10f == _GEN_9121 ? phv_data_271 : _GEN_270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_272 = 9'h110 == _GEN_9121 ? phv_data_272 : _GEN_271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_273 = 9'h111 == _GEN_9121 ? phv_data_273 : _GEN_272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_274 = 9'h112 == _GEN_9121 ? phv_data_274 : _GEN_273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_275 = 9'h113 == _GEN_9121 ? phv_data_275 : _GEN_274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_276 = 9'h114 == _GEN_9121 ? phv_data_276 : _GEN_275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_277 = 9'h115 == _GEN_9121 ? phv_data_277 : _GEN_276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_278 = 9'h116 == _GEN_9121 ? phv_data_278 : _GEN_277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_279 = 9'h117 == _GEN_9121 ? phv_data_279 : _GEN_278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_280 = 9'h118 == _GEN_9121 ? phv_data_280 : _GEN_279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_281 = 9'h119 == _GEN_9121 ? phv_data_281 : _GEN_280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_282 = 9'h11a == _GEN_9121 ? phv_data_282 : _GEN_281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_283 = 9'h11b == _GEN_9121 ? phv_data_283 : _GEN_282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_284 = 9'h11c == _GEN_9121 ? phv_data_284 : _GEN_283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_285 = 9'h11d == _GEN_9121 ? phv_data_285 : _GEN_284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_286 = 9'h11e == _GEN_9121 ? phv_data_286 : _GEN_285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_287 = 9'h11f == _GEN_9121 ? phv_data_287 : _GEN_286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_288 = 9'h120 == _GEN_9121 ? phv_data_288 : _GEN_287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_289 = 9'h121 == _GEN_9121 ? phv_data_289 : _GEN_288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_290 = 9'h122 == _GEN_9121 ? phv_data_290 : _GEN_289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_291 = 9'h123 == _GEN_9121 ? phv_data_291 : _GEN_290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_292 = 9'h124 == _GEN_9121 ? phv_data_292 : _GEN_291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_293 = 9'h125 == _GEN_9121 ? phv_data_293 : _GEN_292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_294 = 9'h126 == _GEN_9121 ? phv_data_294 : _GEN_293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_295 = 9'h127 == _GEN_9121 ? phv_data_295 : _GEN_294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_296 = 9'h128 == _GEN_9121 ? phv_data_296 : _GEN_295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_297 = 9'h129 == _GEN_9121 ? phv_data_297 : _GEN_296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_298 = 9'h12a == _GEN_9121 ? phv_data_298 : _GEN_297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_299 = 9'h12b == _GEN_9121 ? phv_data_299 : _GEN_298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_300 = 9'h12c == _GEN_9121 ? phv_data_300 : _GEN_299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_301 = 9'h12d == _GEN_9121 ? phv_data_301 : _GEN_300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_302 = 9'h12e == _GEN_9121 ? phv_data_302 : _GEN_301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_303 = 9'h12f == _GEN_9121 ? phv_data_303 : _GEN_302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_304 = 9'h130 == _GEN_9121 ? phv_data_304 : _GEN_303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_305 = 9'h131 == _GEN_9121 ? phv_data_305 : _GEN_304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_306 = 9'h132 == _GEN_9121 ? phv_data_306 : _GEN_305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_307 = 9'h133 == _GEN_9121 ? phv_data_307 : _GEN_306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_308 = 9'h134 == _GEN_9121 ? phv_data_308 : _GEN_307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_309 = 9'h135 == _GEN_9121 ? phv_data_309 : _GEN_308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_310 = 9'h136 == _GEN_9121 ? phv_data_310 : _GEN_309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_311 = 9'h137 == _GEN_9121 ? phv_data_311 : _GEN_310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_312 = 9'h138 == _GEN_9121 ? phv_data_312 : _GEN_311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_313 = 9'h139 == _GEN_9121 ? phv_data_313 : _GEN_312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_314 = 9'h13a == _GEN_9121 ? phv_data_314 : _GEN_313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_315 = 9'h13b == _GEN_9121 ? phv_data_315 : _GEN_314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_316 = 9'h13c == _GEN_9121 ? phv_data_316 : _GEN_315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_317 = 9'h13d == _GEN_9121 ? phv_data_317 : _GEN_316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_318 = 9'h13e == _GEN_9121 ? phv_data_318 : _GEN_317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_319 = 9'h13f == _GEN_9121 ? phv_data_319 : _GEN_318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_320 = 9'h140 == _GEN_9121 ? phv_data_320 : _GEN_319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_321 = 9'h141 == _GEN_9121 ? phv_data_321 : _GEN_320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_322 = 9'h142 == _GEN_9121 ? phv_data_322 : _GEN_321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_323 = 9'h143 == _GEN_9121 ? phv_data_323 : _GEN_322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_324 = 9'h144 == _GEN_9121 ? phv_data_324 : _GEN_323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_325 = 9'h145 == _GEN_9121 ? phv_data_325 : _GEN_324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_326 = 9'h146 == _GEN_9121 ? phv_data_326 : _GEN_325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_327 = 9'h147 == _GEN_9121 ? phv_data_327 : _GEN_326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_328 = 9'h148 == _GEN_9121 ? phv_data_328 : _GEN_327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_329 = 9'h149 == _GEN_9121 ? phv_data_329 : _GEN_328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_330 = 9'h14a == _GEN_9121 ? phv_data_330 : _GEN_329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_331 = 9'h14b == _GEN_9121 ? phv_data_331 : _GEN_330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_332 = 9'h14c == _GEN_9121 ? phv_data_332 : _GEN_331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_333 = 9'h14d == _GEN_9121 ? phv_data_333 : _GEN_332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_334 = 9'h14e == _GEN_9121 ? phv_data_334 : _GEN_333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_335 = 9'h14f == _GEN_9121 ? phv_data_335 : _GEN_334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_336 = 9'h150 == _GEN_9121 ? phv_data_336 : _GEN_335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_337 = 9'h151 == _GEN_9121 ? phv_data_337 : _GEN_336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_338 = 9'h152 == _GEN_9121 ? phv_data_338 : _GEN_337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_339 = 9'h153 == _GEN_9121 ? phv_data_339 : _GEN_338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_340 = 9'h154 == _GEN_9121 ? phv_data_340 : _GEN_339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_341 = 9'h155 == _GEN_9121 ? phv_data_341 : _GEN_340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_342 = 9'h156 == _GEN_9121 ? phv_data_342 : _GEN_341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_343 = 9'h157 == _GEN_9121 ? phv_data_343 : _GEN_342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_344 = 9'h158 == _GEN_9121 ? phv_data_344 : _GEN_343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_345 = 9'h159 == _GEN_9121 ? phv_data_345 : _GEN_344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_346 = 9'h15a == _GEN_9121 ? phv_data_346 : _GEN_345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_347 = 9'h15b == _GEN_9121 ? phv_data_347 : _GEN_346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_348 = 9'h15c == _GEN_9121 ? phv_data_348 : _GEN_347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_349 = 9'h15d == _GEN_9121 ? phv_data_349 : _GEN_348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_350 = 9'h15e == _GEN_9121 ? phv_data_350 : _GEN_349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_351 = 9'h15f == _GEN_9121 ? phv_data_351 : _GEN_350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_352 = 9'h160 == _GEN_9121 ? phv_data_352 : _GEN_351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_353 = 9'h161 == _GEN_9121 ? phv_data_353 : _GEN_352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_354 = 9'h162 == _GEN_9121 ? phv_data_354 : _GEN_353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_355 = 9'h163 == _GEN_9121 ? phv_data_355 : _GEN_354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_356 = 9'h164 == _GEN_9121 ? phv_data_356 : _GEN_355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_357 = 9'h165 == _GEN_9121 ? phv_data_357 : _GEN_356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_358 = 9'h166 == _GEN_9121 ? phv_data_358 : _GEN_357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_359 = 9'h167 == _GEN_9121 ? phv_data_359 : _GEN_358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_360 = 9'h168 == _GEN_9121 ? phv_data_360 : _GEN_359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_361 = 9'h169 == _GEN_9121 ? phv_data_361 : _GEN_360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_362 = 9'h16a == _GEN_9121 ? phv_data_362 : _GEN_361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_363 = 9'h16b == _GEN_9121 ? phv_data_363 : _GEN_362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_364 = 9'h16c == _GEN_9121 ? phv_data_364 : _GEN_363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_365 = 9'h16d == _GEN_9121 ? phv_data_365 : _GEN_364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_366 = 9'h16e == _GEN_9121 ? phv_data_366 : _GEN_365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_367 = 9'h16f == _GEN_9121 ? phv_data_367 : _GEN_366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_368 = 9'h170 == _GEN_9121 ? phv_data_368 : _GEN_367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_369 = 9'h171 == _GEN_9121 ? phv_data_369 : _GEN_368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_370 = 9'h172 == _GEN_9121 ? phv_data_370 : _GEN_369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_371 = 9'h173 == _GEN_9121 ? phv_data_371 : _GEN_370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_372 = 9'h174 == _GEN_9121 ? phv_data_372 : _GEN_371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_373 = 9'h175 == _GEN_9121 ? phv_data_373 : _GEN_372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_374 = 9'h176 == _GEN_9121 ? phv_data_374 : _GEN_373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_375 = 9'h177 == _GEN_9121 ? phv_data_375 : _GEN_374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_376 = 9'h178 == _GEN_9121 ? phv_data_376 : _GEN_375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_377 = 9'h179 == _GEN_9121 ? phv_data_377 : _GEN_376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_378 = 9'h17a == _GEN_9121 ? phv_data_378 : _GEN_377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_379 = 9'h17b == _GEN_9121 ? phv_data_379 : _GEN_378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_380 = 9'h17c == _GEN_9121 ? phv_data_380 : _GEN_379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_381 = 9'h17d == _GEN_9121 ? phv_data_381 : _GEN_380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_382 = 9'h17e == _GEN_9121 ? phv_data_382 : _GEN_381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_383 = 9'h17f == _GEN_9121 ? phv_data_383 : _GEN_382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_384 = 9'h180 == _GEN_9121 ? phv_data_384 : _GEN_383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_385 = 9'h181 == _GEN_9121 ? phv_data_385 : _GEN_384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_386 = 9'h182 == _GEN_9121 ? phv_data_386 : _GEN_385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_387 = 9'h183 == _GEN_9121 ? phv_data_387 : _GEN_386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_388 = 9'h184 == _GEN_9121 ? phv_data_388 : _GEN_387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_389 = 9'h185 == _GEN_9121 ? phv_data_389 : _GEN_388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_390 = 9'h186 == _GEN_9121 ? phv_data_390 : _GEN_389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_391 = 9'h187 == _GEN_9121 ? phv_data_391 : _GEN_390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_392 = 9'h188 == _GEN_9121 ? phv_data_392 : _GEN_391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_393 = 9'h189 == _GEN_9121 ? phv_data_393 : _GEN_392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_394 = 9'h18a == _GEN_9121 ? phv_data_394 : _GEN_393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_395 = 9'h18b == _GEN_9121 ? phv_data_395 : _GEN_394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_396 = 9'h18c == _GEN_9121 ? phv_data_396 : _GEN_395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_397 = 9'h18d == _GEN_9121 ? phv_data_397 : _GEN_396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_398 = 9'h18e == _GEN_9121 ? phv_data_398 : _GEN_397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_399 = 9'h18f == _GEN_9121 ? phv_data_399 : _GEN_398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_400 = 9'h190 == _GEN_9121 ? phv_data_400 : _GEN_399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_401 = 9'h191 == _GEN_9121 ? phv_data_401 : _GEN_400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_402 = 9'h192 == _GEN_9121 ? phv_data_402 : _GEN_401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_403 = 9'h193 == _GEN_9121 ? phv_data_403 : _GEN_402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_404 = 9'h194 == _GEN_9121 ? phv_data_404 : _GEN_403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_405 = 9'h195 == _GEN_9121 ? phv_data_405 : _GEN_404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_406 = 9'h196 == _GEN_9121 ? phv_data_406 : _GEN_405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_407 = 9'h197 == _GEN_9121 ? phv_data_407 : _GEN_406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_408 = 9'h198 == _GEN_9121 ? phv_data_408 : _GEN_407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_409 = 9'h199 == _GEN_9121 ? phv_data_409 : _GEN_408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_410 = 9'h19a == _GEN_9121 ? phv_data_410 : _GEN_409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_411 = 9'h19b == _GEN_9121 ? phv_data_411 : _GEN_410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_412 = 9'h19c == _GEN_9121 ? phv_data_412 : _GEN_411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_413 = 9'h19d == _GEN_9121 ? phv_data_413 : _GEN_412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_414 = 9'h19e == _GEN_9121 ? phv_data_414 : _GEN_413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_415 = 9'h19f == _GEN_9121 ? phv_data_415 : _GEN_414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_416 = 9'h1a0 == _GEN_9121 ? phv_data_416 : _GEN_415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_417 = 9'h1a1 == _GEN_9121 ? phv_data_417 : _GEN_416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_418 = 9'h1a2 == _GEN_9121 ? phv_data_418 : _GEN_417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_419 = 9'h1a3 == _GEN_9121 ? phv_data_419 : _GEN_418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_420 = 9'h1a4 == _GEN_9121 ? phv_data_420 : _GEN_419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_421 = 9'h1a5 == _GEN_9121 ? phv_data_421 : _GEN_420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_422 = 9'h1a6 == _GEN_9121 ? phv_data_422 : _GEN_421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_423 = 9'h1a7 == _GEN_9121 ? phv_data_423 : _GEN_422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_424 = 9'h1a8 == _GEN_9121 ? phv_data_424 : _GEN_423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_425 = 9'h1a9 == _GEN_9121 ? phv_data_425 : _GEN_424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_426 = 9'h1aa == _GEN_9121 ? phv_data_426 : _GEN_425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_427 = 9'h1ab == _GEN_9121 ? phv_data_427 : _GEN_426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_428 = 9'h1ac == _GEN_9121 ? phv_data_428 : _GEN_427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_429 = 9'h1ad == _GEN_9121 ? phv_data_429 : _GEN_428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_430 = 9'h1ae == _GEN_9121 ? phv_data_430 : _GEN_429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_431 = 9'h1af == _GEN_9121 ? phv_data_431 : _GEN_430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_432 = 9'h1b0 == _GEN_9121 ? phv_data_432 : _GEN_431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_433 = 9'h1b1 == _GEN_9121 ? phv_data_433 : _GEN_432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_434 = 9'h1b2 == _GEN_9121 ? phv_data_434 : _GEN_433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_435 = 9'h1b3 == _GEN_9121 ? phv_data_435 : _GEN_434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_436 = 9'h1b4 == _GEN_9121 ? phv_data_436 : _GEN_435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_437 = 9'h1b5 == _GEN_9121 ? phv_data_437 : _GEN_436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_438 = 9'h1b6 == _GEN_9121 ? phv_data_438 : _GEN_437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_439 = 9'h1b7 == _GEN_9121 ? phv_data_439 : _GEN_438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_440 = 9'h1b8 == _GEN_9121 ? phv_data_440 : _GEN_439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_441 = 9'h1b9 == _GEN_9121 ? phv_data_441 : _GEN_440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_442 = 9'h1ba == _GEN_9121 ? phv_data_442 : _GEN_441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_443 = 9'h1bb == _GEN_9121 ? phv_data_443 : _GEN_442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_444 = 9'h1bc == _GEN_9121 ? phv_data_444 : _GEN_443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_445 = 9'h1bd == _GEN_9121 ? phv_data_445 : _GEN_444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_446 = 9'h1be == _GEN_9121 ? phv_data_446 : _GEN_445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_447 = 9'h1bf == _GEN_9121 ? phv_data_447 : _GEN_446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_448 = 9'h1c0 == _GEN_9121 ? phv_data_448 : _GEN_447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_449 = 9'h1c1 == _GEN_9121 ? phv_data_449 : _GEN_448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_450 = 9'h1c2 == _GEN_9121 ? phv_data_450 : _GEN_449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_451 = 9'h1c3 == _GEN_9121 ? phv_data_451 : _GEN_450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_452 = 9'h1c4 == _GEN_9121 ? phv_data_452 : _GEN_451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_453 = 9'h1c5 == _GEN_9121 ? phv_data_453 : _GEN_452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_454 = 9'h1c6 == _GEN_9121 ? phv_data_454 : _GEN_453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_455 = 9'h1c7 == _GEN_9121 ? phv_data_455 : _GEN_454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_456 = 9'h1c8 == _GEN_9121 ? phv_data_456 : _GEN_455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_457 = 9'h1c9 == _GEN_9121 ? phv_data_457 : _GEN_456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_458 = 9'h1ca == _GEN_9121 ? phv_data_458 : _GEN_457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_459 = 9'h1cb == _GEN_9121 ? phv_data_459 : _GEN_458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_460 = 9'h1cc == _GEN_9121 ? phv_data_460 : _GEN_459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_461 = 9'h1cd == _GEN_9121 ? phv_data_461 : _GEN_460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_462 = 9'h1ce == _GEN_9121 ? phv_data_462 : _GEN_461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_463 = 9'h1cf == _GEN_9121 ? phv_data_463 : _GEN_462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_464 = 9'h1d0 == _GEN_9121 ? phv_data_464 : _GEN_463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_465 = 9'h1d1 == _GEN_9121 ? phv_data_465 : _GEN_464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_466 = 9'h1d2 == _GEN_9121 ? phv_data_466 : _GEN_465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_467 = 9'h1d3 == _GEN_9121 ? phv_data_467 : _GEN_466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_468 = 9'h1d4 == _GEN_9121 ? phv_data_468 : _GEN_467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_469 = 9'h1d5 == _GEN_9121 ? phv_data_469 : _GEN_468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_470 = 9'h1d6 == _GEN_9121 ? phv_data_470 : _GEN_469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_471 = 9'h1d7 == _GEN_9121 ? phv_data_471 : _GEN_470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_472 = 9'h1d8 == _GEN_9121 ? phv_data_472 : _GEN_471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_473 = 9'h1d9 == _GEN_9121 ? phv_data_473 : _GEN_472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_474 = 9'h1da == _GEN_9121 ? phv_data_474 : _GEN_473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_475 = 9'h1db == _GEN_9121 ? phv_data_475 : _GEN_474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_476 = 9'h1dc == _GEN_9121 ? phv_data_476 : _GEN_475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_477 = 9'h1dd == _GEN_9121 ? phv_data_477 : _GEN_476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_478 = 9'h1de == _GEN_9121 ? phv_data_478 : _GEN_477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_479 = 9'h1df == _GEN_9121 ? phv_data_479 : _GEN_478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_480 = 9'h1e0 == _GEN_9121 ? phv_data_480 : _GEN_479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_481 = 9'h1e1 == _GEN_9121 ? phv_data_481 : _GEN_480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_482 = 9'h1e2 == _GEN_9121 ? phv_data_482 : _GEN_481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_483 = 9'h1e3 == _GEN_9121 ? phv_data_483 : _GEN_482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_484 = 9'h1e4 == _GEN_9121 ? phv_data_484 : _GEN_483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_485 = 9'h1e5 == _GEN_9121 ? phv_data_485 : _GEN_484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_486 = 9'h1e6 == _GEN_9121 ? phv_data_486 : _GEN_485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_487 = 9'h1e7 == _GEN_9121 ? phv_data_487 : _GEN_486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_488 = 9'h1e8 == _GEN_9121 ? phv_data_488 : _GEN_487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_489 = 9'h1e9 == _GEN_9121 ? phv_data_489 : _GEN_488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_490 = 9'h1ea == _GEN_9121 ? phv_data_490 : _GEN_489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_491 = 9'h1eb == _GEN_9121 ? phv_data_491 : _GEN_490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_492 = 9'h1ec == _GEN_9121 ? phv_data_492 : _GEN_491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_493 = 9'h1ed == _GEN_9121 ? phv_data_493 : _GEN_492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_494 = 9'h1ee == _GEN_9121 ? phv_data_494 : _GEN_493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_495 = 9'h1ef == _GEN_9121 ? phv_data_495 : _GEN_494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_496 = 9'h1f0 == _GEN_9121 ? phv_data_496 : _GEN_495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_497 = 9'h1f1 == _GEN_9121 ? phv_data_497 : _GEN_496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_498 = 9'h1f2 == _GEN_9121 ? phv_data_498 : _GEN_497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_499 = 9'h1f3 == _GEN_9121 ? phv_data_499 : _GEN_498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_500 = 9'h1f4 == _GEN_9121 ? phv_data_500 : _GEN_499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_501 = 9'h1f5 == _GEN_9121 ? phv_data_501 : _GEN_500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_502 = 9'h1f6 == _GEN_9121 ? phv_data_502 : _GEN_501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_503 = 9'h1f7 == _GEN_9121 ? phv_data_503 : _GEN_502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_504 = 9'h1f8 == _GEN_9121 ? phv_data_504 : _GEN_503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_505 = 9'h1f9 == _GEN_9121 ? phv_data_505 : _GEN_504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_506 = 9'h1fa == _GEN_9121 ? phv_data_506 : _GEN_505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_507 = 9'h1fb == _GEN_9121 ? phv_data_507 : _GEN_506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_508 = 9'h1fc == _GEN_9121 ? phv_data_508 : _GEN_507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_509 = 9'h1fd == _GEN_9121 ? phv_data_509 : _GEN_508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_510 = 9'h1fe == _GEN_9121 ? phv_data_510 : _GEN_509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__3 = 9'h1ff == _GEN_9121 ? phv_data_511 : _GEN_510; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_3 = ending == 2'h0; // @[executor.scala 199:88]
  wire  mask__3 = 2'h0 >= offset_0[1:0] & (2'h0 < ending | ending == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_1 = {total_offset_hi,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_513 = 8'h1 == total_offset_1 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_514 = 8'h2 == total_offset_1 ? phv_data_2 : _GEN_513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_515 = 8'h3 == total_offset_1 ? phv_data_3 : _GEN_514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_516 = 8'h4 == total_offset_1 ? phv_data_4 : _GEN_515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_517 = 8'h5 == total_offset_1 ? phv_data_5 : _GEN_516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_518 = 8'h6 == total_offset_1 ? phv_data_6 : _GEN_517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_519 = 8'h7 == total_offset_1 ? phv_data_7 : _GEN_518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_520 = 8'h8 == total_offset_1 ? phv_data_8 : _GEN_519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_521 = 8'h9 == total_offset_1 ? phv_data_9 : _GEN_520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_522 = 8'ha == total_offset_1 ? phv_data_10 : _GEN_521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_523 = 8'hb == total_offset_1 ? phv_data_11 : _GEN_522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_524 = 8'hc == total_offset_1 ? phv_data_12 : _GEN_523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_525 = 8'hd == total_offset_1 ? phv_data_13 : _GEN_524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_526 = 8'he == total_offset_1 ? phv_data_14 : _GEN_525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_527 = 8'hf == total_offset_1 ? phv_data_15 : _GEN_526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_528 = 8'h10 == total_offset_1 ? phv_data_16 : _GEN_527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_529 = 8'h11 == total_offset_1 ? phv_data_17 : _GEN_528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_530 = 8'h12 == total_offset_1 ? phv_data_18 : _GEN_529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_531 = 8'h13 == total_offset_1 ? phv_data_19 : _GEN_530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_532 = 8'h14 == total_offset_1 ? phv_data_20 : _GEN_531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_533 = 8'h15 == total_offset_1 ? phv_data_21 : _GEN_532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_534 = 8'h16 == total_offset_1 ? phv_data_22 : _GEN_533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_535 = 8'h17 == total_offset_1 ? phv_data_23 : _GEN_534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_536 = 8'h18 == total_offset_1 ? phv_data_24 : _GEN_535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_537 = 8'h19 == total_offset_1 ? phv_data_25 : _GEN_536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_538 = 8'h1a == total_offset_1 ? phv_data_26 : _GEN_537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_539 = 8'h1b == total_offset_1 ? phv_data_27 : _GEN_538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_540 = 8'h1c == total_offset_1 ? phv_data_28 : _GEN_539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_541 = 8'h1d == total_offset_1 ? phv_data_29 : _GEN_540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_542 = 8'h1e == total_offset_1 ? phv_data_30 : _GEN_541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_543 = 8'h1f == total_offset_1 ? phv_data_31 : _GEN_542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_544 = 8'h20 == total_offset_1 ? phv_data_32 : _GEN_543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_545 = 8'h21 == total_offset_1 ? phv_data_33 : _GEN_544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_546 = 8'h22 == total_offset_1 ? phv_data_34 : _GEN_545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_547 = 8'h23 == total_offset_1 ? phv_data_35 : _GEN_546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_548 = 8'h24 == total_offset_1 ? phv_data_36 : _GEN_547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_549 = 8'h25 == total_offset_1 ? phv_data_37 : _GEN_548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_550 = 8'h26 == total_offset_1 ? phv_data_38 : _GEN_549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_551 = 8'h27 == total_offset_1 ? phv_data_39 : _GEN_550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_552 = 8'h28 == total_offset_1 ? phv_data_40 : _GEN_551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_553 = 8'h29 == total_offset_1 ? phv_data_41 : _GEN_552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_554 = 8'h2a == total_offset_1 ? phv_data_42 : _GEN_553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_555 = 8'h2b == total_offset_1 ? phv_data_43 : _GEN_554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_556 = 8'h2c == total_offset_1 ? phv_data_44 : _GEN_555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_557 = 8'h2d == total_offset_1 ? phv_data_45 : _GEN_556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_558 = 8'h2e == total_offset_1 ? phv_data_46 : _GEN_557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_559 = 8'h2f == total_offset_1 ? phv_data_47 : _GEN_558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_560 = 8'h30 == total_offset_1 ? phv_data_48 : _GEN_559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_561 = 8'h31 == total_offset_1 ? phv_data_49 : _GEN_560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_562 = 8'h32 == total_offset_1 ? phv_data_50 : _GEN_561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_563 = 8'h33 == total_offset_1 ? phv_data_51 : _GEN_562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_564 = 8'h34 == total_offset_1 ? phv_data_52 : _GEN_563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_565 = 8'h35 == total_offset_1 ? phv_data_53 : _GEN_564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_566 = 8'h36 == total_offset_1 ? phv_data_54 : _GEN_565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_567 = 8'h37 == total_offset_1 ? phv_data_55 : _GEN_566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_568 = 8'h38 == total_offset_1 ? phv_data_56 : _GEN_567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_569 = 8'h39 == total_offset_1 ? phv_data_57 : _GEN_568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_570 = 8'h3a == total_offset_1 ? phv_data_58 : _GEN_569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_571 = 8'h3b == total_offset_1 ? phv_data_59 : _GEN_570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_572 = 8'h3c == total_offset_1 ? phv_data_60 : _GEN_571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_573 = 8'h3d == total_offset_1 ? phv_data_61 : _GEN_572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_574 = 8'h3e == total_offset_1 ? phv_data_62 : _GEN_573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_575 = 8'h3f == total_offset_1 ? phv_data_63 : _GEN_574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_576 = 8'h40 == total_offset_1 ? phv_data_64 : _GEN_575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_577 = 8'h41 == total_offset_1 ? phv_data_65 : _GEN_576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_578 = 8'h42 == total_offset_1 ? phv_data_66 : _GEN_577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_579 = 8'h43 == total_offset_1 ? phv_data_67 : _GEN_578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_580 = 8'h44 == total_offset_1 ? phv_data_68 : _GEN_579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_581 = 8'h45 == total_offset_1 ? phv_data_69 : _GEN_580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_582 = 8'h46 == total_offset_1 ? phv_data_70 : _GEN_581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_583 = 8'h47 == total_offset_1 ? phv_data_71 : _GEN_582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_584 = 8'h48 == total_offset_1 ? phv_data_72 : _GEN_583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_585 = 8'h49 == total_offset_1 ? phv_data_73 : _GEN_584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_586 = 8'h4a == total_offset_1 ? phv_data_74 : _GEN_585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_587 = 8'h4b == total_offset_1 ? phv_data_75 : _GEN_586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_588 = 8'h4c == total_offset_1 ? phv_data_76 : _GEN_587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_589 = 8'h4d == total_offset_1 ? phv_data_77 : _GEN_588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_590 = 8'h4e == total_offset_1 ? phv_data_78 : _GEN_589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_591 = 8'h4f == total_offset_1 ? phv_data_79 : _GEN_590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_592 = 8'h50 == total_offset_1 ? phv_data_80 : _GEN_591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_593 = 8'h51 == total_offset_1 ? phv_data_81 : _GEN_592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_594 = 8'h52 == total_offset_1 ? phv_data_82 : _GEN_593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_595 = 8'h53 == total_offset_1 ? phv_data_83 : _GEN_594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_596 = 8'h54 == total_offset_1 ? phv_data_84 : _GEN_595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_597 = 8'h55 == total_offset_1 ? phv_data_85 : _GEN_596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_598 = 8'h56 == total_offset_1 ? phv_data_86 : _GEN_597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_599 = 8'h57 == total_offset_1 ? phv_data_87 : _GEN_598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_600 = 8'h58 == total_offset_1 ? phv_data_88 : _GEN_599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_601 = 8'h59 == total_offset_1 ? phv_data_89 : _GEN_600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_602 = 8'h5a == total_offset_1 ? phv_data_90 : _GEN_601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_603 = 8'h5b == total_offset_1 ? phv_data_91 : _GEN_602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_604 = 8'h5c == total_offset_1 ? phv_data_92 : _GEN_603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_605 = 8'h5d == total_offset_1 ? phv_data_93 : _GEN_604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_606 = 8'h5e == total_offset_1 ? phv_data_94 : _GEN_605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_607 = 8'h5f == total_offset_1 ? phv_data_95 : _GEN_606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_608 = 8'h60 == total_offset_1 ? phv_data_96 : _GEN_607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_609 = 8'h61 == total_offset_1 ? phv_data_97 : _GEN_608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_610 = 8'h62 == total_offset_1 ? phv_data_98 : _GEN_609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_611 = 8'h63 == total_offset_1 ? phv_data_99 : _GEN_610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_612 = 8'h64 == total_offset_1 ? phv_data_100 : _GEN_611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_613 = 8'h65 == total_offset_1 ? phv_data_101 : _GEN_612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_614 = 8'h66 == total_offset_1 ? phv_data_102 : _GEN_613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_615 = 8'h67 == total_offset_1 ? phv_data_103 : _GEN_614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_616 = 8'h68 == total_offset_1 ? phv_data_104 : _GEN_615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_617 = 8'h69 == total_offset_1 ? phv_data_105 : _GEN_616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_618 = 8'h6a == total_offset_1 ? phv_data_106 : _GEN_617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_619 = 8'h6b == total_offset_1 ? phv_data_107 : _GEN_618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_620 = 8'h6c == total_offset_1 ? phv_data_108 : _GEN_619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_621 = 8'h6d == total_offset_1 ? phv_data_109 : _GEN_620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_622 = 8'h6e == total_offset_1 ? phv_data_110 : _GEN_621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_623 = 8'h6f == total_offset_1 ? phv_data_111 : _GEN_622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_624 = 8'h70 == total_offset_1 ? phv_data_112 : _GEN_623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_625 = 8'h71 == total_offset_1 ? phv_data_113 : _GEN_624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_626 = 8'h72 == total_offset_1 ? phv_data_114 : _GEN_625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_627 = 8'h73 == total_offset_1 ? phv_data_115 : _GEN_626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_628 = 8'h74 == total_offset_1 ? phv_data_116 : _GEN_627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_629 = 8'h75 == total_offset_1 ? phv_data_117 : _GEN_628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_630 = 8'h76 == total_offset_1 ? phv_data_118 : _GEN_629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_631 = 8'h77 == total_offset_1 ? phv_data_119 : _GEN_630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_632 = 8'h78 == total_offset_1 ? phv_data_120 : _GEN_631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_633 = 8'h79 == total_offset_1 ? phv_data_121 : _GEN_632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_634 = 8'h7a == total_offset_1 ? phv_data_122 : _GEN_633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_635 = 8'h7b == total_offset_1 ? phv_data_123 : _GEN_634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_636 = 8'h7c == total_offset_1 ? phv_data_124 : _GEN_635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_637 = 8'h7d == total_offset_1 ? phv_data_125 : _GEN_636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_638 = 8'h7e == total_offset_1 ? phv_data_126 : _GEN_637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_639 = 8'h7f == total_offset_1 ? phv_data_127 : _GEN_638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_640 = 8'h80 == total_offset_1 ? phv_data_128 : _GEN_639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_641 = 8'h81 == total_offset_1 ? phv_data_129 : _GEN_640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_642 = 8'h82 == total_offset_1 ? phv_data_130 : _GEN_641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_643 = 8'h83 == total_offset_1 ? phv_data_131 : _GEN_642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_644 = 8'h84 == total_offset_1 ? phv_data_132 : _GEN_643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_645 = 8'h85 == total_offset_1 ? phv_data_133 : _GEN_644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_646 = 8'h86 == total_offset_1 ? phv_data_134 : _GEN_645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_647 = 8'h87 == total_offset_1 ? phv_data_135 : _GEN_646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_648 = 8'h88 == total_offset_1 ? phv_data_136 : _GEN_647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_649 = 8'h89 == total_offset_1 ? phv_data_137 : _GEN_648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_650 = 8'h8a == total_offset_1 ? phv_data_138 : _GEN_649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_651 = 8'h8b == total_offset_1 ? phv_data_139 : _GEN_650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_652 = 8'h8c == total_offset_1 ? phv_data_140 : _GEN_651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_653 = 8'h8d == total_offset_1 ? phv_data_141 : _GEN_652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_654 = 8'h8e == total_offset_1 ? phv_data_142 : _GEN_653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_655 = 8'h8f == total_offset_1 ? phv_data_143 : _GEN_654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_656 = 8'h90 == total_offset_1 ? phv_data_144 : _GEN_655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_657 = 8'h91 == total_offset_1 ? phv_data_145 : _GEN_656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_658 = 8'h92 == total_offset_1 ? phv_data_146 : _GEN_657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_659 = 8'h93 == total_offset_1 ? phv_data_147 : _GEN_658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_660 = 8'h94 == total_offset_1 ? phv_data_148 : _GEN_659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_661 = 8'h95 == total_offset_1 ? phv_data_149 : _GEN_660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_662 = 8'h96 == total_offset_1 ? phv_data_150 : _GEN_661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_663 = 8'h97 == total_offset_1 ? phv_data_151 : _GEN_662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_664 = 8'h98 == total_offset_1 ? phv_data_152 : _GEN_663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_665 = 8'h99 == total_offset_1 ? phv_data_153 : _GEN_664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_666 = 8'h9a == total_offset_1 ? phv_data_154 : _GEN_665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_667 = 8'h9b == total_offset_1 ? phv_data_155 : _GEN_666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_668 = 8'h9c == total_offset_1 ? phv_data_156 : _GEN_667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_669 = 8'h9d == total_offset_1 ? phv_data_157 : _GEN_668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_670 = 8'h9e == total_offset_1 ? phv_data_158 : _GEN_669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_671 = 8'h9f == total_offset_1 ? phv_data_159 : _GEN_670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_672 = 8'ha0 == total_offset_1 ? phv_data_160 : _GEN_671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_673 = 8'ha1 == total_offset_1 ? phv_data_161 : _GEN_672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_674 = 8'ha2 == total_offset_1 ? phv_data_162 : _GEN_673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_675 = 8'ha3 == total_offset_1 ? phv_data_163 : _GEN_674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_676 = 8'ha4 == total_offset_1 ? phv_data_164 : _GEN_675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_677 = 8'ha5 == total_offset_1 ? phv_data_165 : _GEN_676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_678 = 8'ha6 == total_offset_1 ? phv_data_166 : _GEN_677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_679 = 8'ha7 == total_offset_1 ? phv_data_167 : _GEN_678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_680 = 8'ha8 == total_offset_1 ? phv_data_168 : _GEN_679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_681 = 8'ha9 == total_offset_1 ? phv_data_169 : _GEN_680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_682 = 8'haa == total_offset_1 ? phv_data_170 : _GEN_681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_683 = 8'hab == total_offset_1 ? phv_data_171 : _GEN_682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_684 = 8'hac == total_offset_1 ? phv_data_172 : _GEN_683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_685 = 8'had == total_offset_1 ? phv_data_173 : _GEN_684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_686 = 8'hae == total_offset_1 ? phv_data_174 : _GEN_685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_687 = 8'haf == total_offset_1 ? phv_data_175 : _GEN_686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_688 = 8'hb0 == total_offset_1 ? phv_data_176 : _GEN_687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_689 = 8'hb1 == total_offset_1 ? phv_data_177 : _GEN_688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_690 = 8'hb2 == total_offset_1 ? phv_data_178 : _GEN_689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_691 = 8'hb3 == total_offset_1 ? phv_data_179 : _GEN_690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_692 = 8'hb4 == total_offset_1 ? phv_data_180 : _GEN_691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_693 = 8'hb5 == total_offset_1 ? phv_data_181 : _GEN_692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_694 = 8'hb6 == total_offset_1 ? phv_data_182 : _GEN_693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_695 = 8'hb7 == total_offset_1 ? phv_data_183 : _GEN_694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_696 = 8'hb8 == total_offset_1 ? phv_data_184 : _GEN_695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_697 = 8'hb9 == total_offset_1 ? phv_data_185 : _GEN_696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_698 = 8'hba == total_offset_1 ? phv_data_186 : _GEN_697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_699 = 8'hbb == total_offset_1 ? phv_data_187 : _GEN_698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_700 = 8'hbc == total_offset_1 ? phv_data_188 : _GEN_699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_701 = 8'hbd == total_offset_1 ? phv_data_189 : _GEN_700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_702 = 8'hbe == total_offset_1 ? phv_data_190 : _GEN_701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_703 = 8'hbf == total_offset_1 ? phv_data_191 : _GEN_702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_704 = 8'hc0 == total_offset_1 ? phv_data_192 : _GEN_703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_705 = 8'hc1 == total_offset_1 ? phv_data_193 : _GEN_704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_706 = 8'hc2 == total_offset_1 ? phv_data_194 : _GEN_705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_707 = 8'hc3 == total_offset_1 ? phv_data_195 : _GEN_706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_708 = 8'hc4 == total_offset_1 ? phv_data_196 : _GEN_707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_709 = 8'hc5 == total_offset_1 ? phv_data_197 : _GEN_708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_710 = 8'hc6 == total_offset_1 ? phv_data_198 : _GEN_709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_711 = 8'hc7 == total_offset_1 ? phv_data_199 : _GEN_710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_712 = 8'hc8 == total_offset_1 ? phv_data_200 : _GEN_711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_713 = 8'hc9 == total_offset_1 ? phv_data_201 : _GEN_712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_714 = 8'hca == total_offset_1 ? phv_data_202 : _GEN_713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_715 = 8'hcb == total_offset_1 ? phv_data_203 : _GEN_714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_716 = 8'hcc == total_offset_1 ? phv_data_204 : _GEN_715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_717 = 8'hcd == total_offset_1 ? phv_data_205 : _GEN_716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_718 = 8'hce == total_offset_1 ? phv_data_206 : _GEN_717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_719 = 8'hcf == total_offset_1 ? phv_data_207 : _GEN_718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_720 = 8'hd0 == total_offset_1 ? phv_data_208 : _GEN_719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_721 = 8'hd1 == total_offset_1 ? phv_data_209 : _GEN_720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_722 = 8'hd2 == total_offset_1 ? phv_data_210 : _GEN_721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_723 = 8'hd3 == total_offset_1 ? phv_data_211 : _GEN_722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_724 = 8'hd4 == total_offset_1 ? phv_data_212 : _GEN_723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_725 = 8'hd5 == total_offset_1 ? phv_data_213 : _GEN_724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_726 = 8'hd6 == total_offset_1 ? phv_data_214 : _GEN_725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_727 = 8'hd7 == total_offset_1 ? phv_data_215 : _GEN_726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_728 = 8'hd8 == total_offset_1 ? phv_data_216 : _GEN_727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_729 = 8'hd9 == total_offset_1 ? phv_data_217 : _GEN_728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_730 = 8'hda == total_offset_1 ? phv_data_218 : _GEN_729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_731 = 8'hdb == total_offset_1 ? phv_data_219 : _GEN_730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_732 = 8'hdc == total_offset_1 ? phv_data_220 : _GEN_731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_733 = 8'hdd == total_offset_1 ? phv_data_221 : _GEN_732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_734 = 8'hde == total_offset_1 ? phv_data_222 : _GEN_733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_735 = 8'hdf == total_offset_1 ? phv_data_223 : _GEN_734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_736 = 8'he0 == total_offset_1 ? phv_data_224 : _GEN_735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_737 = 8'he1 == total_offset_1 ? phv_data_225 : _GEN_736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_738 = 8'he2 == total_offset_1 ? phv_data_226 : _GEN_737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_739 = 8'he3 == total_offset_1 ? phv_data_227 : _GEN_738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_740 = 8'he4 == total_offset_1 ? phv_data_228 : _GEN_739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_741 = 8'he5 == total_offset_1 ? phv_data_229 : _GEN_740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_742 = 8'he6 == total_offset_1 ? phv_data_230 : _GEN_741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_743 = 8'he7 == total_offset_1 ? phv_data_231 : _GEN_742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_744 = 8'he8 == total_offset_1 ? phv_data_232 : _GEN_743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_745 = 8'he9 == total_offset_1 ? phv_data_233 : _GEN_744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_746 = 8'hea == total_offset_1 ? phv_data_234 : _GEN_745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_747 = 8'heb == total_offset_1 ? phv_data_235 : _GEN_746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_748 = 8'hec == total_offset_1 ? phv_data_236 : _GEN_747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_749 = 8'hed == total_offset_1 ? phv_data_237 : _GEN_748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_750 = 8'hee == total_offset_1 ? phv_data_238 : _GEN_749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_751 = 8'hef == total_offset_1 ? phv_data_239 : _GEN_750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_752 = 8'hf0 == total_offset_1 ? phv_data_240 : _GEN_751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_753 = 8'hf1 == total_offset_1 ? phv_data_241 : _GEN_752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_754 = 8'hf2 == total_offset_1 ? phv_data_242 : _GEN_753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_755 = 8'hf3 == total_offset_1 ? phv_data_243 : _GEN_754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_756 = 8'hf4 == total_offset_1 ? phv_data_244 : _GEN_755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_757 = 8'hf5 == total_offset_1 ? phv_data_245 : _GEN_756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_758 = 8'hf6 == total_offset_1 ? phv_data_246 : _GEN_757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_759 = 8'hf7 == total_offset_1 ? phv_data_247 : _GEN_758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_760 = 8'hf8 == total_offset_1 ? phv_data_248 : _GEN_759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_761 = 8'hf9 == total_offset_1 ? phv_data_249 : _GEN_760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_762 = 8'hfa == total_offset_1 ? phv_data_250 : _GEN_761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_763 = 8'hfb == total_offset_1 ? phv_data_251 : _GEN_762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_764 = 8'hfc == total_offset_1 ? phv_data_252 : _GEN_763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_765 = 8'hfd == total_offset_1 ? phv_data_253 : _GEN_764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_766 = 8'hfe == total_offset_1 ? phv_data_254 : _GEN_765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_767 = 8'hff == total_offset_1 ? phv_data_255 : _GEN_766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_9377 = {{1'd0}, total_offset_1}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_768 = 9'h100 == _GEN_9377 ? phv_data_256 : _GEN_767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_769 = 9'h101 == _GEN_9377 ? phv_data_257 : _GEN_768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_770 = 9'h102 == _GEN_9377 ? phv_data_258 : _GEN_769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_771 = 9'h103 == _GEN_9377 ? phv_data_259 : _GEN_770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_772 = 9'h104 == _GEN_9377 ? phv_data_260 : _GEN_771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_773 = 9'h105 == _GEN_9377 ? phv_data_261 : _GEN_772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_774 = 9'h106 == _GEN_9377 ? phv_data_262 : _GEN_773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_775 = 9'h107 == _GEN_9377 ? phv_data_263 : _GEN_774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_776 = 9'h108 == _GEN_9377 ? phv_data_264 : _GEN_775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_777 = 9'h109 == _GEN_9377 ? phv_data_265 : _GEN_776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_778 = 9'h10a == _GEN_9377 ? phv_data_266 : _GEN_777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_779 = 9'h10b == _GEN_9377 ? phv_data_267 : _GEN_778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_780 = 9'h10c == _GEN_9377 ? phv_data_268 : _GEN_779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_781 = 9'h10d == _GEN_9377 ? phv_data_269 : _GEN_780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_782 = 9'h10e == _GEN_9377 ? phv_data_270 : _GEN_781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_783 = 9'h10f == _GEN_9377 ? phv_data_271 : _GEN_782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_784 = 9'h110 == _GEN_9377 ? phv_data_272 : _GEN_783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_785 = 9'h111 == _GEN_9377 ? phv_data_273 : _GEN_784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_786 = 9'h112 == _GEN_9377 ? phv_data_274 : _GEN_785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_787 = 9'h113 == _GEN_9377 ? phv_data_275 : _GEN_786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_788 = 9'h114 == _GEN_9377 ? phv_data_276 : _GEN_787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_789 = 9'h115 == _GEN_9377 ? phv_data_277 : _GEN_788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_790 = 9'h116 == _GEN_9377 ? phv_data_278 : _GEN_789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_791 = 9'h117 == _GEN_9377 ? phv_data_279 : _GEN_790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_792 = 9'h118 == _GEN_9377 ? phv_data_280 : _GEN_791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_793 = 9'h119 == _GEN_9377 ? phv_data_281 : _GEN_792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_794 = 9'h11a == _GEN_9377 ? phv_data_282 : _GEN_793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_795 = 9'h11b == _GEN_9377 ? phv_data_283 : _GEN_794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_796 = 9'h11c == _GEN_9377 ? phv_data_284 : _GEN_795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_797 = 9'h11d == _GEN_9377 ? phv_data_285 : _GEN_796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_798 = 9'h11e == _GEN_9377 ? phv_data_286 : _GEN_797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_799 = 9'h11f == _GEN_9377 ? phv_data_287 : _GEN_798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_800 = 9'h120 == _GEN_9377 ? phv_data_288 : _GEN_799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_801 = 9'h121 == _GEN_9377 ? phv_data_289 : _GEN_800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_802 = 9'h122 == _GEN_9377 ? phv_data_290 : _GEN_801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_803 = 9'h123 == _GEN_9377 ? phv_data_291 : _GEN_802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_804 = 9'h124 == _GEN_9377 ? phv_data_292 : _GEN_803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_805 = 9'h125 == _GEN_9377 ? phv_data_293 : _GEN_804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_806 = 9'h126 == _GEN_9377 ? phv_data_294 : _GEN_805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_807 = 9'h127 == _GEN_9377 ? phv_data_295 : _GEN_806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_808 = 9'h128 == _GEN_9377 ? phv_data_296 : _GEN_807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_809 = 9'h129 == _GEN_9377 ? phv_data_297 : _GEN_808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_810 = 9'h12a == _GEN_9377 ? phv_data_298 : _GEN_809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_811 = 9'h12b == _GEN_9377 ? phv_data_299 : _GEN_810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_812 = 9'h12c == _GEN_9377 ? phv_data_300 : _GEN_811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_813 = 9'h12d == _GEN_9377 ? phv_data_301 : _GEN_812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_814 = 9'h12e == _GEN_9377 ? phv_data_302 : _GEN_813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_815 = 9'h12f == _GEN_9377 ? phv_data_303 : _GEN_814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_816 = 9'h130 == _GEN_9377 ? phv_data_304 : _GEN_815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_817 = 9'h131 == _GEN_9377 ? phv_data_305 : _GEN_816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_818 = 9'h132 == _GEN_9377 ? phv_data_306 : _GEN_817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_819 = 9'h133 == _GEN_9377 ? phv_data_307 : _GEN_818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_820 = 9'h134 == _GEN_9377 ? phv_data_308 : _GEN_819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_821 = 9'h135 == _GEN_9377 ? phv_data_309 : _GEN_820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_822 = 9'h136 == _GEN_9377 ? phv_data_310 : _GEN_821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_823 = 9'h137 == _GEN_9377 ? phv_data_311 : _GEN_822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_824 = 9'h138 == _GEN_9377 ? phv_data_312 : _GEN_823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_825 = 9'h139 == _GEN_9377 ? phv_data_313 : _GEN_824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_826 = 9'h13a == _GEN_9377 ? phv_data_314 : _GEN_825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_827 = 9'h13b == _GEN_9377 ? phv_data_315 : _GEN_826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_828 = 9'h13c == _GEN_9377 ? phv_data_316 : _GEN_827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_829 = 9'h13d == _GEN_9377 ? phv_data_317 : _GEN_828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_830 = 9'h13e == _GEN_9377 ? phv_data_318 : _GEN_829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_831 = 9'h13f == _GEN_9377 ? phv_data_319 : _GEN_830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_832 = 9'h140 == _GEN_9377 ? phv_data_320 : _GEN_831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_833 = 9'h141 == _GEN_9377 ? phv_data_321 : _GEN_832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_834 = 9'h142 == _GEN_9377 ? phv_data_322 : _GEN_833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_835 = 9'h143 == _GEN_9377 ? phv_data_323 : _GEN_834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_836 = 9'h144 == _GEN_9377 ? phv_data_324 : _GEN_835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_837 = 9'h145 == _GEN_9377 ? phv_data_325 : _GEN_836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_838 = 9'h146 == _GEN_9377 ? phv_data_326 : _GEN_837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_839 = 9'h147 == _GEN_9377 ? phv_data_327 : _GEN_838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_840 = 9'h148 == _GEN_9377 ? phv_data_328 : _GEN_839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_841 = 9'h149 == _GEN_9377 ? phv_data_329 : _GEN_840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_842 = 9'h14a == _GEN_9377 ? phv_data_330 : _GEN_841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_843 = 9'h14b == _GEN_9377 ? phv_data_331 : _GEN_842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_844 = 9'h14c == _GEN_9377 ? phv_data_332 : _GEN_843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_845 = 9'h14d == _GEN_9377 ? phv_data_333 : _GEN_844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_846 = 9'h14e == _GEN_9377 ? phv_data_334 : _GEN_845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_847 = 9'h14f == _GEN_9377 ? phv_data_335 : _GEN_846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_848 = 9'h150 == _GEN_9377 ? phv_data_336 : _GEN_847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_849 = 9'h151 == _GEN_9377 ? phv_data_337 : _GEN_848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_850 = 9'h152 == _GEN_9377 ? phv_data_338 : _GEN_849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_851 = 9'h153 == _GEN_9377 ? phv_data_339 : _GEN_850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_852 = 9'h154 == _GEN_9377 ? phv_data_340 : _GEN_851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_853 = 9'h155 == _GEN_9377 ? phv_data_341 : _GEN_852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_854 = 9'h156 == _GEN_9377 ? phv_data_342 : _GEN_853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_855 = 9'h157 == _GEN_9377 ? phv_data_343 : _GEN_854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_856 = 9'h158 == _GEN_9377 ? phv_data_344 : _GEN_855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_857 = 9'h159 == _GEN_9377 ? phv_data_345 : _GEN_856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_858 = 9'h15a == _GEN_9377 ? phv_data_346 : _GEN_857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_859 = 9'h15b == _GEN_9377 ? phv_data_347 : _GEN_858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_860 = 9'h15c == _GEN_9377 ? phv_data_348 : _GEN_859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_861 = 9'h15d == _GEN_9377 ? phv_data_349 : _GEN_860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_862 = 9'h15e == _GEN_9377 ? phv_data_350 : _GEN_861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_863 = 9'h15f == _GEN_9377 ? phv_data_351 : _GEN_862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_864 = 9'h160 == _GEN_9377 ? phv_data_352 : _GEN_863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_865 = 9'h161 == _GEN_9377 ? phv_data_353 : _GEN_864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_866 = 9'h162 == _GEN_9377 ? phv_data_354 : _GEN_865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_867 = 9'h163 == _GEN_9377 ? phv_data_355 : _GEN_866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_868 = 9'h164 == _GEN_9377 ? phv_data_356 : _GEN_867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_869 = 9'h165 == _GEN_9377 ? phv_data_357 : _GEN_868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_870 = 9'h166 == _GEN_9377 ? phv_data_358 : _GEN_869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_871 = 9'h167 == _GEN_9377 ? phv_data_359 : _GEN_870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_872 = 9'h168 == _GEN_9377 ? phv_data_360 : _GEN_871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_873 = 9'h169 == _GEN_9377 ? phv_data_361 : _GEN_872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_874 = 9'h16a == _GEN_9377 ? phv_data_362 : _GEN_873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_875 = 9'h16b == _GEN_9377 ? phv_data_363 : _GEN_874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_876 = 9'h16c == _GEN_9377 ? phv_data_364 : _GEN_875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_877 = 9'h16d == _GEN_9377 ? phv_data_365 : _GEN_876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_878 = 9'h16e == _GEN_9377 ? phv_data_366 : _GEN_877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_879 = 9'h16f == _GEN_9377 ? phv_data_367 : _GEN_878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_880 = 9'h170 == _GEN_9377 ? phv_data_368 : _GEN_879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_881 = 9'h171 == _GEN_9377 ? phv_data_369 : _GEN_880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_882 = 9'h172 == _GEN_9377 ? phv_data_370 : _GEN_881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_883 = 9'h173 == _GEN_9377 ? phv_data_371 : _GEN_882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_884 = 9'h174 == _GEN_9377 ? phv_data_372 : _GEN_883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_885 = 9'h175 == _GEN_9377 ? phv_data_373 : _GEN_884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_886 = 9'h176 == _GEN_9377 ? phv_data_374 : _GEN_885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_887 = 9'h177 == _GEN_9377 ? phv_data_375 : _GEN_886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_888 = 9'h178 == _GEN_9377 ? phv_data_376 : _GEN_887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_889 = 9'h179 == _GEN_9377 ? phv_data_377 : _GEN_888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_890 = 9'h17a == _GEN_9377 ? phv_data_378 : _GEN_889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_891 = 9'h17b == _GEN_9377 ? phv_data_379 : _GEN_890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_892 = 9'h17c == _GEN_9377 ? phv_data_380 : _GEN_891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_893 = 9'h17d == _GEN_9377 ? phv_data_381 : _GEN_892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_894 = 9'h17e == _GEN_9377 ? phv_data_382 : _GEN_893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_895 = 9'h17f == _GEN_9377 ? phv_data_383 : _GEN_894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_896 = 9'h180 == _GEN_9377 ? phv_data_384 : _GEN_895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_897 = 9'h181 == _GEN_9377 ? phv_data_385 : _GEN_896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_898 = 9'h182 == _GEN_9377 ? phv_data_386 : _GEN_897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_899 = 9'h183 == _GEN_9377 ? phv_data_387 : _GEN_898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_900 = 9'h184 == _GEN_9377 ? phv_data_388 : _GEN_899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_901 = 9'h185 == _GEN_9377 ? phv_data_389 : _GEN_900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_902 = 9'h186 == _GEN_9377 ? phv_data_390 : _GEN_901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_903 = 9'h187 == _GEN_9377 ? phv_data_391 : _GEN_902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_904 = 9'h188 == _GEN_9377 ? phv_data_392 : _GEN_903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_905 = 9'h189 == _GEN_9377 ? phv_data_393 : _GEN_904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_906 = 9'h18a == _GEN_9377 ? phv_data_394 : _GEN_905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_907 = 9'h18b == _GEN_9377 ? phv_data_395 : _GEN_906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_908 = 9'h18c == _GEN_9377 ? phv_data_396 : _GEN_907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_909 = 9'h18d == _GEN_9377 ? phv_data_397 : _GEN_908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_910 = 9'h18e == _GEN_9377 ? phv_data_398 : _GEN_909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_911 = 9'h18f == _GEN_9377 ? phv_data_399 : _GEN_910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_912 = 9'h190 == _GEN_9377 ? phv_data_400 : _GEN_911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_913 = 9'h191 == _GEN_9377 ? phv_data_401 : _GEN_912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_914 = 9'h192 == _GEN_9377 ? phv_data_402 : _GEN_913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_915 = 9'h193 == _GEN_9377 ? phv_data_403 : _GEN_914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_916 = 9'h194 == _GEN_9377 ? phv_data_404 : _GEN_915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_917 = 9'h195 == _GEN_9377 ? phv_data_405 : _GEN_916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_918 = 9'h196 == _GEN_9377 ? phv_data_406 : _GEN_917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_919 = 9'h197 == _GEN_9377 ? phv_data_407 : _GEN_918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_920 = 9'h198 == _GEN_9377 ? phv_data_408 : _GEN_919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_921 = 9'h199 == _GEN_9377 ? phv_data_409 : _GEN_920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_922 = 9'h19a == _GEN_9377 ? phv_data_410 : _GEN_921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_923 = 9'h19b == _GEN_9377 ? phv_data_411 : _GEN_922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_924 = 9'h19c == _GEN_9377 ? phv_data_412 : _GEN_923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_925 = 9'h19d == _GEN_9377 ? phv_data_413 : _GEN_924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_926 = 9'h19e == _GEN_9377 ? phv_data_414 : _GEN_925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_927 = 9'h19f == _GEN_9377 ? phv_data_415 : _GEN_926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_928 = 9'h1a0 == _GEN_9377 ? phv_data_416 : _GEN_927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_929 = 9'h1a1 == _GEN_9377 ? phv_data_417 : _GEN_928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_930 = 9'h1a2 == _GEN_9377 ? phv_data_418 : _GEN_929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_931 = 9'h1a3 == _GEN_9377 ? phv_data_419 : _GEN_930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_932 = 9'h1a4 == _GEN_9377 ? phv_data_420 : _GEN_931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_933 = 9'h1a5 == _GEN_9377 ? phv_data_421 : _GEN_932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_934 = 9'h1a6 == _GEN_9377 ? phv_data_422 : _GEN_933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_935 = 9'h1a7 == _GEN_9377 ? phv_data_423 : _GEN_934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_936 = 9'h1a8 == _GEN_9377 ? phv_data_424 : _GEN_935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_937 = 9'h1a9 == _GEN_9377 ? phv_data_425 : _GEN_936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_938 = 9'h1aa == _GEN_9377 ? phv_data_426 : _GEN_937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_939 = 9'h1ab == _GEN_9377 ? phv_data_427 : _GEN_938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_940 = 9'h1ac == _GEN_9377 ? phv_data_428 : _GEN_939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_941 = 9'h1ad == _GEN_9377 ? phv_data_429 : _GEN_940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_942 = 9'h1ae == _GEN_9377 ? phv_data_430 : _GEN_941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_943 = 9'h1af == _GEN_9377 ? phv_data_431 : _GEN_942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_944 = 9'h1b0 == _GEN_9377 ? phv_data_432 : _GEN_943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_945 = 9'h1b1 == _GEN_9377 ? phv_data_433 : _GEN_944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_946 = 9'h1b2 == _GEN_9377 ? phv_data_434 : _GEN_945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_947 = 9'h1b3 == _GEN_9377 ? phv_data_435 : _GEN_946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_948 = 9'h1b4 == _GEN_9377 ? phv_data_436 : _GEN_947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_949 = 9'h1b5 == _GEN_9377 ? phv_data_437 : _GEN_948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_950 = 9'h1b6 == _GEN_9377 ? phv_data_438 : _GEN_949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_951 = 9'h1b7 == _GEN_9377 ? phv_data_439 : _GEN_950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_952 = 9'h1b8 == _GEN_9377 ? phv_data_440 : _GEN_951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_953 = 9'h1b9 == _GEN_9377 ? phv_data_441 : _GEN_952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_954 = 9'h1ba == _GEN_9377 ? phv_data_442 : _GEN_953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_955 = 9'h1bb == _GEN_9377 ? phv_data_443 : _GEN_954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_956 = 9'h1bc == _GEN_9377 ? phv_data_444 : _GEN_955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_957 = 9'h1bd == _GEN_9377 ? phv_data_445 : _GEN_956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_958 = 9'h1be == _GEN_9377 ? phv_data_446 : _GEN_957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_959 = 9'h1bf == _GEN_9377 ? phv_data_447 : _GEN_958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_960 = 9'h1c0 == _GEN_9377 ? phv_data_448 : _GEN_959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_961 = 9'h1c1 == _GEN_9377 ? phv_data_449 : _GEN_960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_962 = 9'h1c2 == _GEN_9377 ? phv_data_450 : _GEN_961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_963 = 9'h1c3 == _GEN_9377 ? phv_data_451 : _GEN_962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_964 = 9'h1c4 == _GEN_9377 ? phv_data_452 : _GEN_963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_965 = 9'h1c5 == _GEN_9377 ? phv_data_453 : _GEN_964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_966 = 9'h1c6 == _GEN_9377 ? phv_data_454 : _GEN_965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_967 = 9'h1c7 == _GEN_9377 ? phv_data_455 : _GEN_966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_968 = 9'h1c8 == _GEN_9377 ? phv_data_456 : _GEN_967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_969 = 9'h1c9 == _GEN_9377 ? phv_data_457 : _GEN_968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_970 = 9'h1ca == _GEN_9377 ? phv_data_458 : _GEN_969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_971 = 9'h1cb == _GEN_9377 ? phv_data_459 : _GEN_970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_972 = 9'h1cc == _GEN_9377 ? phv_data_460 : _GEN_971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_973 = 9'h1cd == _GEN_9377 ? phv_data_461 : _GEN_972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_974 = 9'h1ce == _GEN_9377 ? phv_data_462 : _GEN_973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_975 = 9'h1cf == _GEN_9377 ? phv_data_463 : _GEN_974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_976 = 9'h1d0 == _GEN_9377 ? phv_data_464 : _GEN_975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_977 = 9'h1d1 == _GEN_9377 ? phv_data_465 : _GEN_976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_978 = 9'h1d2 == _GEN_9377 ? phv_data_466 : _GEN_977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_979 = 9'h1d3 == _GEN_9377 ? phv_data_467 : _GEN_978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_980 = 9'h1d4 == _GEN_9377 ? phv_data_468 : _GEN_979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_981 = 9'h1d5 == _GEN_9377 ? phv_data_469 : _GEN_980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_982 = 9'h1d6 == _GEN_9377 ? phv_data_470 : _GEN_981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_983 = 9'h1d7 == _GEN_9377 ? phv_data_471 : _GEN_982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_984 = 9'h1d8 == _GEN_9377 ? phv_data_472 : _GEN_983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_985 = 9'h1d9 == _GEN_9377 ? phv_data_473 : _GEN_984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_986 = 9'h1da == _GEN_9377 ? phv_data_474 : _GEN_985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_987 = 9'h1db == _GEN_9377 ? phv_data_475 : _GEN_986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_988 = 9'h1dc == _GEN_9377 ? phv_data_476 : _GEN_987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_989 = 9'h1dd == _GEN_9377 ? phv_data_477 : _GEN_988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_990 = 9'h1de == _GEN_9377 ? phv_data_478 : _GEN_989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_991 = 9'h1df == _GEN_9377 ? phv_data_479 : _GEN_990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_992 = 9'h1e0 == _GEN_9377 ? phv_data_480 : _GEN_991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_993 = 9'h1e1 == _GEN_9377 ? phv_data_481 : _GEN_992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_994 = 9'h1e2 == _GEN_9377 ? phv_data_482 : _GEN_993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_995 = 9'h1e3 == _GEN_9377 ? phv_data_483 : _GEN_994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_996 = 9'h1e4 == _GEN_9377 ? phv_data_484 : _GEN_995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_997 = 9'h1e5 == _GEN_9377 ? phv_data_485 : _GEN_996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_998 = 9'h1e6 == _GEN_9377 ? phv_data_486 : _GEN_997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_999 = 9'h1e7 == _GEN_9377 ? phv_data_487 : _GEN_998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1000 = 9'h1e8 == _GEN_9377 ? phv_data_488 : _GEN_999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1001 = 9'h1e9 == _GEN_9377 ? phv_data_489 : _GEN_1000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1002 = 9'h1ea == _GEN_9377 ? phv_data_490 : _GEN_1001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1003 = 9'h1eb == _GEN_9377 ? phv_data_491 : _GEN_1002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1004 = 9'h1ec == _GEN_9377 ? phv_data_492 : _GEN_1003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1005 = 9'h1ed == _GEN_9377 ? phv_data_493 : _GEN_1004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1006 = 9'h1ee == _GEN_9377 ? phv_data_494 : _GEN_1005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1007 = 9'h1ef == _GEN_9377 ? phv_data_495 : _GEN_1006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1008 = 9'h1f0 == _GEN_9377 ? phv_data_496 : _GEN_1007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1009 = 9'h1f1 == _GEN_9377 ? phv_data_497 : _GEN_1008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1010 = 9'h1f2 == _GEN_9377 ? phv_data_498 : _GEN_1009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1011 = 9'h1f3 == _GEN_9377 ? phv_data_499 : _GEN_1010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1012 = 9'h1f4 == _GEN_9377 ? phv_data_500 : _GEN_1011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1013 = 9'h1f5 == _GEN_9377 ? phv_data_501 : _GEN_1012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1014 = 9'h1f6 == _GEN_9377 ? phv_data_502 : _GEN_1013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1015 = 9'h1f7 == _GEN_9377 ? phv_data_503 : _GEN_1014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1016 = 9'h1f8 == _GEN_9377 ? phv_data_504 : _GEN_1015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1017 = 9'h1f9 == _GEN_9377 ? phv_data_505 : _GEN_1016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1018 = 9'h1fa == _GEN_9377 ? phv_data_506 : _GEN_1017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1019 = 9'h1fb == _GEN_9377 ? phv_data_507 : _GEN_1018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1020 = 9'h1fc == _GEN_9377 ? phv_data_508 : _GEN_1019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1021 = 9'h1fd == _GEN_9377 ? phv_data_509 : _GEN_1020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1022 = 9'h1fe == _GEN_9377 ? phv_data_510 : _GEN_1021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__2 = 9'h1ff == _GEN_9377 ? phv_data_511 : _GEN_1022; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask__2 = 2'h1 >= offset_0[1:0] & (2'h1 < ending | ending == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_2 = {total_offset_hi,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1025 = 8'h1 == total_offset_2 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1026 = 8'h2 == total_offset_2 ? phv_data_2 : _GEN_1025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1027 = 8'h3 == total_offset_2 ? phv_data_3 : _GEN_1026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1028 = 8'h4 == total_offset_2 ? phv_data_4 : _GEN_1027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1029 = 8'h5 == total_offset_2 ? phv_data_5 : _GEN_1028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1030 = 8'h6 == total_offset_2 ? phv_data_6 : _GEN_1029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1031 = 8'h7 == total_offset_2 ? phv_data_7 : _GEN_1030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1032 = 8'h8 == total_offset_2 ? phv_data_8 : _GEN_1031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1033 = 8'h9 == total_offset_2 ? phv_data_9 : _GEN_1032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1034 = 8'ha == total_offset_2 ? phv_data_10 : _GEN_1033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1035 = 8'hb == total_offset_2 ? phv_data_11 : _GEN_1034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1036 = 8'hc == total_offset_2 ? phv_data_12 : _GEN_1035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1037 = 8'hd == total_offset_2 ? phv_data_13 : _GEN_1036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1038 = 8'he == total_offset_2 ? phv_data_14 : _GEN_1037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1039 = 8'hf == total_offset_2 ? phv_data_15 : _GEN_1038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1040 = 8'h10 == total_offset_2 ? phv_data_16 : _GEN_1039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1041 = 8'h11 == total_offset_2 ? phv_data_17 : _GEN_1040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1042 = 8'h12 == total_offset_2 ? phv_data_18 : _GEN_1041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1043 = 8'h13 == total_offset_2 ? phv_data_19 : _GEN_1042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1044 = 8'h14 == total_offset_2 ? phv_data_20 : _GEN_1043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1045 = 8'h15 == total_offset_2 ? phv_data_21 : _GEN_1044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1046 = 8'h16 == total_offset_2 ? phv_data_22 : _GEN_1045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1047 = 8'h17 == total_offset_2 ? phv_data_23 : _GEN_1046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1048 = 8'h18 == total_offset_2 ? phv_data_24 : _GEN_1047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1049 = 8'h19 == total_offset_2 ? phv_data_25 : _GEN_1048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1050 = 8'h1a == total_offset_2 ? phv_data_26 : _GEN_1049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1051 = 8'h1b == total_offset_2 ? phv_data_27 : _GEN_1050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1052 = 8'h1c == total_offset_2 ? phv_data_28 : _GEN_1051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1053 = 8'h1d == total_offset_2 ? phv_data_29 : _GEN_1052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1054 = 8'h1e == total_offset_2 ? phv_data_30 : _GEN_1053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1055 = 8'h1f == total_offset_2 ? phv_data_31 : _GEN_1054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1056 = 8'h20 == total_offset_2 ? phv_data_32 : _GEN_1055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1057 = 8'h21 == total_offset_2 ? phv_data_33 : _GEN_1056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1058 = 8'h22 == total_offset_2 ? phv_data_34 : _GEN_1057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1059 = 8'h23 == total_offset_2 ? phv_data_35 : _GEN_1058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1060 = 8'h24 == total_offset_2 ? phv_data_36 : _GEN_1059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1061 = 8'h25 == total_offset_2 ? phv_data_37 : _GEN_1060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1062 = 8'h26 == total_offset_2 ? phv_data_38 : _GEN_1061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1063 = 8'h27 == total_offset_2 ? phv_data_39 : _GEN_1062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1064 = 8'h28 == total_offset_2 ? phv_data_40 : _GEN_1063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1065 = 8'h29 == total_offset_2 ? phv_data_41 : _GEN_1064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1066 = 8'h2a == total_offset_2 ? phv_data_42 : _GEN_1065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1067 = 8'h2b == total_offset_2 ? phv_data_43 : _GEN_1066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1068 = 8'h2c == total_offset_2 ? phv_data_44 : _GEN_1067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1069 = 8'h2d == total_offset_2 ? phv_data_45 : _GEN_1068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1070 = 8'h2e == total_offset_2 ? phv_data_46 : _GEN_1069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1071 = 8'h2f == total_offset_2 ? phv_data_47 : _GEN_1070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1072 = 8'h30 == total_offset_2 ? phv_data_48 : _GEN_1071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1073 = 8'h31 == total_offset_2 ? phv_data_49 : _GEN_1072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1074 = 8'h32 == total_offset_2 ? phv_data_50 : _GEN_1073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1075 = 8'h33 == total_offset_2 ? phv_data_51 : _GEN_1074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1076 = 8'h34 == total_offset_2 ? phv_data_52 : _GEN_1075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1077 = 8'h35 == total_offset_2 ? phv_data_53 : _GEN_1076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1078 = 8'h36 == total_offset_2 ? phv_data_54 : _GEN_1077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1079 = 8'h37 == total_offset_2 ? phv_data_55 : _GEN_1078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1080 = 8'h38 == total_offset_2 ? phv_data_56 : _GEN_1079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1081 = 8'h39 == total_offset_2 ? phv_data_57 : _GEN_1080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1082 = 8'h3a == total_offset_2 ? phv_data_58 : _GEN_1081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1083 = 8'h3b == total_offset_2 ? phv_data_59 : _GEN_1082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1084 = 8'h3c == total_offset_2 ? phv_data_60 : _GEN_1083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1085 = 8'h3d == total_offset_2 ? phv_data_61 : _GEN_1084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1086 = 8'h3e == total_offset_2 ? phv_data_62 : _GEN_1085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1087 = 8'h3f == total_offset_2 ? phv_data_63 : _GEN_1086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1088 = 8'h40 == total_offset_2 ? phv_data_64 : _GEN_1087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1089 = 8'h41 == total_offset_2 ? phv_data_65 : _GEN_1088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1090 = 8'h42 == total_offset_2 ? phv_data_66 : _GEN_1089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1091 = 8'h43 == total_offset_2 ? phv_data_67 : _GEN_1090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1092 = 8'h44 == total_offset_2 ? phv_data_68 : _GEN_1091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1093 = 8'h45 == total_offset_2 ? phv_data_69 : _GEN_1092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1094 = 8'h46 == total_offset_2 ? phv_data_70 : _GEN_1093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1095 = 8'h47 == total_offset_2 ? phv_data_71 : _GEN_1094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1096 = 8'h48 == total_offset_2 ? phv_data_72 : _GEN_1095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1097 = 8'h49 == total_offset_2 ? phv_data_73 : _GEN_1096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1098 = 8'h4a == total_offset_2 ? phv_data_74 : _GEN_1097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1099 = 8'h4b == total_offset_2 ? phv_data_75 : _GEN_1098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1100 = 8'h4c == total_offset_2 ? phv_data_76 : _GEN_1099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1101 = 8'h4d == total_offset_2 ? phv_data_77 : _GEN_1100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1102 = 8'h4e == total_offset_2 ? phv_data_78 : _GEN_1101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1103 = 8'h4f == total_offset_2 ? phv_data_79 : _GEN_1102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1104 = 8'h50 == total_offset_2 ? phv_data_80 : _GEN_1103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1105 = 8'h51 == total_offset_2 ? phv_data_81 : _GEN_1104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1106 = 8'h52 == total_offset_2 ? phv_data_82 : _GEN_1105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1107 = 8'h53 == total_offset_2 ? phv_data_83 : _GEN_1106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1108 = 8'h54 == total_offset_2 ? phv_data_84 : _GEN_1107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1109 = 8'h55 == total_offset_2 ? phv_data_85 : _GEN_1108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1110 = 8'h56 == total_offset_2 ? phv_data_86 : _GEN_1109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1111 = 8'h57 == total_offset_2 ? phv_data_87 : _GEN_1110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1112 = 8'h58 == total_offset_2 ? phv_data_88 : _GEN_1111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1113 = 8'h59 == total_offset_2 ? phv_data_89 : _GEN_1112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1114 = 8'h5a == total_offset_2 ? phv_data_90 : _GEN_1113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1115 = 8'h5b == total_offset_2 ? phv_data_91 : _GEN_1114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1116 = 8'h5c == total_offset_2 ? phv_data_92 : _GEN_1115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1117 = 8'h5d == total_offset_2 ? phv_data_93 : _GEN_1116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1118 = 8'h5e == total_offset_2 ? phv_data_94 : _GEN_1117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1119 = 8'h5f == total_offset_2 ? phv_data_95 : _GEN_1118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1120 = 8'h60 == total_offset_2 ? phv_data_96 : _GEN_1119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1121 = 8'h61 == total_offset_2 ? phv_data_97 : _GEN_1120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1122 = 8'h62 == total_offset_2 ? phv_data_98 : _GEN_1121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1123 = 8'h63 == total_offset_2 ? phv_data_99 : _GEN_1122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1124 = 8'h64 == total_offset_2 ? phv_data_100 : _GEN_1123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1125 = 8'h65 == total_offset_2 ? phv_data_101 : _GEN_1124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1126 = 8'h66 == total_offset_2 ? phv_data_102 : _GEN_1125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1127 = 8'h67 == total_offset_2 ? phv_data_103 : _GEN_1126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1128 = 8'h68 == total_offset_2 ? phv_data_104 : _GEN_1127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1129 = 8'h69 == total_offset_2 ? phv_data_105 : _GEN_1128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1130 = 8'h6a == total_offset_2 ? phv_data_106 : _GEN_1129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1131 = 8'h6b == total_offset_2 ? phv_data_107 : _GEN_1130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1132 = 8'h6c == total_offset_2 ? phv_data_108 : _GEN_1131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1133 = 8'h6d == total_offset_2 ? phv_data_109 : _GEN_1132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1134 = 8'h6e == total_offset_2 ? phv_data_110 : _GEN_1133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1135 = 8'h6f == total_offset_2 ? phv_data_111 : _GEN_1134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1136 = 8'h70 == total_offset_2 ? phv_data_112 : _GEN_1135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1137 = 8'h71 == total_offset_2 ? phv_data_113 : _GEN_1136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1138 = 8'h72 == total_offset_2 ? phv_data_114 : _GEN_1137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1139 = 8'h73 == total_offset_2 ? phv_data_115 : _GEN_1138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1140 = 8'h74 == total_offset_2 ? phv_data_116 : _GEN_1139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1141 = 8'h75 == total_offset_2 ? phv_data_117 : _GEN_1140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1142 = 8'h76 == total_offset_2 ? phv_data_118 : _GEN_1141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1143 = 8'h77 == total_offset_2 ? phv_data_119 : _GEN_1142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1144 = 8'h78 == total_offset_2 ? phv_data_120 : _GEN_1143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1145 = 8'h79 == total_offset_2 ? phv_data_121 : _GEN_1144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1146 = 8'h7a == total_offset_2 ? phv_data_122 : _GEN_1145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1147 = 8'h7b == total_offset_2 ? phv_data_123 : _GEN_1146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1148 = 8'h7c == total_offset_2 ? phv_data_124 : _GEN_1147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1149 = 8'h7d == total_offset_2 ? phv_data_125 : _GEN_1148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1150 = 8'h7e == total_offset_2 ? phv_data_126 : _GEN_1149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1151 = 8'h7f == total_offset_2 ? phv_data_127 : _GEN_1150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1152 = 8'h80 == total_offset_2 ? phv_data_128 : _GEN_1151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1153 = 8'h81 == total_offset_2 ? phv_data_129 : _GEN_1152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1154 = 8'h82 == total_offset_2 ? phv_data_130 : _GEN_1153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1155 = 8'h83 == total_offset_2 ? phv_data_131 : _GEN_1154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1156 = 8'h84 == total_offset_2 ? phv_data_132 : _GEN_1155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1157 = 8'h85 == total_offset_2 ? phv_data_133 : _GEN_1156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1158 = 8'h86 == total_offset_2 ? phv_data_134 : _GEN_1157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1159 = 8'h87 == total_offset_2 ? phv_data_135 : _GEN_1158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1160 = 8'h88 == total_offset_2 ? phv_data_136 : _GEN_1159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1161 = 8'h89 == total_offset_2 ? phv_data_137 : _GEN_1160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1162 = 8'h8a == total_offset_2 ? phv_data_138 : _GEN_1161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1163 = 8'h8b == total_offset_2 ? phv_data_139 : _GEN_1162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1164 = 8'h8c == total_offset_2 ? phv_data_140 : _GEN_1163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1165 = 8'h8d == total_offset_2 ? phv_data_141 : _GEN_1164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1166 = 8'h8e == total_offset_2 ? phv_data_142 : _GEN_1165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1167 = 8'h8f == total_offset_2 ? phv_data_143 : _GEN_1166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1168 = 8'h90 == total_offset_2 ? phv_data_144 : _GEN_1167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1169 = 8'h91 == total_offset_2 ? phv_data_145 : _GEN_1168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1170 = 8'h92 == total_offset_2 ? phv_data_146 : _GEN_1169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1171 = 8'h93 == total_offset_2 ? phv_data_147 : _GEN_1170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1172 = 8'h94 == total_offset_2 ? phv_data_148 : _GEN_1171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1173 = 8'h95 == total_offset_2 ? phv_data_149 : _GEN_1172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1174 = 8'h96 == total_offset_2 ? phv_data_150 : _GEN_1173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1175 = 8'h97 == total_offset_2 ? phv_data_151 : _GEN_1174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1176 = 8'h98 == total_offset_2 ? phv_data_152 : _GEN_1175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1177 = 8'h99 == total_offset_2 ? phv_data_153 : _GEN_1176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1178 = 8'h9a == total_offset_2 ? phv_data_154 : _GEN_1177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1179 = 8'h9b == total_offset_2 ? phv_data_155 : _GEN_1178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1180 = 8'h9c == total_offset_2 ? phv_data_156 : _GEN_1179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1181 = 8'h9d == total_offset_2 ? phv_data_157 : _GEN_1180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1182 = 8'h9e == total_offset_2 ? phv_data_158 : _GEN_1181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1183 = 8'h9f == total_offset_2 ? phv_data_159 : _GEN_1182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1184 = 8'ha0 == total_offset_2 ? phv_data_160 : _GEN_1183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1185 = 8'ha1 == total_offset_2 ? phv_data_161 : _GEN_1184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1186 = 8'ha2 == total_offset_2 ? phv_data_162 : _GEN_1185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1187 = 8'ha3 == total_offset_2 ? phv_data_163 : _GEN_1186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1188 = 8'ha4 == total_offset_2 ? phv_data_164 : _GEN_1187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1189 = 8'ha5 == total_offset_2 ? phv_data_165 : _GEN_1188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1190 = 8'ha6 == total_offset_2 ? phv_data_166 : _GEN_1189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1191 = 8'ha7 == total_offset_2 ? phv_data_167 : _GEN_1190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1192 = 8'ha8 == total_offset_2 ? phv_data_168 : _GEN_1191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1193 = 8'ha9 == total_offset_2 ? phv_data_169 : _GEN_1192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1194 = 8'haa == total_offset_2 ? phv_data_170 : _GEN_1193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1195 = 8'hab == total_offset_2 ? phv_data_171 : _GEN_1194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1196 = 8'hac == total_offset_2 ? phv_data_172 : _GEN_1195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1197 = 8'had == total_offset_2 ? phv_data_173 : _GEN_1196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1198 = 8'hae == total_offset_2 ? phv_data_174 : _GEN_1197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1199 = 8'haf == total_offset_2 ? phv_data_175 : _GEN_1198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1200 = 8'hb0 == total_offset_2 ? phv_data_176 : _GEN_1199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1201 = 8'hb1 == total_offset_2 ? phv_data_177 : _GEN_1200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1202 = 8'hb2 == total_offset_2 ? phv_data_178 : _GEN_1201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1203 = 8'hb3 == total_offset_2 ? phv_data_179 : _GEN_1202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1204 = 8'hb4 == total_offset_2 ? phv_data_180 : _GEN_1203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1205 = 8'hb5 == total_offset_2 ? phv_data_181 : _GEN_1204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1206 = 8'hb6 == total_offset_2 ? phv_data_182 : _GEN_1205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1207 = 8'hb7 == total_offset_2 ? phv_data_183 : _GEN_1206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1208 = 8'hb8 == total_offset_2 ? phv_data_184 : _GEN_1207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1209 = 8'hb9 == total_offset_2 ? phv_data_185 : _GEN_1208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1210 = 8'hba == total_offset_2 ? phv_data_186 : _GEN_1209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1211 = 8'hbb == total_offset_2 ? phv_data_187 : _GEN_1210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1212 = 8'hbc == total_offset_2 ? phv_data_188 : _GEN_1211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1213 = 8'hbd == total_offset_2 ? phv_data_189 : _GEN_1212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1214 = 8'hbe == total_offset_2 ? phv_data_190 : _GEN_1213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1215 = 8'hbf == total_offset_2 ? phv_data_191 : _GEN_1214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1216 = 8'hc0 == total_offset_2 ? phv_data_192 : _GEN_1215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1217 = 8'hc1 == total_offset_2 ? phv_data_193 : _GEN_1216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1218 = 8'hc2 == total_offset_2 ? phv_data_194 : _GEN_1217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1219 = 8'hc3 == total_offset_2 ? phv_data_195 : _GEN_1218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1220 = 8'hc4 == total_offset_2 ? phv_data_196 : _GEN_1219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1221 = 8'hc5 == total_offset_2 ? phv_data_197 : _GEN_1220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1222 = 8'hc6 == total_offset_2 ? phv_data_198 : _GEN_1221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1223 = 8'hc7 == total_offset_2 ? phv_data_199 : _GEN_1222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1224 = 8'hc8 == total_offset_2 ? phv_data_200 : _GEN_1223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1225 = 8'hc9 == total_offset_2 ? phv_data_201 : _GEN_1224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1226 = 8'hca == total_offset_2 ? phv_data_202 : _GEN_1225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1227 = 8'hcb == total_offset_2 ? phv_data_203 : _GEN_1226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1228 = 8'hcc == total_offset_2 ? phv_data_204 : _GEN_1227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1229 = 8'hcd == total_offset_2 ? phv_data_205 : _GEN_1228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1230 = 8'hce == total_offset_2 ? phv_data_206 : _GEN_1229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1231 = 8'hcf == total_offset_2 ? phv_data_207 : _GEN_1230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1232 = 8'hd0 == total_offset_2 ? phv_data_208 : _GEN_1231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1233 = 8'hd1 == total_offset_2 ? phv_data_209 : _GEN_1232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1234 = 8'hd2 == total_offset_2 ? phv_data_210 : _GEN_1233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1235 = 8'hd3 == total_offset_2 ? phv_data_211 : _GEN_1234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1236 = 8'hd4 == total_offset_2 ? phv_data_212 : _GEN_1235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1237 = 8'hd5 == total_offset_2 ? phv_data_213 : _GEN_1236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1238 = 8'hd6 == total_offset_2 ? phv_data_214 : _GEN_1237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1239 = 8'hd7 == total_offset_2 ? phv_data_215 : _GEN_1238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1240 = 8'hd8 == total_offset_2 ? phv_data_216 : _GEN_1239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1241 = 8'hd9 == total_offset_2 ? phv_data_217 : _GEN_1240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1242 = 8'hda == total_offset_2 ? phv_data_218 : _GEN_1241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1243 = 8'hdb == total_offset_2 ? phv_data_219 : _GEN_1242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1244 = 8'hdc == total_offset_2 ? phv_data_220 : _GEN_1243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1245 = 8'hdd == total_offset_2 ? phv_data_221 : _GEN_1244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1246 = 8'hde == total_offset_2 ? phv_data_222 : _GEN_1245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1247 = 8'hdf == total_offset_2 ? phv_data_223 : _GEN_1246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1248 = 8'he0 == total_offset_2 ? phv_data_224 : _GEN_1247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1249 = 8'he1 == total_offset_2 ? phv_data_225 : _GEN_1248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1250 = 8'he2 == total_offset_2 ? phv_data_226 : _GEN_1249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1251 = 8'he3 == total_offset_2 ? phv_data_227 : _GEN_1250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1252 = 8'he4 == total_offset_2 ? phv_data_228 : _GEN_1251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1253 = 8'he5 == total_offset_2 ? phv_data_229 : _GEN_1252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1254 = 8'he6 == total_offset_2 ? phv_data_230 : _GEN_1253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1255 = 8'he7 == total_offset_2 ? phv_data_231 : _GEN_1254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1256 = 8'he8 == total_offset_2 ? phv_data_232 : _GEN_1255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1257 = 8'he9 == total_offset_2 ? phv_data_233 : _GEN_1256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1258 = 8'hea == total_offset_2 ? phv_data_234 : _GEN_1257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1259 = 8'heb == total_offset_2 ? phv_data_235 : _GEN_1258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1260 = 8'hec == total_offset_2 ? phv_data_236 : _GEN_1259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1261 = 8'hed == total_offset_2 ? phv_data_237 : _GEN_1260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1262 = 8'hee == total_offset_2 ? phv_data_238 : _GEN_1261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1263 = 8'hef == total_offset_2 ? phv_data_239 : _GEN_1262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1264 = 8'hf0 == total_offset_2 ? phv_data_240 : _GEN_1263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1265 = 8'hf1 == total_offset_2 ? phv_data_241 : _GEN_1264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1266 = 8'hf2 == total_offset_2 ? phv_data_242 : _GEN_1265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1267 = 8'hf3 == total_offset_2 ? phv_data_243 : _GEN_1266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1268 = 8'hf4 == total_offset_2 ? phv_data_244 : _GEN_1267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1269 = 8'hf5 == total_offset_2 ? phv_data_245 : _GEN_1268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1270 = 8'hf6 == total_offset_2 ? phv_data_246 : _GEN_1269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1271 = 8'hf7 == total_offset_2 ? phv_data_247 : _GEN_1270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1272 = 8'hf8 == total_offset_2 ? phv_data_248 : _GEN_1271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1273 = 8'hf9 == total_offset_2 ? phv_data_249 : _GEN_1272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1274 = 8'hfa == total_offset_2 ? phv_data_250 : _GEN_1273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1275 = 8'hfb == total_offset_2 ? phv_data_251 : _GEN_1274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1276 = 8'hfc == total_offset_2 ? phv_data_252 : _GEN_1275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1277 = 8'hfd == total_offset_2 ? phv_data_253 : _GEN_1276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1278 = 8'hfe == total_offset_2 ? phv_data_254 : _GEN_1277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1279 = 8'hff == total_offset_2 ? phv_data_255 : _GEN_1278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_9633 = {{1'd0}, total_offset_2}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1280 = 9'h100 == _GEN_9633 ? phv_data_256 : _GEN_1279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1281 = 9'h101 == _GEN_9633 ? phv_data_257 : _GEN_1280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1282 = 9'h102 == _GEN_9633 ? phv_data_258 : _GEN_1281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1283 = 9'h103 == _GEN_9633 ? phv_data_259 : _GEN_1282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1284 = 9'h104 == _GEN_9633 ? phv_data_260 : _GEN_1283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1285 = 9'h105 == _GEN_9633 ? phv_data_261 : _GEN_1284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1286 = 9'h106 == _GEN_9633 ? phv_data_262 : _GEN_1285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1287 = 9'h107 == _GEN_9633 ? phv_data_263 : _GEN_1286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1288 = 9'h108 == _GEN_9633 ? phv_data_264 : _GEN_1287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1289 = 9'h109 == _GEN_9633 ? phv_data_265 : _GEN_1288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1290 = 9'h10a == _GEN_9633 ? phv_data_266 : _GEN_1289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1291 = 9'h10b == _GEN_9633 ? phv_data_267 : _GEN_1290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1292 = 9'h10c == _GEN_9633 ? phv_data_268 : _GEN_1291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1293 = 9'h10d == _GEN_9633 ? phv_data_269 : _GEN_1292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1294 = 9'h10e == _GEN_9633 ? phv_data_270 : _GEN_1293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1295 = 9'h10f == _GEN_9633 ? phv_data_271 : _GEN_1294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1296 = 9'h110 == _GEN_9633 ? phv_data_272 : _GEN_1295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1297 = 9'h111 == _GEN_9633 ? phv_data_273 : _GEN_1296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1298 = 9'h112 == _GEN_9633 ? phv_data_274 : _GEN_1297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1299 = 9'h113 == _GEN_9633 ? phv_data_275 : _GEN_1298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1300 = 9'h114 == _GEN_9633 ? phv_data_276 : _GEN_1299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1301 = 9'h115 == _GEN_9633 ? phv_data_277 : _GEN_1300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1302 = 9'h116 == _GEN_9633 ? phv_data_278 : _GEN_1301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1303 = 9'h117 == _GEN_9633 ? phv_data_279 : _GEN_1302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1304 = 9'h118 == _GEN_9633 ? phv_data_280 : _GEN_1303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1305 = 9'h119 == _GEN_9633 ? phv_data_281 : _GEN_1304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1306 = 9'h11a == _GEN_9633 ? phv_data_282 : _GEN_1305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1307 = 9'h11b == _GEN_9633 ? phv_data_283 : _GEN_1306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1308 = 9'h11c == _GEN_9633 ? phv_data_284 : _GEN_1307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1309 = 9'h11d == _GEN_9633 ? phv_data_285 : _GEN_1308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1310 = 9'h11e == _GEN_9633 ? phv_data_286 : _GEN_1309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1311 = 9'h11f == _GEN_9633 ? phv_data_287 : _GEN_1310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1312 = 9'h120 == _GEN_9633 ? phv_data_288 : _GEN_1311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1313 = 9'h121 == _GEN_9633 ? phv_data_289 : _GEN_1312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1314 = 9'h122 == _GEN_9633 ? phv_data_290 : _GEN_1313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1315 = 9'h123 == _GEN_9633 ? phv_data_291 : _GEN_1314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1316 = 9'h124 == _GEN_9633 ? phv_data_292 : _GEN_1315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1317 = 9'h125 == _GEN_9633 ? phv_data_293 : _GEN_1316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1318 = 9'h126 == _GEN_9633 ? phv_data_294 : _GEN_1317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1319 = 9'h127 == _GEN_9633 ? phv_data_295 : _GEN_1318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1320 = 9'h128 == _GEN_9633 ? phv_data_296 : _GEN_1319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1321 = 9'h129 == _GEN_9633 ? phv_data_297 : _GEN_1320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1322 = 9'h12a == _GEN_9633 ? phv_data_298 : _GEN_1321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1323 = 9'h12b == _GEN_9633 ? phv_data_299 : _GEN_1322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1324 = 9'h12c == _GEN_9633 ? phv_data_300 : _GEN_1323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1325 = 9'h12d == _GEN_9633 ? phv_data_301 : _GEN_1324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1326 = 9'h12e == _GEN_9633 ? phv_data_302 : _GEN_1325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1327 = 9'h12f == _GEN_9633 ? phv_data_303 : _GEN_1326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1328 = 9'h130 == _GEN_9633 ? phv_data_304 : _GEN_1327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1329 = 9'h131 == _GEN_9633 ? phv_data_305 : _GEN_1328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1330 = 9'h132 == _GEN_9633 ? phv_data_306 : _GEN_1329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1331 = 9'h133 == _GEN_9633 ? phv_data_307 : _GEN_1330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1332 = 9'h134 == _GEN_9633 ? phv_data_308 : _GEN_1331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1333 = 9'h135 == _GEN_9633 ? phv_data_309 : _GEN_1332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1334 = 9'h136 == _GEN_9633 ? phv_data_310 : _GEN_1333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1335 = 9'h137 == _GEN_9633 ? phv_data_311 : _GEN_1334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1336 = 9'h138 == _GEN_9633 ? phv_data_312 : _GEN_1335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1337 = 9'h139 == _GEN_9633 ? phv_data_313 : _GEN_1336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1338 = 9'h13a == _GEN_9633 ? phv_data_314 : _GEN_1337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1339 = 9'h13b == _GEN_9633 ? phv_data_315 : _GEN_1338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1340 = 9'h13c == _GEN_9633 ? phv_data_316 : _GEN_1339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1341 = 9'h13d == _GEN_9633 ? phv_data_317 : _GEN_1340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1342 = 9'h13e == _GEN_9633 ? phv_data_318 : _GEN_1341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1343 = 9'h13f == _GEN_9633 ? phv_data_319 : _GEN_1342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1344 = 9'h140 == _GEN_9633 ? phv_data_320 : _GEN_1343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1345 = 9'h141 == _GEN_9633 ? phv_data_321 : _GEN_1344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1346 = 9'h142 == _GEN_9633 ? phv_data_322 : _GEN_1345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1347 = 9'h143 == _GEN_9633 ? phv_data_323 : _GEN_1346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1348 = 9'h144 == _GEN_9633 ? phv_data_324 : _GEN_1347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1349 = 9'h145 == _GEN_9633 ? phv_data_325 : _GEN_1348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1350 = 9'h146 == _GEN_9633 ? phv_data_326 : _GEN_1349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1351 = 9'h147 == _GEN_9633 ? phv_data_327 : _GEN_1350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1352 = 9'h148 == _GEN_9633 ? phv_data_328 : _GEN_1351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1353 = 9'h149 == _GEN_9633 ? phv_data_329 : _GEN_1352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1354 = 9'h14a == _GEN_9633 ? phv_data_330 : _GEN_1353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1355 = 9'h14b == _GEN_9633 ? phv_data_331 : _GEN_1354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1356 = 9'h14c == _GEN_9633 ? phv_data_332 : _GEN_1355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1357 = 9'h14d == _GEN_9633 ? phv_data_333 : _GEN_1356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1358 = 9'h14e == _GEN_9633 ? phv_data_334 : _GEN_1357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1359 = 9'h14f == _GEN_9633 ? phv_data_335 : _GEN_1358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1360 = 9'h150 == _GEN_9633 ? phv_data_336 : _GEN_1359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1361 = 9'h151 == _GEN_9633 ? phv_data_337 : _GEN_1360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1362 = 9'h152 == _GEN_9633 ? phv_data_338 : _GEN_1361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1363 = 9'h153 == _GEN_9633 ? phv_data_339 : _GEN_1362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1364 = 9'h154 == _GEN_9633 ? phv_data_340 : _GEN_1363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1365 = 9'h155 == _GEN_9633 ? phv_data_341 : _GEN_1364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1366 = 9'h156 == _GEN_9633 ? phv_data_342 : _GEN_1365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1367 = 9'h157 == _GEN_9633 ? phv_data_343 : _GEN_1366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1368 = 9'h158 == _GEN_9633 ? phv_data_344 : _GEN_1367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1369 = 9'h159 == _GEN_9633 ? phv_data_345 : _GEN_1368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1370 = 9'h15a == _GEN_9633 ? phv_data_346 : _GEN_1369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1371 = 9'h15b == _GEN_9633 ? phv_data_347 : _GEN_1370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1372 = 9'h15c == _GEN_9633 ? phv_data_348 : _GEN_1371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1373 = 9'h15d == _GEN_9633 ? phv_data_349 : _GEN_1372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1374 = 9'h15e == _GEN_9633 ? phv_data_350 : _GEN_1373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1375 = 9'h15f == _GEN_9633 ? phv_data_351 : _GEN_1374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1376 = 9'h160 == _GEN_9633 ? phv_data_352 : _GEN_1375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1377 = 9'h161 == _GEN_9633 ? phv_data_353 : _GEN_1376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1378 = 9'h162 == _GEN_9633 ? phv_data_354 : _GEN_1377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1379 = 9'h163 == _GEN_9633 ? phv_data_355 : _GEN_1378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1380 = 9'h164 == _GEN_9633 ? phv_data_356 : _GEN_1379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1381 = 9'h165 == _GEN_9633 ? phv_data_357 : _GEN_1380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1382 = 9'h166 == _GEN_9633 ? phv_data_358 : _GEN_1381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1383 = 9'h167 == _GEN_9633 ? phv_data_359 : _GEN_1382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1384 = 9'h168 == _GEN_9633 ? phv_data_360 : _GEN_1383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1385 = 9'h169 == _GEN_9633 ? phv_data_361 : _GEN_1384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1386 = 9'h16a == _GEN_9633 ? phv_data_362 : _GEN_1385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1387 = 9'h16b == _GEN_9633 ? phv_data_363 : _GEN_1386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1388 = 9'h16c == _GEN_9633 ? phv_data_364 : _GEN_1387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1389 = 9'h16d == _GEN_9633 ? phv_data_365 : _GEN_1388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1390 = 9'h16e == _GEN_9633 ? phv_data_366 : _GEN_1389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1391 = 9'h16f == _GEN_9633 ? phv_data_367 : _GEN_1390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1392 = 9'h170 == _GEN_9633 ? phv_data_368 : _GEN_1391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1393 = 9'h171 == _GEN_9633 ? phv_data_369 : _GEN_1392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1394 = 9'h172 == _GEN_9633 ? phv_data_370 : _GEN_1393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1395 = 9'h173 == _GEN_9633 ? phv_data_371 : _GEN_1394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1396 = 9'h174 == _GEN_9633 ? phv_data_372 : _GEN_1395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1397 = 9'h175 == _GEN_9633 ? phv_data_373 : _GEN_1396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1398 = 9'h176 == _GEN_9633 ? phv_data_374 : _GEN_1397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1399 = 9'h177 == _GEN_9633 ? phv_data_375 : _GEN_1398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1400 = 9'h178 == _GEN_9633 ? phv_data_376 : _GEN_1399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1401 = 9'h179 == _GEN_9633 ? phv_data_377 : _GEN_1400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1402 = 9'h17a == _GEN_9633 ? phv_data_378 : _GEN_1401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1403 = 9'h17b == _GEN_9633 ? phv_data_379 : _GEN_1402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1404 = 9'h17c == _GEN_9633 ? phv_data_380 : _GEN_1403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1405 = 9'h17d == _GEN_9633 ? phv_data_381 : _GEN_1404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1406 = 9'h17e == _GEN_9633 ? phv_data_382 : _GEN_1405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1407 = 9'h17f == _GEN_9633 ? phv_data_383 : _GEN_1406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1408 = 9'h180 == _GEN_9633 ? phv_data_384 : _GEN_1407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1409 = 9'h181 == _GEN_9633 ? phv_data_385 : _GEN_1408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1410 = 9'h182 == _GEN_9633 ? phv_data_386 : _GEN_1409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1411 = 9'h183 == _GEN_9633 ? phv_data_387 : _GEN_1410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1412 = 9'h184 == _GEN_9633 ? phv_data_388 : _GEN_1411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1413 = 9'h185 == _GEN_9633 ? phv_data_389 : _GEN_1412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1414 = 9'h186 == _GEN_9633 ? phv_data_390 : _GEN_1413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1415 = 9'h187 == _GEN_9633 ? phv_data_391 : _GEN_1414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1416 = 9'h188 == _GEN_9633 ? phv_data_392 : _GEN_1415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1417 = 9'h189 == _GEN_9633 ? phv_data_393 : _GEN_1416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1418 = 9'h18a == _GEN_9633 ? phv_data_394 : _GEN_1417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1419 = 9'h18b == _GEN_9633 ? phv_data_395 : _GEN_1418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1420 = 9'h18c == _GEN_9633 ? phv_data_396 : _GEN_1419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1421 = 9'h18d == _GEN_9633 ? phv_data_397 : _GEN_1420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1422 = 9'h18e == _GEN_9633 ? phv_data_398 : _GEN_1421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1423 = 9'h18f == _GEN_9633 ? phv_data_399 : _GEN_1422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1424 = 9'h190 == _GEN_9633 ? phv_data_400 : _GEN_1423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1425 = 9'h191 == _GEN_9633 ? phv_data_401 : _GEN_1424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1426 = 9'h192 == _GEN_9633 ? phv_data_402 : _GEN_1425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1427 = 9'h193 == _GEN_9633 ? phv_data_403 : _GEN_1426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1428 = 9'h194 == _GEN_9633 ? phv_data_404 : _GEN_1427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1429 = 9'h195 == _GEN_9633 ? phv_data_405 : _GEN_1428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1430 = 9'h196 == _GEN_9633 ? phv_data_406 : _GEN_1429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1431 = 9'h197 == _GEN_9633 ? phv_data_407 : _GEN_1430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1432 = 9'h198 == _GEN_9633 ? phv_data_408 : _GEN_1431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1433 = 9'h199 == _GEN_9633 ? phv_data_409 : _GEN_1432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1434 = 9'h19a == _GEN_9633 ? phv_data_410 : _GEN_1433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1435 = 9'h19b == _GEN_9633 ? phv_data_411 : _GEN_1434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1436 = 9'h19c == _GEN_9633 ? phv_data_412 : _GEN_1435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1437 = 9'h19d == _GEN_9633 ? phv_data_413 : _GEN_1436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1438 = 9'h19e == _GEN_9633 ? phv_data_414 : _GEN_1437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1439 = 9'h19f == _GEN_9633 ? phv_data_415 : _GEN_1438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1440 = 9'h1a0 == _GEN_9633 ? phv_data_416 : _GEN_1439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1441 = 9'h1a1 == _GEN_9633 ? phv_data_417 : _GEN_1440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1442 = 9'h1a2 == _GEN_9633 ? phv_data_418 : _GEN_1441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1443 = 9'h1a3 == _GEN_9633 ? phv_data_419 : _GEN_1442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1444 = 9'h1a4 == _GEN_9633 ? phv_data_420 : _GEN_1443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1445 = 9'h1a5 == _GEN_9633 ? phv_data_421 : _GEN_1444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1446 = 9'h1a6 == _GEN_9633 ? phv_data_422 : _GEN_1445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1447 = 9'h1a7 == _GEN_9633 ? phv_data_423 : _GEN_1446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1448 = 9'h1a8 == _GEN_9633 ? phv_data_424 : _GEN_1447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1449 = 9'h1a9 == _GEN_9633 ? phv_data_425 : _GEN_1448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1450 = 9'h1aa == _GEN_9633 ? phv_data_426 : _GEN_1449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1451 = 9'h1ab == _GEN_9633 ? phv_data_427 : _GEN_1450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1452 = 9'h1ac == _GEN_9633 ? phv_data_428 : _GEN_1451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1453 = 9'h1ad == _GEN_9633 ? phv_data_429 : _GEN_1452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1454 = 9'h1ae == _GEN_9633 ? phv_data_430 : _GEN_1453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1455 = 9'h1af == _GEN_9633 ? phv_data_431 : _GEN_1454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1456 = 9'h1b0 == _GEN_9633 ? phv_data_432 : _GEN_1455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1457 = 9'h1b1 == _GEN_9633 ? phv_data_433 : _GEN_1456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1458 = 9'h1b2 == _GEN_9633 ? phv_data_434 : _GEN_1457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1459 = 9'h1b3 == _GEN_9633 ? phv_data_435 : _GEN_1458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1460 = 9'h1b4 == _GEN_9633 ? phv_data_436 : _GEN_1459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1461 = 9'h1b5 == _GEN_9633 ? phv_data_437 : _GEN_1460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1462 = 9'h1b6 == _GEN_9633 ? phv_data_438 : _GEN_1461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1463 = 9'h1b7 == _GEN_9633 ? phv_data_439 : _GEN_1462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1464 = 9'h1b8 == _GEN_9633 ? phv_data_440 : _GEN_1463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1465 = 9'h1b9 == _GEN_9633 ? phv_data_441 : _GEN_1464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1466 = 9'h1ba == _GEN_9633 ? phv_data_442 : _GEN_1465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1467 = 9'h1bb == _GEN_9633 ? phv_data_443 : _GEN_1466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1468 = 9'h1bc == _GEN_9633 ? phv_data_444 : _GEN_1467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1469 = 9'h1bd == _GEN_9633 ? phv_data_445 : _GEN_1468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1470 = 9'h1be == _GEN_9633 ? phv_data_446 : _GEN_1469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1471 = 9'h1bf == _GEN_9633 ? phv_data_447 : _GEN_1470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1472 = 9'h1c0 == _GEN_9633 ? phv_data_448 : _GEN_1471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1473 = 9'h1c1 == _GEN_9633 ? phv_data_449 : _GEN_1472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1474 = 9'h1c2 == _GEN_9633 ? phv_data_450 : _GEN_1473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1475 = 9'h1c3 == _GEN_9633 ? phv_data_451 : _GEN_1474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1476 = 9'h1c4 == _GEN_9633 ? phv_data_452 : _GEN_1475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1477 = 9'h1c5 == _GEN_9633 ? phv_data_453 : _GEN_1476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1478 = 9'h1c6 == _GEN_9633 ? phv_data_454 : _GEN_1477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1479 = 9'h1c7 == _GEN_9633 ? phv_data_455 : _GEN_1478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1480 = 9'h1c8 == _GEN_9633 ? phv_data_456 : _GEN_1479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1481 = 9'h1c9 == _GEN_9633 ? phv_data_457 : _GEN_1480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1482 = 9'h1ca == _GEN_9633 ? phv_data_458 : _GEN_1481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1483 = 9'h1cb == _GEN_9633 ? phv_data_459 : _GEN_1482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1484 = 9'h1cc == _GEN_9633 ? phv_data_460 : _GEN_1483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1485 = 9'h1cd == _GEN_9633 ? phv_data_461 : _GEN_1484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1486 = 9'h1ce == _GEN_9633 ? phv_data_462 : _GEN_1485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1487 = 9'h1cf == _GEN_9633 ? phv_data_463 : _GEN_1486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1488 = 9'h1d0 == _GEN_9633 ? phv_data_464 : _GEN_1487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1489 = 9'h1d1 == _GEN_9633 ? phv_data_465 : _GEN_1488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1490 = 9'h1d2 == _GEN_9633 ? phv_data_466 : _GEN_1489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1491 = 9'h1d3 == _GEN_9633 ? phv_data_467 : _GEN_1490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1492 = 9'h1d4 == _GEN_9633 ? phv_data_468 : _GEN_1491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1493 = 9'h1d5 == _GEN_9633 ? phv_data_469 : _GEN_1492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1494 = 9'h1d6 == _GEN_9633 ? phv_data_470 : _GEN_1493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1495 = 9'h1d7 == _GEN_9633 ? phv_data_471 : _GEN_1494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1496 = 9'h1d8 == _GEN_9633 ? phv_data_472 : _GEN_1495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1497 = 9'h1d9 == _GEN_9633 ? phv_data_473 : _GEN_1496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1498 = 9'h1da == _GEN_9633 ? phv_data_474 : _GEN_1497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1499 = 9'h1db == _GEN_9633 ? phv_data_475 : _GEN_1498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1500 = 9'h1dc == _GEN_9633 ? phv_data_476 : _GEN_1499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1501 = 9'h1dd == _GEN_9633 ? phv_data_477 : _GEN_1500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1502 = 9'h1de == _GEN_9633 ? phv_data_478 : _GEN_1501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1503 = 9'h1df == _GEN_9633 ? phv_data_479 : _GEN_1502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1504 = 9'h1e0 == _GEN_9633 ? phv_data_480 : _GEN_1503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1505 = 9'h1e1 == _GEN_9633 ? phv_data_481 : _GEN_1504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1506 = 9'h1e2 == _GEN_9633 ? phv_data_482 : _GEN_1505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1507 = 9'h1e3 == _GEN_9633 ? phv_data_483 : _GEN_1506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1508 = 9'h1e4 == _GEN_9633 ? phv_data_484 : _GEN_1507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1509 = 9'h1e5 == _GEN_9633 ? phv_data_485 : _GEN_1508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1510 = 9'h1e6 == _GEN_9633 ? phv_data_486 : _GEN_1509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1511 = 9'h1e7 == _GEN_9633 ? phv_data_487 : _GEN_1510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1512 = 9'h1e8 == _GEN_9633 ? phv_data_488 : _GEN_1511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1513 = 9'h1e9 == _GEN_9633 ? phv_data_489 : _GEN_1512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1514 = 9'h1ea == _GEN_9633 ? phv_data_490 : _GEN_1513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1515 = 9'h1eb == _GEN_9633 ? phv_data_491 : _GEN_1514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1516 = 9'h1ec == _GEN_9633 ? phv_data_492 : _GEN_1515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1517 = 9'h1ed == _GEN_9633 ? phv_data_493 : _GEN_1516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1518 = 9'h1ee == _GEN_9633 ? phv_data_494 : _GEN_1517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1519 = 9'h1ef == _GEN_9633 ? phv_data_495 : _GEN_1518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1520 = 9'h1f0 == _GEN_9633 ? phv_data_496 : _GEN_1519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1521 = 9'h1f1 == _GEN_9633 ? phv_data_497 : _GEN_1520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1522 = 9'h1f2 == _GEN_9633 ? phv_data_498 : _GEN_1521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1523 = 9'h1f3 == _GEN_9633 ? phv_data_499 : _GEN_1522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1524 = 9'h1f4 == _GEN_9633 ? phv_data_500 : _GEN_1523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1525 = 9'h1f5 == _GEN_9633 ? phv_data_501 : _GEN_1524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1526 = 9'h1f6 == _GEN_9633 ? phv_data_502 : _GEN_1525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1527 = 9'h1f7 == _GEN_9633 ? phv_data_503 : _GEN_1526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1528 = 9'h1f8 == _GEN_9633 ? phv_data_504 : _GEN_1527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1529 = 9'h1f9 == _GEN_9633 ? phv_data_505 : _GEN_1528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1530 = 9'h1fa == _GEN_9633 ? phv_data_506 : _GEN_1529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1531 = 9'h1fb == _GEN_9633 ? phv_data_507 : _GEN_1530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1532 = 9'h1fc == _GEN_9633 ? phv_data_508 : _GEN_1531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1533 = 9'h1fd == _GEN_9633 ? phv_data_509 : _GEN_1532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1534 = 9'h1fe == _GEN_9633 ? phv_data_510 : _GEN_1533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__1 = 9'h1ff == _GEN_9633 ? phv_data_511 : _GEN_1534; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask__1 = 2'h2 >= offset_0[1:0] & (2'h2 < ending | ending == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_3 = {total_offset_hi,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_1537 = 8'h1 == total_offset_3 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1538 = 8'h2 == total_offset_3 ? phv_data_2 : _GEN_1537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1539 = 8'h3 == total_offset_3 ? phv_data_3 : _GEN_1538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1540 = 8'h4 == total_offset_3 ? phv_data_4 : _GEN_1539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1541 = 8'h5 == total_offset_3 ? phv_data_5 : _GEN_1540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1542 = 8'h6 == total_offset_3 ? phv_data_6 : _GEN_1541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1543 = 8'h7 == total_offset_3 ? phv_data_7 : _GEN_1542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1544 = 8'h8 == total_offset_3 ? phv_data_8 : _GEN_1543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1545 = 8'h9 == total_offset_3 ? phv_data_9 : _GEN_1544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1546 = 8'ha == total_offset_3 ? phv_data_10 : _GEN_1545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1547 = 8'hb == total_offset_3 ? phv_data_11 : _GEN_1546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1548 = 8'hc == total_offset_3 ? phv_data_12 : _GEN_1547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1549 = 8'hd == total_offset_3 ? phv_data_13 : _GEN_1548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1550 = 8'he == total_offset_3 ? phv_data_14 : _GEN_1549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1551 = 8'hf == total_offset_3 ? phv_data_15 : _GEN_1550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1552 = 8'h10 == total_offset_3 ? phv_data_16 : _GEN_1551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1553 = 8'h11 == total_offset_3 ? phv_data_17 : _GEN_1552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1554 = 8'h12 == total_offset_3 ? phv_data_18 : _GEN_1553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1555 = 8'h13 == total_offset_3 ? phv_data_19 : _GEN_1554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1556 = 8'h14 == total_offset_3 ? phv_data_20 : _GEN_1555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1557 = 8'h15 == total_offset_3 ? phv_data_21 : _GEN_1556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1558 = 8'h16 == total_offset_3 ? phv_data_22 : _GEN_1557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1559 = 8'h17 == total_offset_3 ? phv_data_23 : _GEN_1558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1560 = 8'h18 == total_offset_3 ? phv_data_24 : _GEN_1559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1561 = 8'h19 == total_offset_3 ? phv_data_25 : _GEN_1560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1562 = 8'h1a == total_offset_3 ? phv_data_26 : _GEN_1561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1563 = 8'h1b == total_offset_3 ? phv_data_27 : _GEN_1562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1564 = 8'h1c == total_offset_3 ? phv_data_28 : _GEN_1563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1565 = 8'h1d == total_offset_3 ? phv_data_29 : _GEN_1564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1566 = 8'h1e == total_offset_3 ? phv_data_30 : _GEN_1565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1567 = 8'h1f == total_offset_3 ? phv_data_31 : _GEN_1566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1568 = 8'h20 == total_offset_3 ? phv_data_32 : _GEN_1567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1569 = 8'h21 == total_offset_3 ? phv_data_33 : _GEN_1568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1570 = 8'h22 == total_offset_3 ? phv_data_34 : _GEN_1569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1571 = 8'h23 == total_offset_3 ? phv_data_35 : _GEN_1570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1572 = 8'h24 == total_offset_3 ? phv_data_36 : _GEN_1571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1573 = 8'h25 == total_offset_3 ? phv_data_37 : _GEN_1572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1574 = 8'h26 == total_offset_3 ? phv_data_38 : _GEN_1573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1575 = 8'h27 == total_offset_3 ? phv_data_39 : _GEN_1574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1576 = 8'h28 == total_offset_3 ? phv_data_40 : _GEN_1575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1577 = 8'h29 == total_offset_3 ? phv_data_41 : _GEN_1576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1578 = 8'h2a == total_offset_3 ? phv_data_42 : _GEN_1577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1579 = 8'h2b == total_offset_3 ? phv_data_43 : _GEN_1578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1580 = 8'h2c == total_offset_3 ? phv_data_44 : _GEN_1579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1581 = 8'h2d == total_offset_3 ? phv_data_45 : _GEN_1580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1582 = 8'h2e == total_offset_3 ? phv_data_46 : _GEN_1581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1583 = 8'h2f == total_offset_3 ? phv_data_47 : _GEN_1582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1584 = 8'h30 == total_offset_3 ? phv_data_48 : _GEN_1583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1585 = 8'h31 == total_offset_3 ? phv_data_49 : _GEN_1584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1586 = 8'h32 == total_offset_3 ? phv_data_50 : _GEN_1585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1587 = 8'h33 == total_offset_3 ? phv_data_51 : _GEN_1586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1588 = 8'h34 == total_offset_3 ? phv_data_52 : _GEN_1587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1589 = 8'h35 == total_offset_3 ? phv_data_53 : _GEN_1588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1590 = 8'h36 == total_offset_3 ? phv_data_54 : _GEN_1589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1591 = 8'h37 == total_offset_3 ? phv_data_55 : _GEN_1590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1592 = 8'h38 == total_offset_3 ? phv_data_56 : _GEN_1591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1593 = 8'h39 == total_offset_3 ? phv_data_57 : _GEN_1592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1594 = 8'h3a == total_offset_3 ? phv_data_58 : _GEN_1593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1595 = 8'h3b == total_offset_3 ? phv_data_59 : _GEN_1594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1596 = 8'h3c == total_offset_3 ? phv_data_60 : _GEN_1595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1597 = 8'h3d == total_offset_3 ? phv_data_61 : _GEN_1596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1598 = 8'h3e == total_offset_3 ? phv_data_62 : _GEN_1597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1599 = 8'h3f == total_offset_3 ? phv_data_63 : _GEN_1598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1600 = 8'h40 == total_offset_3 ? phv_data_64 : _GEN_1599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1601 = 8'h41 == total_offset_3 ? phv_data_65 : _GEN_1600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1602 = 8'h42 == total_offset_3 ? phv_data_66 : _GEN_1601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1603 = 8'h43 == total_offset_3 ? phv_data_67 : _GEN_1602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1604 = 8'h44 == total_offset_3 ? phv_data_68 : _GEN_1603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1605 = 8'h45 == total_offset_3 ? phv_data_69 : _GEN_1604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1606 = 8'h46 == total_offset_3 ? phv_data_70 : _GEN_1605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1607 = 8'h47 == total_offset_3 ? phv_data_71 : _GEN_1606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1608 = 8'h48 == total_offset_3 ? phv_data_72 : _GEN_1607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1609 = 8'h49 == total_offset_3 ? phv_data_73 : _GEN_1608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1610 = 8'h4a == total_offset_3 ? phv_data_74 : _GEN_1609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1611 = 8'h4b == total_offset_3 ? phv_data_75 : _GEN_1610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1612 = 8'h4c == total_offset_3 ? phv_data_76 : _GEN_1611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1613 = 8'h4d == total_offset_3 ? phv_data_77 : _GEN_1612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1614 = 8'h4e == total_offset_3 ? phv_data_78 : _GEN_1613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1615 = 8'h4f == total_offset_3 ? phv_data_79 : _GEN_1614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1616 = 8'h50 == total_offset_3 ? phv_data_80 : _GEN_1615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1617 = 8'h51 == total_offset_3 ? phv_data_81 : _GEN_1616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1618 = 8'h52 == total_offset_3 ? phv_data_82 : _GEN_1617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1619 = 8'h53 == total_offset_3 ? phv_data_83 : _GEN_1618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1620 = 8'h54 == total_offset_3 ? phv_data_84 : _GEN_1619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1621 = 8'h55 == total_offset_3 ? phv_data_85 : _GEN_1620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1622 = 8'h56 == total_offset_3 ? phv_data_86 : _GEN_1621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1623 = 8'h57 == total_offset_3 ? phv_data_87 : _GEN_1622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1624 = 8'h58 == total_offset_3 ? phv_data_88 : _GEN_1623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1625 = 8'h59 == total_offset_3 ? phv_data_89 : _GEN_1624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1626 = 8'h5a == total_offset_3 ? phv_data_90 : _GEN_1625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1627 = 8'h5b == total_offset_3 ? phv_data_91 : _GEN_1626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1628 = 8'h5c == total_offset_3 ? phv_data_92 : _GEN_1627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1629 = 8'h5d == total_offset_3 ? phv_data_93 : _GEN_1628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1630 = 8'h5e == total_offset_3 ? phv_data_94 : _GEN_1629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1631 = 8'h5f == total_offset_3 ? phv_data_95 : _GEN_1630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1632 = 8'h60 == total_offset_3 ? phv_data_96 : _GEN_1631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1633 = 8'h61 == total_offset_3 ? phv_data_97 : _GEN_1632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1634 = 8'h62 == total_offset_3 ? phv_data_98 : _GEN_1633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1635 = 8'h63 == total_offset_3 ? phv_data_99 : _GEN_1634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1636 = 8'h64 == total_offset_3 ? phv_data_100 : _GEN_1635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1637 = 8'h65 == total_offset_3 ? phv_data_101 : _GEN_1636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1638 = 8'h66 == total_offset_3 ? phv_data_102 : _GEN_1637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1639 = 8'h67 == total_offset_3 ? phv_data_103 : _GEN_1638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1640 = 8'h68 == total_offset_3 ? phv_data_104 : _GEN_1639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1641 = 8'h69 == total_offset_3 ? phv_data_105 : _GEN_1640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1642 = 8'h6a == total_offset_3 ? phv_data_106 : _GEN_1641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1643 = 8'h6b == total_offset_3 ? phv_data_107 : _GEN_1642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1644 = 8'h6c == total_offset_3 ? phv_data_108 : _GEN_1643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1645 = 8'h6d == total_offset_3 ? phv_data_109 : _GEN_1644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1646 = 8'h6e == total_offset_3 ? phv_data_110 : _GEN_1645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1647 = 8'h6f == total_offset_3 ? phv_data_111 : _GEN_1646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1648 = 8'h70 == total_offset_3 ? phv_data_112 : _GEN_1647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1649 = 8'h71 == total_offset_3 ? phv_data_113 : _GEN_1648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1650 = 8'h72 == total_offset_3 ? phv_data_114 : _GEN_1649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1651 = 8'h73 == total_offset_3 ? phv_data_115 : _GEN_1650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1652 = 8'h74 == total_offset_3 ? phv_data_116 : _GEN_1651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1653 = 8'h75 == total_offset_3 ? phv_data_117 : _GEN_1652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1654 = 8'h76 == total_offset_3 ? phv_data_118 : _GEN_1653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1655 = 8'h77 == total_offset_3 ? phv_data_119 : _GEN_1654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1656 = 8'h78 == total_offset_3 ? phv_data_120 : _GEN_1655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1657 = 8'h79 == total_offset_3 ? phv_data_121 : _GEN_1656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1658 = 8'h7a == total_offset_3 ? phv_data_122 : _GEN_1657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1659 = 8'h7b == total_offset_3 ? phv_data_123 : _GEN_1658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1660 = 8'h7c == total_offset_3 ? phv_data_124 : _GEN_1659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1661 = 8'h7d == total_offset_3 ? phv_data_125 : _GEN_1660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1662 = 8'h7e == total_offset_3 ? phv_data_126 : _GEN_1661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1663 = 8'h7f == total_offset_3 ? phv_data_127 : _GEN_1662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1664 = 8'h80 == total_offset_3 ? phv_data_128 : _GEN_1663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1665 = 8'h81 == total_offset_3 ? phv_data_129 : _GEN_1664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1666 = 8'h82 == total_offset_3 ? phv_data_130 : _GEN_1665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1667 = 8'h83 == total_offset_3 ? phv_data_131 : _GEN_1666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1668 = 8'h84 == total_offset_3 ? phv_data_132 : _GEN_1667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1669 = 8'h85 == total_offset_3 ? phv_data_133 : _GEN_1668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1670 = 8'h86 == total_offset_3 ? phv_data_134 : _GEN_1669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1671 = 8'h87 == total_offset_3 ? phv_data_135 : _GEN_1670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1672 = 8'h88 == total_offset_3 ? phv_data_136 : _GEN_1671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1673 = 8'h89 == total_offset_3 ? phv_data_137 : _GEN_1672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1674 = 8'h8a == total_offset_3 ? phv_data_138 : _GEN_1673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1675 = 8'h8b == total_offset_3 ? phv_data_139 : _GEN_1674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1676 = 8'h8c == total_offset_3 ? phv_data_140 : _GEN_1675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1677 = 8'h8d == total_offset_3 ? phv_data_141 : _GEN_1676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1678 = 8'h8e == total_offset_3 ? phv_data_142 : _GEN_1677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1679 = 8'h8f == total_offset_3 ? phv_data_143 : _GEN_1678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1680 = 8'h90 == total_offset_3 ? phv_data_144 : _GEN_1679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1681 = 8'h91 == total_offset_3 ? phv_data_145 : _GEN_1680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1682 = 8'h92 == total_offset_3 ? phv_data_146 : _GEN_1681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1683 = 8'h93 == total_offset_3 ? phv_data_147 : _GEN_1682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1684 = 8'h94 == total_offset_3 ? phv_data_148 : _GEN_1683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1685 = 8'h95 == total_offset_3 ? phv_data_149 : _GEN_1684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1686 = 8'h96 == total_offset_3 ? phv_data_150 : _GEN_1685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1687 = 8'h97 == total_offset_3 ? phv_data_151 : _GEN_1686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1688 = 8'h98 == total_offset_3 ? phv_data_152 : _GEN_1687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1689 = 8'h99 == total_offset_3 ? phv_data_153 : _GEN_1688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1690 = 8'h9a == total_offset_3 ? phv_data_154 : _GEN_1689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1691 = 8'h9b == total_offset_3 ? phv_data_155 : _GEN_1690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1692 = 8'h9c == total_offset_3 ? phv_data_156 : _GEN_1691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1693 = 8'h9d == total_offset_3 ? phv_data_157 : _GEN_1692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1694 = 8'h9e == total_offset_3 ? phv_data_158 : _GEN_1693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1695 = 8'h9f == total_offset_3 ? phv_data_159 : _GEN_1694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1696 = 8'ha0 == total_offset_3 ? phv_data_160 : _GEN_1695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1697 = 8'ha1 == total_offset_3 ? phv_data_161 : _GEN_1696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1698 = 8'ha2 == total_offset_3 ? phv_data_162 : _GEN_1697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1699 = 8'ha3 == total_offset_3 ? phv_data_163 : _GEN_1698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1700 = 8'ha4 == total_offset_3 ? phv_data_164 : _GEN_1699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1701 = 8'ha5 == total_offset_3 ? phv_data_165 : _GEN_1700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1702 = 8'ha6 == total_offset_3 ? phv_data_166 : _GEN_1701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1703 = 8'ha7 == total_offset_3 ? phv_data_167 : _GEN_1702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1704 = 8'ha8 == total_offset_3 ? phv_data_168 : _GEN_1703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1705 = 8'ha9 == total_offset_3 ? phv_data_169 : _GEN_1704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1706 = 8'haa == total_offset_3 ? phv_data_170 : _GEN_1705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1707 = 8'hab == total_offset_3 ? phv_data_171 : _GEN_1706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1708 = 8'hac == total_offset_3 ? phv_data_172 : _GEN_1707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1709 = 8'had == total_offset_3 ? phv_data_173 : _GEN_1708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1710 = 8'hae == total_offset_3 ? phv_data_174 : _GEN_1709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1711 = 8'haf == total_offset_3 ? phv_data_175 : _GEN_1710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1712 = 8'hb0 == total_offset_3 ? phv_data_176 : _GEN_1711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1713 = 8'hb1 == total_offset_3 ? phv_data_177 : _GEN_1712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1714 = 8'hb2 == total_offset_3 ? phv_data_178 : _GEN_1713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1715 = 8'hb3 == total_offset_3 ? phv_data_179 : _GEN_1714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1716 = 8'hb4 == total_offset_3 ? phv_data_180 : _GEN_1715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1717 = 8'hb5 == total_offset_3 ? phv_data_181 : _GEN_1716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1718 = 8'hb6 == total_offset_3 ? phv_data_182 : _GEN_1717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1719 = 8'hb7 == total_offset_3 ? phv_data_183 : _GEN_1718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1720 = 8'hb8 == total_offset_3 ? phv_data_184 : _GEN_1719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1721 = 8'hb9 == total_offset_3 ? phv_data_185 : _GEN_1720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1722 = 8'hba == total_offset_3 ? phv_data_186 : _GEN_1721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1723 = 8'hbb == total_offset_3 ? phv_data_187 : _GEN_1722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1724 = 8'hbc == total_offset_3 ? phv_data_188 : _GEN_1723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1725 = 8'hbd == total_offset_3 ? phv_data_189 : _GEN_1724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1726 = 8'hbe == total_offset_3 ? phv_data_190 : _GEN_1725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1727 = 8'hbf == total_offset_3 ? phv_data_191 : _GEN_1726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1728 = 8'hc0 == total_offset_3 ? phv_data_192 : _GEN_1727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1729 = 8'hc1 == total_offset_3 ? phv_data_193 : _GEN_1728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1730 = 8'hc2 == total_offset_3 ? phv_data_194 : _GEN_1729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1731 = 8'hc3 == total_offset_3 ? phv_data_195 : _GEN_1730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1732 = 8'hc4 == total_offset_3 ? phv_data_196 : _GEN_1731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1733 = 8'hc5 == total_offset_3 ? phv_data_197 : _GEN_1732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1734 = 8'hc6 == total_offset_3 ? phv_data_198 : _GEN_1733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1735 = 8'hc7 == total_offset_3 ? phv_data_199 : _GEN_1734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1736 = 8'hc8 == total_offset_3 ? phv_data_200 : _GEN_1735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1737 = 8'hc9 == total_offset_3 ? phv_data_201 : _GEN_1736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1738 = 8'hca == total_offset_3 ? phv_data_202 : _GEN_1737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1739 = 8'hcb == total_offset_3 ? phv_data_203 : _GEN_1738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1740 = 8'hcc == total_offset_3 ? phv_data_204 : _GEN_1739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1741 = 8'hcd == total_offset_3 ? phv_data_205 : _GEN_1740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1742 = 8'hce == total_offset_3 ? phv_data_206 : _GEN_1741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1743 = 8'hcf == total_offset_3 ? phv_data_207 : _GEN_1742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1744 = 8'hd0 == total_offset_3 ? phv_data_208 : _GEN_1743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1745 = 8'hd1 == total_offset_3 ? phv_data_209 : _GEN_1744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1746 = 8'hd2 == total_offset_3 ? phv_data_210 : _GEN_1745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1747 = 8'hd3 == total_offset_3 ? phv_data_211 : _GEN_1746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1748 = 8'hd4 == total_offset_3 ? phv_data_212 : _GEN_1747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1749 = 8'hd5 == total_offset_3 ? phv_data_213 : _GEN_1748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1750 = 8'hd6 == total_offset_3 ? phv_data_214 : _GEN_1749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1751 = 8'hd7 == total_offset_3 ? phv_data_215 : _GEN_1750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1752 = 8'hd8 == total_offset_3 ? phv_data_216 : _GEN_1751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1753 = 8'hd9 == total_offset_3 ? phv_data_217 : _GEN_1752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1754 = 8'hda == total_offset_3 ? phv_data_218 : _GEN_1753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1755 = 8'hdb == total_offset_3 ? phv_data_219 : _GEN_1754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1756 = 8'hdc == total_offset_3 ? phv_data_220 : _GEN_1755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1757 = 8'hdd == total_offset_3 ? phv_data_221 : _GEN_1756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1758 = 8'hde == total_offset_3 ? phv_data_222 : _GEN_1757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1759 = 8'hdf == total_offset_3 ? phv_data_223 : _GEN_1758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1760 = 8'he0 == total_offset_3 ? phv_data_224 : _GEN_1759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1761 = 8'he1 == total_offset_3 ? phv_data_225 : _GEN_1760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1762 = 8'he2 == total_offset_3 ? phv_data_226 : _GEN_1761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1763 = 8'he3 == total_offset_3 ? phv_data_227 : _GEN_1762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1764 = 8'he4 == total_offset_3 ? phv_data_228 : _GEN_1763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1765 = 8'he5 == total_offset_3 ? phv_data_229 : _GEN_1764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1766 = 8'he6 == total_offset_3 ? phv_data_230 : _GEN_1765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1767 = 8'he7 == total_offset_3 ? phv_data_231 : _GEN_1766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1768 = 8'he8 == total_offset_3 ? phv_data_232 : _GEN_1767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1769 = 8'he9 == total_offset_3 ? phv_data_233 : _GEN_1768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1770 = 8'hea == total_offset_3 ? phv_data_234 : _GEN_1769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1771 = 8'heb == total_offset_3 ? phv_data_235 : _GEN_1770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1772 = 8'hec == total_offset_3 ? phv_data_236 : _GEN_1771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1773 = 8'hed == total_offset_3 ? phv_data_237 : _GEN_1772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1774 = 8'hee == total_offset_3 ? phv_data_238 : _GEN_1773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1775 = 8'hef == total_offset_3 ? phv_data_239 : _GEN_1774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1776 = 8'hf0 == total_offset_3 ? phv_data_240 : _GEN_1775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1777 = 8'hf1 == total_offset_3 ? phv_data_241 : _GEN_1776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1778 = 8'hf2 == total_offset_3 ? phv_data_242 : _GEN_1777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1779 = 8'hf3 == total_offset_3 ? phv_data_243 : _GEN_1778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1780 = 8'hf4 == total_offset_3 ? phv_data_244 : _GEN_1779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1781 = 8'hf5 == total_offset_3 ? phv_data_245 : _GEN_1780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1782 = 8'hf6 == total_offset_3 ? phv_data_246 : _GEN_1781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1783 = 8'hf7 == total_offset_3 ? phv_data_247 : _GEN_1782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1784 = 8'hf8 == total_offset_3 ? phv_data_248 : _GEN_1783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1785 = 8'hf9 == total_offset_3 ? phv_data_249 : _GEN_1784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1786 = 8'hfa == total_offset_3 ? phv_data_250 : _GEN_1785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1787 = 8'hfb == total_offset_3 ? phv_data_251 : _GEN_1786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1788 = 8'hfc == total_offset_3 ? phv_data_252 : _GEN_1787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1789 = 8'hfd == total_offset_3 ? phv_data_253 : _GEN_1788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1790 = 8'hfe == total_offset_3 ? phv_data_254 : _GEN_1789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1791 = 8'hff == total_offset_3 ? phv_data_255 : _GEN_1790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_9889 = {{1'd0}, total_offset_3}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1792 = 9'h100 == _GEN_9889 ? phv_data_256 : _GEN_1791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1793 = 9'h101 == _GEN_9889 ? phv_data_257 : _GEN_1792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1794 = 9'h102 == _GEN_9889 ? phv_data_258 : _GEN_1793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1795 = 9'h103 == _GEN_9889 ? phv_data_259 : _GEN_1794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1796 = 9'h104 == _GEN_9889 ? phv_data_260 : _GEN_1795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1797 = 9'h105 == _GEN_9889 ? phv_data_261 : _GEN_1796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1798 = 9'h106 == _GEN_9889 ? phv_data_262 : _GEN_1797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1799 = 9'h107 == _GEN_9889 ? phv_data_263 : _GEN_1798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1800 = 9'h108 == _GEN_9889 ? phv_data_264 : _GEN_1799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1801 = 9'h109 == _GEN_9889 ? phv_data_265 : _GEN_1800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1802 = 9'h10a == _GEN_9889 ? phv_data_266 : _GEN_1801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1803 = 9'h10b == _GEN_9889 ? phv_data_267 : _GEN_1802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1804 = 9'h10c == _GEN_9889 ? phv_data_268 : _GEN_1803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1805 = 9'h10d == _GEN_9889 ? phv_data_269 : _GEN_1804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1806 = 9'h10e == _GEN_9889 ? phv_data_270 : _GEN_1805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1807 = 9'h10f == _GEN_9889 ? phv_data_271 : _GEN_1806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1808 = 9'h110 == _GEN_9889 ? phv_data_272 : _GEN_1807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1809 = 9'h111 == _GEN_9889 ? phv_data_273 : _GEN_1808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1810 = 9'h112 == _GEN_9889 ? phv_data_274 : _GEN_1809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1811 = 9'h113 == _GEN_9889 ? phv_data_275 : _GEN_1810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1812 = 9'h114 == _GEN_9889 ? phv_data_276 : _GEN_1811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1813 = 9'h115 == _GEN_9889 ? phv_data_277 : _GEN_1812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1814 = 9'h116 == _GEN_9889 ? phv_data_278 : _GEN_1813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1815 = 9'h117 == _GEN_9889 ? phv_data_279 : _GEN_1814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1816 = 9'h118 == _GEN_9889 ? phv_data_280 : _GEN_1815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1817 = 9'h119 == _GEN_9889 ? phv_data_281 : _GEN_1816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1818 = 9'h11a == _GEN_9889 ? phv_data_282 : _GEN_1817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1819 = 9'h11b == _GEN_9889 ? phv_data_283 : _GEN_1818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1820 = 9'h11c == _GEN_9889 ? phv_data_284 : _GEN_1819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1821 = 9'h11d == _GEN_9889 ? phv_data_285 : _GEN_1820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1822 = 9'h11e == _GEN_9889 ? phv_data_286 : _GEN_1821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1823 = 9'h11f == _GEN_9889 ? phv_data_287 : _GEN_1822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1824 = 9'h120 == _GEN_9889 ? phv_data_288 : _GEN_1823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1825 = 9'h121 == _GEN_9889 ? phv_data_289 : _GEN_1824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1826 = 9'h122 == _GEN_9889 ? phv_data_290 : _GEN_1825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1827 = 9'h123 == _GEN_9889 ? phv_data_291 : _GEN_1826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1828 = 9'h124 == _GEN_9889 ? phv_data_292 : _GEN_1827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1829 = 9'h125 == _GEN_9889 ? phv_data_293 : _GEN_1828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1830 = 9'h126 == _GEN_9889 ? phv_data_294 : _GEN_1829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1831 = 9'h127 == _GEN_9889 ? phv_data_295 : _GEN_1830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1832 = 9'h128 == _GEN_9889 ? phv_data_296 : _GEN_1831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1833 = 9'h129 == _GEN_9889 ? phv_data_297 : _GEN_1832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1834 = 9'h12a == _GEN_9889 ? phv_data_298 : _GEN_1833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1835 = 9'h12b == _GEN_9889 ? phv_data_299 : _GEN_1834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1836 = 9'h12c == _GEN_9889 ? phv_data_300 : _GEN_1835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1837 = 9'h12d == _GEN_9889 ? phv_data_301 : _GEN_1836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1838 = 9'h12e == _GEN_9889 ? phv_data_302 : _GEN_1837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1839 = 9'h12f == _GEN_9889 ? phv_data_303 : _GEN_1838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1840 = 9'h130 == _GEN_9889 ? phv_data_304 : _GEN_1839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1841 = 9'h131 == _GEN_9889 ? phv_data_305 : _GEN_1840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1842 = 9'h132 == _GEN_9889 ? phv_data_306 : _GEN_1841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1843 = 9'h133 == _GEN_9889 ? phv_data_307 : _GEN_1842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1844 = 9'h134 == _GEN_9889 ? phv_data_308 : _GEN_1843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1845 = 9'h135 == _GEN_9889 ? phv_data_309 : _GEN_1844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1846 = 9'h136 == _GEN_9889 ? phv_data_310 : _GEN_1845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1847 = 9'h137 == _GEN_9889 ? phv_data_311 : _GEN_1846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1848 = 9'h138 == _GEN_9889 ? phv_data_312 : _GEN_1847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1849 = 9'h139 == _GEN_9889 ? phv_data_313 : _GEN_1848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1850 = 9'h13a == _GEN_9889 ? phv_data_314 : _GEN_1849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1851 = 9'h13b == _GEN_9889 ? phv_data_315 : _GEN_1850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1852 = 9'h13c == _GEN_9889 ? phv_data_316 : _GEN_1851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1853 = 9'h13d == _GEN_9889 ? phv_data_317 : _GEN_1852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1854 = 9'h13e == _GEN_9889 ? phv_data_318 : _GEN_1853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1855 = 9'h13f == _GEN_9889 ? phv_data_319 : _GEN_1854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1856 = 9'h140 == _GEN_9889 ? phv_data_320 : _GEN_1855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1857 = 9'h141 == _GEN_9889 ? phv_data_321 : _GEN_1856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1858 = 9'h142 == _GEN_9889 ? phv_data_322 : _GEN_1857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1859 = 9'h143 == _GEN_9889 ? phv_data_323 : _GEN_1858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1860 = 9'h144 == _GEN_9889 ? phv_data_324 : _GEN_1859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1861 = 9'h145 == _GEN_9889 ? phv_data_325 : _GEN_1860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1862 = 9'h146 == _GEN_9889 ? phv_data_326 : _GEN_1861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1863 = 9'h147 == _GEN_9889 ? phv_data_327 : _GEN_1862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1864 = 9'h148 == _GEN_9889 ? phv_data_328 : _GEN_1863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1865 = 9'h149 == _GEN_9889 ? phv_data_329 : _GEN_1864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1866 = 9'h14a == _GEN_9889 ? phv_data_330 : _GEN_1865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1867 = 9'h14b == _GEN_9889 ? phv_data_331 : _GEN_1866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1868 = 9'h14c == _GEN_9889 ? phv_data_332 : _GEN_1867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1869 = 9'h14d == _GEN_9889 ? phv_data_333 : _GEN_1868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1870 = 9'h14e == _GEN_9889 ? phv_data_334 : _GEN_1869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1871 = 9'h14f == _GEN_9889 ? phv_data_335 : _GEN_1870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1872 = 9'h150 == _GEN_9889 ? phv_data_336 : _GEN_1871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1873 = 9'h151 == _GEN_9889 ? phv_data_337 : _GEN_1872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1874 = 9'h152 == _GEN_9889 ? phv_data_338 : _GEN_1873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1875 = 9'h153 == _GEN_9889 ? phv_data_339 : _GEN_1874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1876 = 9'h154 == _GEN_9889 ? phv_data_340 : _GEN_1875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1877 = 9'h155 == _GEN_9889 ? phv_data_341 : _GEN_1876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1878 = 9'h156 == _GEN_9889 ? phv_data_342 : _GEN_1877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1879 = 9'h157 == _GEN_9889 ? phv_data_343 : _GEN_1878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1880 = 9'h158 == _GEN_9889 ? phv_data_344 : _GEN_1879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1881 = 9'h159 == _GEN_9889 ? phv_data_345 : _GEN_1880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1882 = 9'h15a == _GEN_9889 ? phv_data_346 : _GEN_1881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1883 = 9'h15b == _GEN_9889 ? phv_data_347 : _GEN_1882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1884 = 9'h15c == _GEN_9889 ? phv_data_348 : _GEN_1883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1885 = 9'h15d == _GEN_9889 ? phv_data_349 : _GEN_1884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1886 = 9'h15e == _GEN_9889 ? phv_data_350 : _GEN_1885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1887 = 9'h15f == _GEN_9889 ? phv_data_351 : _GEN_1886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1888 = 9'h160 == _GEN_9889 ? phv_data_352 : _GEN_1887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1889 = 9'h161 == _GEN_9889 ? phv_data_353 : _GEN_1888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1890 = 9'h162 == _GEN_9889 ? phv_data_354 : _GEN_1889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1891 = 9'h163 == _GEN_9889 ? phv_data_355 : _GEN_1890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1892 = 9'h164 == _GEN_9889 ? phv_data_356 : _GEN_1891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1893 = 9'h165 == _GEN_9889 ? phv_data_357 : _GEN_1892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1894 = 9'h166 == _GEN_9889 ? phv_data_358 : _GEN_1893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1895 = 9'h167 == _GEN_9889 ? phv_data_359 : _GEN_1894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1896 = 9'h168 == _GEN_9889 ? phv_data_360 : _GEN_1895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1897 = 9'h169 == _GEN_9889 ? phv_data_361 : _GEN_1896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1898 = 9'h16a == _GEN_9889 ? phv_data_362 : _GEN_1897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1899 = 9'h16b == _GEN_9889 ? phv_data_363 : _GEN_1898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1900 = 9'h16c == _GEN_9889 ? phv_data_364 : _GEN_1899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1901 = 9'h16d == _GEN_9889 ? phv_data_365 : _GEN_1900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1902 = 9'h16e == _GEN_9889 ? phv_data_366 : _GEN_1901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1903 = 9'h16f == _GEN_9889 ? phv_data_367 : _GEN_1902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1904 = 9'h170 == _GEN_9889 ? phv_data_368 : _GEN_1903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1905 = 9'h171 == _GEN_9889 ? phv_data_369 : _GEN_1904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1906 = 9'h172 == _GEN_9889 ? phv_data_370 : _GEN_1905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1907 = 9'h173 == _GEN_9889 ? phv_data_371 : _GEN_1906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1908 = 9'h174 == _GEN_9889 ? phv_data_372 : _GEN_1907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1909 = 9'h175 == _GEN_9889 ? phv_data_373 : _GEN_1908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1910 = 9'h176 == _GEN_9889 ? phv_data_374 : _GEN_1909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1911 = 9'h177 == _GEN_9889 ? phv_data_375 : _GEN_1910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1912 = 9'h178 == _GEN_9889 ? phv_data_376 : _GEN_1911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1913 = 9'h179 == _GEN_9889 ? phv_data_377 : _GEN_1912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1914 = 9'h17a == _GEN_9889 ? phv_data_378 : _GEN_1913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1915 = 9'h17b == _GEN_9889 ? phv_data_379 : _GEN_1914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1916 = 9'h17c == _GEN_9889 ? phv_data_380 : _GEN_1915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1917 = 9'h17d == _GEN_9889 ? phv_data_381 : _GEN_1916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1918 = 9'h17e == _GEN_9889 ? phv_data_382 : _GEN_1917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1919 = 9'h17f == _GEN_9889 ? phv_data_383 : _GEN_1918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1920 = 9'h180 == _GEN_9889 ? phv_data_384 : _GEN_1919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1921 = 9'h181 == _GEN_9889 ? phv_data_385 : _GEN_1920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1922 = 9'h182 == _GEN_9889 ? phv_data_386 : _GEN_1921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1923 = 9'h183 == _GEN_9889 ? phv_data_387 : _GEN_1922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1924 = 9'h184 == _GEN_9889 ? phv_data_388 : _GEN_1923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1925 = 9'h185 == _GEN_9889 ? phv_data_389 : _GEN_1924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1926 = 9'h186 == _GEN_9889 ? phv_data_390 : _GEN_1925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1927 = 9'h187 == _GEN_9889 ? phv_data_391 : _GEN_1926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1928 = 9'h188 == _GEN_9889 ? phv_data_392 : _GEN_1927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1929 = 9'h189 == _GEN_9889 ? phv_data_393 : _GEN_1928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1930 = 9'h18a == _GEN_9889 ? phv_data_394 : _GEN_1929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1931 = 9'h18b == _GEN_9889 ? phv_data_395 : _GEN_1930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1932 = 9'h18c == _GEN_9889 ? phv_data_396 : _GEN_1931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1933 = 9'h18d == _GEN_9889 ? phv_data_397 : _GEN_1932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1934 = 9'h18e == _GEN_9889 ? phv_data_398 : _GEN_1933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1935 = 9'h18f == _GEN_9889 ? phv_data_399 : _GEN_1934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1936 = 9'h190 == _GEN_9889 ? phv_data_400 : _GEN_1935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1937 = 9'h191 == _GEN_9889 ? phv_data_401 : _GEN_1936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1938 = 9'h192 == _GEN_9889 ? phv_data_402 : _GEN_1937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1939 = 9'h193 == _GEN_9889 ? phv_data_403 : _GEN_1938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1940 = 9'h194 == _GEN_9889 ? phv_data_404 : _GEN_1939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1941 = 9'h195 == _GEN_9889 ? phv_data_405 : _GEN_1940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1942 = 9'h196 == _GEN_9889 ? phv_data_406 : _GEN_1941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1943 = 9'h197 == _GEN_9889 ? phv_data_407 : _GEN_1942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1944 = 9'h198 == _GEN_9889 ? phv_data_408 : _GEN_1943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1945 = 9'h199 == _GEN_9889 ? phv_data_409 : _GEN_1944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1946 = 9'h19a == _GEN_9889 ? phv_data_410 : _GEN_1945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1947 = 9'h19b == _GEN_9889 ? phv_data_411 : _GEN_1946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1948 = 9'h19c == _GEN_9889 ? phv_data_412 : _GEN_1947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1949 = 9'h19d == _GEN_9889 ? phv_data_413 : _GEN_1948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1950 = 9'h19e == _GEN_9889 ? phv_data_414 : _GEN_1949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1951 = 9'h19f == _GEN_9889 ? phv_data_415 : _GEN_1950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1952 = 9'h1a0 == _GEN_9889 ? phv_data_416 : _GEN_1951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1953 = 9'h1a1 == _GEN_9889 ? phv_data_417 : _GEN_1952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1954 = 9'h1a2 == _GEN_9889 ? phv_data_418 : _GEN_1953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1955 = 9'h1a3 == _GEN_9889 ? phv_data_419 : _GEN_1954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1956 = 9'h1a4 == _GEN_9889 ? phv_data_420 : _GEN_1955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1957 = 9'h1a5 == _GEN_9889 ? phv_data_421 : _GEN_1956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1958 = 9'h1a6 == _GEN_9889 ? phv_data_422 : _GEN_1957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1959 = 9'h1a7 == _GEN_9889 ? phv_data_423 : _GEN_1958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1960 = 9'h1a8 == _GEN_9889 ? phv_data_424 : _GEN_1959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1961 = 9'h1a9 == _GEN_9889 ? phv_data_425 : _GEN_1960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1962 = 9'h1aa == _GEN_9889 ? phv_data_426 : _GEN_1961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1963 = 9'h1ab == _GEN_9889 ? phv_data_427 : _GEN_1962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1964 = 9'h1ac == _GEN_9889 ? phv_data_428 : _GEN_1963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1965 = 9'h1ad == _GEN_9889 ? phv_data_429 : _GEN_1964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1966 = 9'h1ae == _GEN_9889 ? phv_data_430 : _GEN_1965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1967 = 9'h1af == _GEN_9889 ? phv_data_431 : _GEN_1966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1968 = 9'h1b0 == _GEN_9889 ? phv_data_432 : _GEN_1967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1969 = 9'h1b1 == _GEN_9889 ? phv_data_433 : _GEN_1968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1970 = 9'h1b2 == _GEN_9889 ? phv_data_434 : _GEN_1969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1971 = 9'h1b3 == _GEN_9889 ? phv_data_435 : _GEN_1970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1972 = 9'h1b4 == _GEN_9889 ? phv_data_436 : _GEN_1971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1973 = 9'h1b5 == _GEN_9889 ? phv_data_437 : _GEN_1972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1974 = 9'h1b6 == _GEN_9889 ? phv_data_438 : _GEN_1973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1975 = 9'h1b7 == _GEN_9889 ? phv_data_439 : _GEN_1974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1976 = 9'h1b8 == _GEN_9889 ? phv_data_440 : _GEN_1975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1977 = 9'h1b9 == _GEN_9889 ? phv_data_441 : _GEN_1976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1978 = 9'h1ba == _GEN_9889 ? phv_data_442 : _GEN_1977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1979 = 9'h1bb == _GEN_9889 ? phv_data_443 : _GEN_1978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1980 = 9'h1bc == _GEN_9889 ? phv_data_444 : _GEN_1979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1981 = 9'h1bd == _GEN_9889 ? phv_data_445 : _GEN_1980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1982 = 9'h1be == _GEN_9889 ? phv_data_446 : _GEN_1981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1983 = 9'h1bf == _GEN_9889 ? phv_data_447 : _GEN_1982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1984 = 9'h1c0 == _GEN_9889 ? phv_data_448 : _GEN_1983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1985 = 9'h1c1 == _GEN_9889 ? phv_data_449 : _GEN_1984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1986 = 9'h1c2 == _GEN_9889 ? phv_data_450 : _GEN_1985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1987 = 9'h1c3 == _GEN_9889 ? phv_data_451 : _GEN_1986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1988 = 9'h1c4 == _GEN_9889 ? phv_data_452 : _GEN_1987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1989 = 9'h1c5 == _GEN_9889 ? phv_data_453 : _GEN_1988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1990 = 9'h1c6 == _GEN_9889 ? phv_data_454 : _GEN_1989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1991 = 9'h1c7 == _GEN_9889 ? phv_data_455 : _GEN_1990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1992 = 9'h1c8 == _GEN_9889 ? phv_data_456 : _GEN_1991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1993 = 9'h1c9 == _GEN_9889 ? phv_data_457 : _GEN_1992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1994 = 9'h1ca == _GEN_9889 ? phv_data_458 : _GEN_1993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1995 = 9'h1cb == _GEN_9889 ? phv_data_459 : _GEN_1994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1996 = 9'h1cc == _GEN_9889 ? phv_data_460 : _GEN_1995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1997 = 9'h1cd == _GEN_9889 ? phv_data_461 : _GEN_1996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1998 = 9'h1ce == _GEN_9889 ? phv_data_462 : _GEN_1997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_1999 = 9'h1cf == _GEN_9889 ? phv_data_463 : _GEN_1998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2000 = 9'h1d0 == _GEN_9889 ? phv_data_464 : _GEN_1999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2001 = 9'h1d1 == _GEN_9889 ? phv_data_465 : _GEN_2000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2002 = 9'h1d2 == _GEN_9889 ? phv_data_466 : _GEN_2001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2003 = 9'h1d3 == _GEN_9889 ? phv_data_467 : _GEN_2002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2004 = 9'h1d4 == _GEN_9889 ? phv_data_468 : _GEN_2003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2005 = 9'h1d5 == _GEN_9889 ? phv_data_469 : _GEN_2004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2006 = 9'h1d6 == _GEN_9889 ? phv_data_470 : _GEN_2005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2007 = 9'h1d7 == _GEN_9889 ? phv_data_471 : _GEN_2006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2008 = 9'h1d8 == _GEN_9889 ? phv_data_472 : _GEN_2007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2009 = 9'h1d9 == _GEN_9889 ? phv_data_473 : _GEN_2008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2010 = 9'h1da == _GEN_9889 ? phv_data_474 : _GEN_2009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2011 = 9'h1db == _GEN_9889 ? phv_data_475 : _GEN_2010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2012 = 9'h1dc == _GEN_9889 ? phv_data_476 : _GEN_2011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2013 = 9'h1dd == _GEN_9889 ? phv_data_477 : _GEN_2012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2014 = 9'h1de == _GEN_9889 ? phv_data_478 : _GEN_2013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2015 = 9'h1df == _GEN_9889 ? phv_data_479 : _GEN_2014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2016 = 9'h1e0 == _GEN_9889 ? phv_data_480 : _GEN_2015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2017 = 9'h1e1 == _GEN_9889 ? phv_data_481 : _GEN_2016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2018 = 9'h1e2 == _GEN_9889 ? phv_data_482 : _GEN_2017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2019 = 9'h1e3 == _GEN_9889 ? phv_data_483 : _GEN_2018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2020 = 9'h1e4 == _GEN_9889 ? phv_data_484 : _GEN_2019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2021 = 9'h1e5 == _GEN_9889 ? phv_data_485 : _GEN_2020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2022 = 9'h1e6 == _GEN_9889 ? phv_data_486 : _GEN_2021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2023 = 9'h1e7 == _GEN_9889 ? phv_data_487 : _GEN_2022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2024 = 9'h1e8 == _GEN_9889 ? phv_data_488 : _GEN_2023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2025 = 9'h1e9 == _GEN_9889 ? phv_data_489 : _GEN_2024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2026 = 9'h1ea == _GEN_9889 ? phv_data_490 : _GEN_2025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2027 = 9'h1eb == _GEN_9889 ? phv_data_491 : _GEN_2026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2028 = 9'h1ec == _GEN_9889 ? phv_data_492 : _GEN_2027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2029 = 9'h1ed == _GEN_9889 ? phv_data_493 : _GEN_2028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2030 = 9'h1ee == _GEN_9889 ? phv_data_494 : _GEN_2029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2031 = 9'h1ef == _GEN_9889 ? phv_data_495 : _GEN_2030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2032 = 9'h1f0 == _GEN_9889 ? phv_data_496 : _GEN_2031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2033 = 9'h1f1 == _GEN_9889 ? phv_data_497 : _GEN_2032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2034 = 9'h1f2 == _GEN_9889 ? phv_data_498 : _GEN_2033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2035 = 9'h1f3 == _GEN_9889 ? phv_data_499 : _GEN_2034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2036 = 9'h1f4 == _GEN_9889 ? phv_data_500 : _GEN_2035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2037 = 9'h1f5 == _GEN_9889 ? phv_data_501 : _GEN_2036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2038 = 9'h1f6 == _GEN_9889 ? phv_data_502 : _GEN_2037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2039 = 9'h1f7 == _GEN_9889 ? phv_data_503 : _GEN_2038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2040 = 9'h1f8 == _GEN_9889 ? phv_data_504 : _GEN_2039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2041 = 9'h1f9 == _GEN_9889 ? phv_data_505 : _GEN_2040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2042 = 9'h1fa == _GEN_9889 ? phv_data_506 : _GEN_2041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2043 = 9'h1fb == _GEN_9889 ? phv_data_507 : _GEN_2042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2044 = 9'h1fc == _GEN_9889 ? phv_data_508 : _GEN_2043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2045 = 9'h1fd == _GEN_9889 ? phv_data_509 : _GEN_2044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2046 = 9'h1fe == _GEN_9889 ? phv_data_510 : _GEN_2045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes__0 = 9'h1ff == _GEN_9889 ? phv_data_511 : _GEN_2046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_0_T = {bytes__0,bytes__1,bytes__2,bytes__3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_0_T = {_mask_3_T_3,mask__1,mask__2,mask__3}; // @[Cat.scala 30:58]
  wire [2:0] args_offset = io_field_out_0_lo[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length = io_field_out_0_lo[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _local_offset_T_1 = {{1'd0}, args_offset}; // @[executor.scala 222:61]
  wire [2:0] local_offset = _local_offset_T_1[2:0]; // @[executor.scala 222:61]
  wire [7:0] _GEN_2049 = 3'h1 == local_offset ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2050 = 3'h2 == local_offset ? args_2 : _GEN_2049; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2051 = 3'h3 == local_offset ? args_3 : _GEN_2050; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2052 = 3'h4 == local_offset ? args_4 : _GEN_2051; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2053 = 3'h5 == local_offset ? args_5 : _GEN_2052; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2054 = 3'h6 == local_offset ? args_6 : _GEN_2053; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2055 = 3'h1 == args_length ? _GEN_2054 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [2:0] local_offset_1 = 3'h1 + args_offset; // @[executor.scala 222:61]
  wire [7:0] _GEN_2057 = 3'h1 == local_offset_1 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2058 = 3'h2 == local_offset_1 ? args_2 : _GEN_2057; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2059 = 3'h3 == local_offset_1 ? args_3 : _GEN_2058; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2060 = 3'h4 == local_offset_1 ? args_4 : _GEN_2059; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2061 = 3'h5 == local_offset_1 ? args_5 : _GEN_2060; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2062 = 3'h6 == local_offset_1 ? args_6 : _GEN_2061; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2063 = 3'h2 == args_length ? _GEN_2062 : _GEN_2055; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_2 = 3'h2 + args_offset; // @[executor.scala 222:61]
  wire [7:0] _GEN_2065 = 3'h1 == local_offset_2 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2066 = 3'h2 == local_offset_2 ? args_2 : _GEN_2065; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2067 = 3'h3 == local_offset_2 ? args_3 : _GEN_2066; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2068 = 3'h4 == local_offset_2 ? args_4 : _GEN_2067; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2069 = 3'h5 == local_offset_2 ? args_5 : _GEN_2068; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2070 = 3'h6 == local_offset_2 ? args_6 : _GEN_2069; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2071 = 3'h3 == args_length ? _GEN_2070 : _GEN_2063; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_3 = 3'h3 + args_offset; // @[executor.scala 222:61]
  wire [7:0] _GEN_2073 = 3'h1 == local_offset_3 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2074 = 3'h2 == local_offset_3 ? args_2 : _GEN_2073; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2075 = 3'h3 == local_offset_3 ? args_3 : _GEN_2074; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2076 = 3'h4 == local_offset_3 ? args_4 : _GEN_2075; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2077 = 3'h5 == local_offset_3 ? args_5 : _GEN_2076; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2078 = 3'h6 == local_offset_3 ? args_6 : _GEN_2077; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2079 = 3'h4 == args_length ? _GEN_2078 : _GEN_2071; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_4 = 3'h4 + args_offset; // @[executor.scala 222:61]
  wire [7:0] _GEN_2081 = 3'h1 == local_offset_4 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2082 = 3'h2 == local_offset_4 ? args_2 : _GEN_2081; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2083 = 3'h3 == local_offset_4 ? args_3 : _GEN_2082; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2084 = 3'h4 == local_offset_4 ? args_4 : _GEN_2083; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2085 = 3'h5 == local_offset_4 ? args_5 : _GEN_2084; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2086 = 3'h6 == local_offset_4 ? args_6 : _GEN_2085; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2087 = 3'h5 == args_length ? _GEN_2086 : _GEN_2079; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_5 = 3'h5 + args_offset; // @[executor.scala 222:61]
  wire [7:0] _GEN_2089 = 3'h1 == local_offset_5 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2090 = 3'h2 == local_offset_5 ? args_2 : _GEN_2089; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2091 = 3'h3 == local_offset_5 ? args_3 : _GEN_2090; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2092 = 3'h4 == local_offset_5 ? args_4 : _GEN_2091; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2093 = 3'h5 == local_offset_5 ? args_5 : _GEN_2092; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2094 = 3'h6 == local_offset_5 ? args_6 : _GEN_2093; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2095 = 3'h6 == args_length ? _GEN_2094 : _GEN_2087; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_6 = 3'h6 + args_offset; // @[executor.scala 222:61]
  wire [7:0] _GEN_2097 = 3'h1 == local_offset_6 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2098 = 3'h2 == local_offset_6 ? args_2 : _GEN_2097; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2099 = 3'h3 == local_offset_6 ? args_3 : _GEN_2098; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2100 = 3'h4 == local_offset_6 ? args_4 : _GEN_2099; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2101 = 3'h5 == local_offset_6 ? args_5 : _GEN_2100; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_2102 = 3'h6 == local_offset_6 ? args_6 : _GEN_2101; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] field_bytes_1_0 = 3'h7 == args_length ? _GEN_2102 : _GEN_2095; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2111 = 3'h2 == args_length ? _GEN_2054 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_2119 = 3'h3 == args_length ? _GEN_2062 : _GEN_2111; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2127 = 3'h4 == args_length ? _GEN_2070 : _GEN_2119; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2135 = 3'h5 == args_length ? _GEN_2078 : _GEN_2127; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2143 = 3'h6 == args_length ? _GEN_2086 : _GEN_2135; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2151 = 3'h7 == args_length ? _GEN_2094 : _GEN_2143; // @[executor.scala 223:66 executor.scala 224:52]
  wire [3:0] _GEN_10145 = {{1'd0}, args_length}; // @[executor.scala 223:49]
  wire [7:0] field_bytes_1_1 = 4'h8 == _GEN_10145 ? _GEN_2102 : _GEN_2151; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2167 = 3'h3 == args_length ? _GEN_2054 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_2175 = 3'h4 == args_length ? _GEN_2062 : _GEN_2167; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2183 = 3'h5 == args_length ? _GEN_2070 : _GEN_2175; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2191 = 3'h6 == args_length ? _GEN_2078 : _GEN_2183; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2199 = 3'h7 == args_length ? _GEN_2086 : _GEN_2191; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2207 = 4'h8 == _GEN_10145 ? _GEN_2094 : _GEN_2199; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_1_2 = 4'h9 == _GEN_10145 ? _GEN_2102 : _GEN_2207; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2223 = 3'h4 == args_length ? _GEN_2054 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_2231 = 3'h5 == args_length ? _GEN_2062 : _GEN_2223; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2239 = 3'h6 == args_length ? _GEN_2070 : _GEN_2231; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2247 = 3'h7 == args_length ? _GEN_2078 : _GEN_2239; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2255 = 4'h8 == _GEN_10145 ? _GEN_2086 : _GEN_2247; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_2263 = 4'h9 == _GEN_10145 ? _GEN_2094 : _GEN_2255; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_1_3 = 4'ha == _GEN_10145 ? _GEN_2102 : _GEN_2263; // @[executor.scala 223:66 executor.scala 224:52]
  wire [31:0] _io_field_out_0_T_1 = {field_bytes_1_0,field_bytes_1_1,field_bytes_1_2,field_bytes_1_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2272 = 4'ha == opcode ? _io_field_out_0_T_1 : 32'h0; // @[executor.scala 207:55 executor.scala 228:41 executor.scala 172:29]
  wire [17:0] io_field_out_0_hi_4 = io_field_out_0_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_0_T_4 = {io_field_out_0_hi_4,io_field_out_0_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_2273 = 4'hb == opcode ? _io_field_out_0_T_4 : _GEN_2272; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_2274 = from_header ? bias : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_2275 = from_header ? _io_field_out_0_T : _GEN_2273; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_2276 = from_header ? _io_mask_out_0_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  wire [3:0] opcode_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_1_lo = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire  from_header_1 = length_1 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi_1 = offset_1[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_3 = offset_1 + length_1; // @[executor.scala 193:46]
  wire [1:0] ending_1 = _ending_T_3[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_10151 = {{2'd0}, ending_1}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_3 = 4'h4 - _GEN_10151; // @[executor.scala 194:45]
  wire [1:0] bias_1 = _bias_T_3[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset_4 = {total_offset_hi_1,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2281 = 8'h1 == total_offset_4 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2282 = 8'h2 == total_offset_4 ? phv_data_2 : _GEN_2281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2283 = 8'h3 == total_offset_4 ? phv_data_3 : _GEN_2282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2284 = 8'h4 == total_offset_4 ? phv_data_4 : _GEN_2283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2285 = 8'h5 == total_offset_4 ? phv_data_5 : _GEN_2284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2286 = 8'h6 == total_offset_4 ? phv_data_6 : _GEN_2285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2287 = 8'h7 == total_offset_4 ? phv_data_7 : _GEN_2286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2288 = 8'h8 == total_offset_4 ? phv_data_8 : _GEN_2287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2289 = 8'h9 == total_offset_4 ? phv_data_9 : _GEN_2288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2290 = 8'ha == total_offset_4 ? phv_data_10 : _GEN_2289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2291 = 8'hb == total_offset_4 ? phv_data_11 : _GEN_2290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2292 = 8'hc == total_offset_4 ? phv_data_12 : _GEN_2291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2293 = 8'hd == total_offset_4 ? phv_data_13 : _GEN_2292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2294 = 8'he == total_offset_4 ? phv_data_14 : _GEN_2293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2295 = 8'hf == total_offset_4 ? phv_data_15 : _GEN_2294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2296 = 8'h10 == total_offset_4 ? phv_data_16 : _GEN_2295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2297 = 8'h11 == total_offset_4 ? phv_data_17 : _GEN_2296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2298 = 8'h12 == total_offset_4 ? phv_data_18 : _GEN_2297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2299 = 8'h13 == total_offset_4 ? phv_data_19 : _GEN_2298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2300 = 8'h14 == total_offset_4 ? phv_data_20 : _GEN_2299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2301 = 8'h15 == total_offset_4 ? phv_data_21 : _GEN_2300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2302 = 8'h16 == total_offset_4 ? phv_data_22 : _GEN_2301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2303 = 8'h17 == total_offset_4 ? phv_data_23 : _GEN_2302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2304 = 8'h18 == total_offset_4 ? phv_data_24 : _GEN_2303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2305 = 8'h19 == total_offset_4 ? phv_data_25 : _GEN_2304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2306 = 8'h1a == total_offset_4 ? phv_data_26 : _GEN_2305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2307 = 8'h1b == total_offset_4 ? phv_data_27 : _GEN_2306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2308 = 8'h1c == total_offset_4 ? phv_data_28 : _GEN_2307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2309 = 8'h1d == total_offset_4 ? phv_data_29 : _GEN_2308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2310 = 8'h1e == total_offset_4 ? phv_data_30 : _GEN_2309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2311 = 8'h1f == total_offset_4 ? phv_data_31 : _GEN_2310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2312 = 8'h20 == total_offset_4 ? phv_data_32 : _GEN_2311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2313 = 8'h21 == total_offset_4 ? phv_data_33 : _GEN_2312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2314 = 8'h22 == total_offset_4 ? phv_data_34 : _GEN_2313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2315 = 8'h23 == total_offset_4 ? phv_data_35 : _GEN_2314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2316 = 8'h24 == total_offset_4 ? phv_data_36 : _GEN_2315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2317 = 8'h25 == total_offset_4 ? phv_data_37 : _GEN_2316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2318 = 8'h26 == total_offset_4 ? phv_data_38 : _GEN_2317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2319 = 8'h27 == total_offset_4 ? phv_data_39 : _GEN_2318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2320 = 8'h28 == total_offset_4 ? phv_data_40 : _GEN_2319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2321 = 8'h29 == total_offset_4 ? phv_data_41 : _GEN_2320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2322 = 8'h2a == total_offset_4 ? phv_data_42 : _GEN_2321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2323 = 8'h2b == total_offset_4 ? phv_data_43 : _GEN_2322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2324 = 8'h2c == total_offset_4 ? phv_data_44 : _GEN_2323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2325 = 8'h2d == total_offset_4 ? phv_data_45 : _GEN_2324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2326 = 8'h2e == total_offset_4 ? phv_data_46 : _GEN_2325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2327 = 8'h2f == total_offset_4 ? phv_data_47 : _GEN_2326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2328 = 8'h30 == total_offset_4 ? phv_data_48 : _GEN_2327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2329 = 8'h31 == total_offset_4 ? phv_data_49 : _GEN_2328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2330 = 8'h32 == total_offset_4 ? phv_data_50 : _GEN_2329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2331 = 8'h33 == total_offset_4 ? phv_data_51 : _GEN_2330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2332 = 8'h34 == total_offset_4 ? phv_data_52 : _GEN_2331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2333 = 8'h35 == total_offset_4 ? phv_data_53 : _GEN_2332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2334 = 8'h36 == total_offset_4 ? phv_data_54 : _GEN_2333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2335 = 8'h37 == total_offset_4 ? phv_data_55 : _GEN_2334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2336 = 8'h38 == total_offset_4 ? phv_data_56 : _GEN_2335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2337 = 8'h39 == total_offset_4 ? phv_data_57 : _GEN_2336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2338 = 8'h3a == total_offset_4 ? phv_data_58 : _GEN_2337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2339 = 8'h3b == total_offset_4 ? phv_data_59 : _GEN_2338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2340 = 8'h3c == total_offset_4 ? phv_data_60 : _GEN_2339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2341 = 8'h3d == total_offset_4 ? phv_data_61 : _GEN_2340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2342 = 8'h3e == total_offset_4 ? phv_data_62 : _GEN_2341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2343 = 8'h3f == total_offset_4 ? phv_data_63 : _GEN_2342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2344 = 8'h40 == total_offset_4 ? phv_data_64 : _GEN_2343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2345 = 8'h41 == total_offset_4 ? phv_data_65 : _GEN_2344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2346 = 8'h42 == total_offset_4 ? phv_data_66 : _GEN_2345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2347 = 8'h43 == total_offset_4 ? phv_data_67 : _GEN_2346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2348 = 8'h44 == total_offset_4 ? phv_data_68 : _GEN_2347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2349 = 8'h45 == total_offset_4 ? phv_data_69 : _GEN_2348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2350 = 8'h46 == total_offset_4 ? phv_data_70 : _GEN_2349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2351 = 8'h47 == total_offset_4 ? phv_data_71 : _GEN_2350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2352 = 8'h48 == total_offset_4 ? phv_data_72 : _GEN_2351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2353 = 8'h49 == total_offset_4 ? phv_data_73 : _GEN_2352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2354 = 8'h4a == total_offset_4 ? phv_data_74 : _GEN_2353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2355 = 8'h4b == total_offset_4 ? phv_data_75 : _GEN_2354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2356 = 8'h4c == total_offset_4 ? phv_data_76 : _GEN_2355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2357 = 8'h4d == total_offset_4 ? phv_data_77 : _GEN_2356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2358 = 8'h4e == total_offset_4 ? phv_data_78 : _GEN_2357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2359 = 8'h4f == total_offset_4 ? phv_data_79 : _GEN_2358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2360 = 8'h50 == total_offset_4 ? phv_data_80 : _GEN_2359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2361 = 8'h51 == total_offset_4 ? phv_data_81 : _GEN_2360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2362 = 8'h52 == total_offset_4 ? phv_data_82 : _GEN_2361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2363 = 8'h53 == total_offset_4 ? phv_data_83 : _GEN_2362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2364 = 8'h54 == total_offset_4 ? phv_data_84 : _GEN_2363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2365 = 8'h55 == total_offset_4 ? phv_data_85 : _GEN_2364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2366 = 8'h56 == total_offset_4 ? phv_data_86 : _GEN_2365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2367 = 8'h57 == total_offset_4 ? phv_data_87 : _GEN_2366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2368 = 8'h58 == total_offset_4 ? phv_data_88 : _GEN_2367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2369 = 8'h59 == total_offset_4 ? phv_data_89 : _GEN_2368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2370 = 8'h5a == total_offset_4 ? phv_data_90 : _GEN_2369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2371 = 8'h5b == total_offset_4 ? phv_data_91 : _GEN_2370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2372 = 8'h5c == total_offset_4 ? phv_data_92 : _GEN_2371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2373 = 8'h5d == total_offset_4 ? phv_data_93 : _GEN_2372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2374 = 8'h5e == total_offset_4 ? phv_data_94 : _GEN_2373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2375 = 8'h5f == total_offset_4 ? phv_data_95 : _GEN_2374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2376 = 8'h60 == total_offset_4 ? phv_data_96 : _GEN_2375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2377 = 8'h61 == total_offset_4 ? phv_data_97 : _GEN_2376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2378 = 8'h62 == total_offset_4 ? phv_data_98 : _GEN_2377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2379 = 8'h63 == total_offset_4 ? phv_data_99 : _GEN_2378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2380 = 8'h64 == total_offset_4 ? phv_data_100 : _GEN_2379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2381 = 8'h65 == total_offset_4 ? phv_data_101 : _GEN_2380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2382 = 8'h66 == total_offset_4 ? phv_data_102 : _GEN_2381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2383 = 8'h67 == total_offset_4 ? phv_data_103 : _GEN_2382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2384 = 8'h68 == total_offset_4 ? phv_data_104 : _GEN_2383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2385 = 8'h69 == total_offset_4 ? phv_data_105 : _GEN_2384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2386 = 8'h6a == total_offset_4 ? phv_data_106 : _GEN_2385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2387 = 8'h6b == total_offset_4 ? phv_data_107 : _GEN_2386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2388 = 8'h6c == total_offset_4 ? phv_data_108 : _GEN_2387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2389 = 8'h6d == total_offset_4 ? phv_data_109 : _GEN_2388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2390 = 8'h6e == total_offset_4 ? phv_data_110 : _GEN_2389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2391 = 8'h6f == total_offset_4 ? phv_data_111 : _GEN_2390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2392 = 8'h70 == total_offset_4 ? phv_data_112 : _GEN_2391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2393 = 8'h71 == total_offset_4 ? phv_data_113 : _GEN_2392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2394 = 8'h72 == total_offset_4 ? phv_data_114 : _GEN_2393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2395 = 8'h73 == total_offset_4 ? phv_data_115 : _GEN_2394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2396 = 8'h74 == total_offset_4 ? phv_data_116 : _GEN_2395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2397 = 8'h75 == total_offset_4 ? phv_data_117 : _GEN_2396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2398 = 8'h76 == total_offset_4 ? phv_data_118 : _GEN_2397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2399 = 8'h77 == total_offset_4 ? phv_data_119 : _GEN_2398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2400 = 8'h78 == total_offset_4 ? phv_data_120 : _GEN_2399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2401 = 8'h79 == total_offset_4 ? phv_data_121 : _GEN_2400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2402 = 8'h7a == total_offset_4 ? phv_data_122 : _GEN_2401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2403 = 8'h7b == total_offset_4 ? phv_data_123 : _GEN_2402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2404 = 8'h7c == total_offset_4 ? phv_data_124 : _GEN_2403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2405 = 8'h7d == total_offset_4 ? phv_data_125 : _GEN_2404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2406 = 8'h7e == total_offset_4 ? phv_data_126 : _GEN_2405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2407 = 8'h7f == total_offset_4 ? phv_data_127 : _GEN_2406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2408 = 8'h80 == total_offset_4 ? phv_data_128 : _GEN_2407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2409 = 8'h81 == total_offset_4 ? phv_data_129 : _GEN_2408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2410 = 8'h82 == total_offset_4 ? phv_data_130 : _GEN_2409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2411 = 8'h83 == total_offset_4 ? phv_data_131 : _GEN_2410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2412 = 8'h84 == total_offset_4 ? phv_data_132 : _GEN_2411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2413 = 8'h85 == total_offset_4 ? phv_data_133 : _GEN_2412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2414 = 8'h86 == total_offset_4 ? phv_data_134 : _GEN_2413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2415 = 8'h87 == total_offset_4 ? phv_data_135 : _GEN_2414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2416 = 8'h88 == total_offset_4 ? phv_data_136 : _GEN_2415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2417 = 8'h89 == total_offset_4 ? phv_data_137 : _GEN_2416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2418 = 8'h8a == total_offset_4 ? phv_data_138 : _GEN_2417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2419 = 8'h8b == total_offset_4 ? phv_data_139 : _GEN_2418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2420 = 8'h8c == total_offset_4 ? phv_data_140 : _GEN_2419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2421 = 8'h8d == total_offset_4 ? phv_data_141 : _GEN_2420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2422 = 8'h8e == total_offset_4 ? phv_data_142 : _GEN_2421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2423 = 8'h8f == total_offset_4 ? phv_data_143 : _GEN_2422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2424 = 8'h90 == total_offset_4 ? phv_data_144 : _GEN_2423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2425 = 8'h91 == total_offset_4 ? phv_data_145 : _GEN_2424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2426 = 8'h92 == total_offset_4 ? phv_data_146 : _GEN_2425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2427 = 8'h93 == total_offset_4 ? phv_data_147 : _GEN_2426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2428 = 8'h94 == total_offset_4 ? phv_data_148 : _GEN_2427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2429 = 8'h95 == total_offset_4 ? phv_data_149 : _GEN_2428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2430 = 8'h96 == total_offset_4 ? phv_data_150 : _GEN_2429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2431 = 8'h97 == total_offset_4 ? phv_data_151 : _GEN_2430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2432 = 8'h98 == total_offset_4 ? phv_data_152 : _GEN_2431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2433 = 8'h99 == total_offset_4 ? phv_data_153 : _GEN_2432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2434 = 8'h9a == total_offset_4 ? phv_data_154 : _GEN_2433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2435 = 8'h9b == total_offset_4 ? phv_data_155 : _GEN_2434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2436 = 8'h9c == total_offset_4 ? phv_data_156 : _GEN_2435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2437 = 8'h9d == total_offset_4 ? phv_data_157 : _GEN_2436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2438 = 8'h9e == total_offset_4 ? phv_data_158 : _GEN_2437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2439 = 8'h9f == total_offset_4 ? phv_data_159 : _GEN_2438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2440 = 8'ha0 == total_offset_4 ? phv_data_160 : _GEN_2439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2441 = 8'ha1 == total_offset_4 ? phv_data_161 : _GEN_2440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2442 = 8'ha2 == total_offset_4 ? phv_data_162 : _GEN_2441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2443 = 8'ha3 == total_offset_4 ? phv_data_163 : _GEN_2442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2444 = 8'ha4 == total_offset_4 ? phv_data_164 : _GEN_2443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2445 = 8'ha5 == total_offset_4 ? phv_data_165 : _GEN_2444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2446 = 8'ha6 == total_offset_4 ? phv_data_166 : _GEN_2445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2447 = 8'ha7 == total_offset_4 ? phv_data_167 : _GEN_2446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2448 = 8'ha8 == total_offset_4 ? phv_data_168 : _GEN_2447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2449 = 8'ha9 == total_offset_4 ? phv_data_169 : _GEN_2448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2450 = 8'haa == total_offset_4 ? phv_data_170 : _GEN_2449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2451 = 8'hab == total_offset_4 ? phv_data_171 : _GEN_2450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2452 = 8'hac == total_offset_4 ? phv_data_172 : _GEN_2451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2453 = 8'had == total_offset_4 ? phv_data_173 : _GEN_2452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2454 = 8'hae == total_offset_4 ? phv_data_174 : _GEN_2453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2455 = 8'haf == total_offset_4 ? phv_data_175 : _GEN_2454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2456 = 8'hb0 == total_offset_4 ? phv_data_176 : _GEN_2455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2457 = 8'hb1 == total_offset_4 ? phv_data_177 : _GEN_2456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2458 = 8'hb2 == total_offset_4 ? phv_data_178 : _GEN_2457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2459 = 8'hb3 == total_offset_4 ? phv_data_179 : _GEN_2458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2460 = 8'hb4 == total_offset_4 ? phv_data_180 : _GEN_2459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2461 = 8'hb5 == total_offset_4 ? phv_data_181 : _GEN_2460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2462 = 8'hb6 == total_offset_4 ? phv_data_182 : _GEN_2461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2463 = 8'hb7 == total_offset_4 ? phv_data_183 : _GEN_2462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2464 = 8'hb8 == total_offset_4 ? phv_data_184 : _GEN_2463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2465 = 8'hb9 == total_offset_4 ? phv_data_185 : _GEN_2464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2466 = 8'hba == total_offset_4 ? phv_data_186 : _GEN_2465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2467 = 8'hbb == total_offset_4 ? phv_data_187 : _GEN_2466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2468 = 8'hbc == total_offset_4 ? phv_data_188 : _GEN_2467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2469 = 8'hbd == total_offset_4 ? phv_data_189 : _GEN_2468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2470 = 8'hbe == total_offset_4 ? phv_data_190 : _GEN_2469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2471 = 8'hbf == total_offset_4 ? phv_data_191 : _GEN_2470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2472 = 8'hc0 == total_offset_4 ? phv_data_192 : _GEN_2471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2473 = 8'hc1 == total_offset_4 ? phv_data_193 : _GEN_2472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2474 = 8'hc2 == total_offset_4 ? phv_data_194 : _GEN_2473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2475 = 8'hc3 == total_offset_4 ? phv_data_195 : _GEN_2474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2476 = 8'hc4 == total_offset_4 ? phv_data_196 : _GEN_2475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2477 = 8'hc5 == total_offset_4 ? phv_data_197 : _GEN_2476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2478 = 8'hc6 == total_offset_4 ? phv_data_198 : _GEN_2477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2479 = 8'hc7 == total_offset_4 ? phv_data_199 : _GEN_2478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2480 = 8'hc8 == total_offset_4 ? phv_data_200 : _GEN_2479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2481 = 8'hc9 == total_offset_4 ? phv_data_201 : _GEN_2480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2482 = 8'hca == total_offset_4 ? phv_data_202 : _GEN_2481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2483 = 8'hcb == total_offset_4 ? phv_data_203 : _GEN_2482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2484 = 8'hcc == total_offset_4 ? phv_data_204 : _GEN_2483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2485 = 8'hcd == total_offset_4 ? phv_data_205 : _GEN_2484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2486 = 8'hce == total_offset_4 ? phv_data_206 : _GEN_2485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2487 = 8'hcf == total_offset_4 ? phv_data_207 : _GEN_2486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2488 = 8'hd0 == total_offset_4 ? phv_data_208 : _GEN_2487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2489 = 8'hd1 == total_offset_4 ? phv_data_209 : _GEN_2488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2490 = 8'hd2 == total_offset_4 ? phv_data_210 : _GEN_2489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2491 = 8'hd3 == total_offset_4 ? phv_data_211 : _GEN_2490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2492 = 8'hd4 == total_offset_4 ? phv_data_212 : _GEN_2491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2493 = 8'hd5 == total_offset_4 ? phv_data_213 : _GEN_2492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2494 = 8'hd6 == total_offset_4 ? phv_data_214 : _GEN_2493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2495 = 8'hd7 == total_offset_4 ? phv_data_215 : _GEN_2494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2496 = 8'hd8 == total_offset_4 ? phv_data_216 : _GEN_2495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2497 = 8'hd9 == total_offset_4 ? phv_data_217 : _GEN_2496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2498 = 8'hda == total_offset_4 ? phv_data_218 : _GEN_2497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2499 = 8'hdb == total_offset_4 ? phv_data_219 : _GEN_2498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2500 = 8'hdc == total_offset_4 ? phv_data_220 : _GEN_2499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2501 = 8'hdd == total_offset_4 ? phv_data_221 : _GEN_2500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2502 = 8'hde == total_offset_4 ? phv_data_222 : _GEN_2501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2503 = 8'hdf == total_offset_4 ? phv_data_223 : _GEN_2502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2504 = 8'he0 == total_offset_4 ? phv_data_224 : _GEN_2503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2505 = 8'he1 == total_offset_4 ? phv_data_225 : _GEN_2504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2506 = 8'he2 == total_offset_4 ? phv_data_226 : _GEN_2505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2507 = 8'he3 == total_offset_4 ? phv_data_227 : _GEN_2506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2508 = 8'he4 == total_offset_4 ? phv_data_228 : _GEN_2507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2509 = 8'he5 == total_offset_4 ? phv_data_229 : _GEN_2508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2510 = 8'he6 == total_offset_4 ? phv_data_230 : _GEN_2509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2511 = 8'he7 == total_offset_4 ? phv_data_231 : _GEN_2510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2512 = 8'he8 == total_offset_4 ? phv_data_232 : _GEN_2511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2513 = 8'he9 == total_offset_4 ? phv_data_233 : _GEN_2512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2514 = 8'hea == total_offset_4 ? phv_data_234 : _GEN_2513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2515 = 8'heb == total_offset_4 ? phv_data_235 : _GEN_2514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2516 = 8'hec == total_offset_4 ? phv_data_236 : _GEN_2515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2517 = 8'hed == total_offset_4 ? phv_data_237 : _GEN_2516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2518 = 8'hee == total_offset_4 ? phv_data_238 : _GEN_2517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2519 = 8'hef == total_offset_4 ? phv_data_239 : _GEN_2518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2520 = 8'hf0 == total_offset_4 ? phv_data_240 : _GEN_2519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2521 = 8'hf1 == total_offset_4 ? phv_data_241 : _GEN_2520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2522 = 8'hf2 == total_offset_4 ? phv_data_242 : _GEN_2521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2523 = 8'hf3 == total_offset_4 ? phv_data_243 : _GEN_2522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2524 = 8'hf4 == total_offset_4 ? phv_data_244 : _GEN_2523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2525 = 8'hf5 == total_offset_4 ? phv_data_245 : _GEN_2524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2526 = 8'hf6 == total_offset_4 ? phv_data_246 : _GEN_2525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2527 = 8'hf7 == total_offset_4 ? phv_data_247 : _GEN_2526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2528 = 8'hf8 == total_offset_4 ? phv_data_248 : _GEN_2527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2529 = 8'hf9 == total_offset_4 ? phv_data_249 : _GEN_2528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2530 = 8'hfa == total_offset_4 ? phv_data_250 : _GEN_2529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2531 = 8'hfb == total_offset_4 ? phv_data_251 : _GEN_2530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2532 = 8'hfc == total_offset_4 ? phv_data_252 : _GEN_2531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2533 = 8'hfd == total_offset_4 ? phv_data_253 : _GEN_2532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2534 = 8'hfe == total_offset_4 ? phv_data_254 : _GEN_2533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2535 = 8'hff == total_offset_4 ? phv_data_255 : _GEN_2534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_10152 = {{1'd0}, total_offset_4}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2536 = 9'h100 == _GEN_10152 ? phv_data_256 : _GEN_2535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2537 = 9'h101 == _GEN_10152 ? phv_data_257 : _GEN_2536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2538 = 9'h102 == _GEN_10152 ? phv_data_258 : _GEN_2537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2539 = 9'h103 == _GEN_10152 ? phv_data_259 : _GEN_2538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2540 = 9'h104 == _GEN_10152 ? phv_data_260 : _GEN_2539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2541 = 9'h105 == _GEN_10152 ? phv_data_261 : _GEN_2540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2542 = 9'h106 == _GEN_10152 ? phv_data_262 : _GEN_2541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2543 = 9'h107 == _GEN_10152 ? phv_data_263 : _GEN_2542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2544 = 9'h108 == _GEN_10152 ? phv_data_264 : _GEN_2543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2545 = 9'h109 == _GEN_10152 ? phv_data_265 : _GEN_2544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2546 = 9'h10a == _GEN_10152 ? phv_data_266 : _GEN_2545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2547 = 9'h10b == _GEN_10152 ? phv_data_267 : _GEN_2546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2548 = 9'h10c == _GEN_10152 ? phv_data_268 : _GEN_2547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2549 = 9'h10d == _GEN_10152 ? phv_data_269 : _GEN_2548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2550 = 9'h10e == _GEN_10152 ? phv_data_270 : _GEN_2549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2551 = 9'h10f == _GEN_10152 ? phv_data_271 : _GEN_2550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2552 = 9'h110 == _GEN_10152 ? phv_data_272 : _GEN_2551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2553 = 9'h111 == _GEN_10152 ? phv_data_273 : _GEN_2552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2554 = 9'h112 == _GEN_10152 ? phv_data_274 : _GEN_2553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2555 = 9'h113 == _GEN_10152 ? phv_data_275 : _GEN_2554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2556 = 9'h114 == _GEN_10152 ? phv_data_276 : _GEN_2555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2557 = 9'h115 == _GEN_10152 ? phv_data_277 : _GEN_2556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2558 = 9'h116 == _GEN_10152 ? phv_data_278 : _GEN_2557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2559 = 9'h117 == _GEN_10152 ? phv_data_279 : _GEN_2558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2560 = 9'h118 == _GEN_10152 ? phv_data_280 : _GEN_2559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2561 = 9'h119 == _GEN_10152 ? phv_data_281 : _GEN_2560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2562 = 9'h11a == _GEN_10152 ? phv_data_282 : _GEN_2561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2563 = 9'h11b == _GEN_10152 ? phv_data_283 : _GEN_2562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2564 = 9'h11c == _GEN_10152 ? phv_data_284 : _GEN_2563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2565 = 9'h11d == _GEN_10152 ? phv_data_285 : _GEN_2564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2566 = 9'h11e == _GEN_10152 ? phv_data_286 : _GEN_2565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2567 = 9'h11f == _GEN_10152 ? phv_data_287 : _GEN_2566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2568 = 9'h120 == _GEN_10152 ? phv_data_288 : _GEN_2567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2569 = 9'h121 == _GEN_10152 ? phv_data_289 : _GEN_2568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2570 = 9'h122 == _GEN_10152 ? phv_data_290 : _GEN_2569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2571 = 9'h123 == _GEN_10152 ? phv_data_291 : _GEN_2570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2572 = 9'h124 == _GEN_10152 ? phv_data_292 : _GEN_2571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2573 = 9'h125 == _GEN_10152 ? phv_data_293 : _GEN_2572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2574 = 9'h126 == _GEN_10152 ? phv_data_294 : _GEN_2573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2575 = 9'h127 == _GEN_10152 ? phv_data_295 : _GEN_2574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2576 = 9'h128 == _GEN_10152 ? phv_data_296 : _GEN_2575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2577 = 9'h129 == _GEN_10152 ? phv_data_297 : _GEN_2576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2578 = 9'h12a == _GEN_10152 ? phv_data_298 : _GEN_2577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2579 = 9'h12b == _GEN_10152 ? phv_data_299 : _GEN_2578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2580 = 9'h12c == _GEN_10152 ? phv_data_300 : _GEN_2579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2581 = 9'h12d == _GEN_10152 ? phv_data_301 : _GEN_2580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2582 = 9'h12e == _GEN_10152 ? phv_data_302 : _GEN_2581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2583 = 9'h12f == _GEN_10152 ? phv_data_303 : _GEN_2582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2584 = 9'h130 == _GEN_10152 ? phv_data_304 : _GEN_2583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2585 = 9'h131 == _GEN_10152 ? phv_data_305 : _GEN_2584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2586 = 9'h132 == _GEN_10152 ? phv_data_306 : _GEN_2585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2587 = 9'h133 == _GEN_10152 ? phv_data_307 : _GEN_2586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2588 = 9'h134 == _GEN_10152 ? phv_data_308 : _GEN_2587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2589 = 9'h135 == _GEN_10152 ? phv_data_309 : _GEN_2588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2590 = 9'h136 == _GEN_10152 ? phv_data_310 : _GEN_2589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2591 = 9'h137 == _GEN_10152 ? phv_data_311 : _GEN_2590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2592 = 9'h138 == _GEN_10152 ? phv_data_312 : _GEN_2591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2593 = 9'h139 == _GEN_10152 ? phv_data_313 : _GEN_2592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2594 = 9'h13a == _GEN_10152 ? phv_data_314 : _GEN_2593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2595 = 9'h13b == _GEN_10152 ? phv_data_315 : _GEN_2594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2596 = 9'h13c == _GEN_10152 ? phv_data_316 : _GEN_2595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2597 = 9'h13d == _GEN_10152 ? phv_data_317 : _GEN_2596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2598 = 9'h13e == _GEN_10152 ? phv_data_318 : _GEN_2597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2599 = 9'h13f == _GEN_10152 ? phv_data_319 : _GEN_2598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2600 = 9'h140 == _GEN_10152 ? phv_data_320 : _GEN_2599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2601 = 9'h141 == _GEN_10152 ? phv_data_321 : _GEN_2600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2602 = 9'h142 == _GEN_10152 ? phv_data_322 : _GEN_2601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2603 = 9'h143 == _GEN_10152 ? phv_data_323 : _GEN_2602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2604 = 9'h144 == _GEN_10152 ? phv_data_324 : _GEN_2603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2605 = 9'h145 == _GEN_10152 ? phv_data_325 : _GEN_2604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2606 = 9'h146 == _GEN_10152 ? phv_data_326 : _GEN_2605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2607 = 9'h147 == _GEN_10152 ? phv_data_327 : _GEN_2606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2608 = 9'h148 == _GEN_10152 ? phv_data_328 : _GEN_2607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2609 = 9'h149 == _GEN_10152 ? phv_data_329 : _GEN_2608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2610 = 9'h14a == _GEN_10152 ? phv_data_330 : _GEN_2609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2611 = 9'h14b == _GEN_10152 ? phv_data_331 : _GEN_2610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2612 = 9'h14c == _GEN_10152 ? phv_data_332 : _GEN_2611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2613 = 9'h14d == _GEN_10152 ? phv_data_333 : _GEN_2612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2614 = 9'h14e == _GEN_10152 ? phv_data_334 : _GEN_2613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2615 = 9'h14f == _GEN_10152 ? phv_data_335 : _GEN_2614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2616 = 9'h150 == _GEN_10152 ? phv_data_336 : _GEN_2615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2617 = 9'h151 == _GEN_10152 ? phv_data_337 : _GEN_2616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2618 = 9'h152 == _GEN_10152 ? phv_data_338 : _GEN_2617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2619 = 9'h153 == _GEN_10152 ? phv_data_339 : _GEN_2618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2620 = 9'h154 == _GEN_10152 ? phv_data_340 : _GEN_2619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2621 = 9'h155 == _GEN_10152 ? phv_data_341 : _GEN_2620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2622 = 9'h156 == _GEN_10152 ? phv_data_342 : _GEN_2621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2623 = 9'h157 == _GEN_10152 ? phv_data_343 : _GEN_2622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2624 = 9'h158 == _GEN_10152 ? phv_data_344 : _GEN_2623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2625 = 9'h159 == _GEN_10152 ? phv_data_345 : _GEN_2624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2626 = 9'h15a == _GEN_10152 ? phv_data_346 : _GEN_2625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2627 = 9'h15b == _GEN_10152 ? phv_data_347 : _GEN_2626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2628 = 9'h15c == _GEN_10152 ? phv_data_348 : _GEN_2627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2629 = 9'h15d == _GEN_10152 ? phv_data_349 : _GEN_2628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2630 = 9'h15e == _GEN_10152 ? phv_data_350 : _GEN_2629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2631 = 9'h15f == _GEN_10152 ? phv_data_351 : _GEN_2630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2632 = 9'h160 == _GEN_10152 ? phv_data_352 : _GEN_2631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2633 = 9'h161 == _GEN_10152 ? phv_data_353 : _GEN_2632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2634 = 9'h162 == _GEN_10152 ? phv_data_354 : _GEN_2633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2635 = 9'h163 == _GEN_10152 ? phv_data_355 : _GEN_2634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2636 = 9'h164 == _GEN_10152 ? phv_data_356 : _GEN_2635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2637 = 9'h165 == _GEN_10152 ? phv_data_357 : _GEN_2636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2638 = 9'h166 == _GEN_10152 ? phv_data_358 : _GEN_2637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2639 = 9'h167 == _GEN_10152 ? phv_data_359 : _GEN_2638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2640 = 9'h168 == _GEN_10152 ? phv_data_360 : _GEN_2639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2641 = 9'h169 == _GEN_10152 ? phv_data_361 : _GEN_2640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2642 = 9'h16a == _GEN_10152 ? phv_data_362 : _GEN_2641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2643 = 9'h16b == _GEN_10152 ? phv_data_363 : _GEN_2642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2644 = 9'h16c == _GEN_10152 ? phv_data_364 : _GEN_2643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2645 = 9'h16d == _GEN_10152 ? phv_data_365 : _GEN_2644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2646 = 9'h16e == _GEN_10152 ? phv_data_366 : _GEN_2645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2647 = 9'h16f == _GEN_10152 ? phv_data_367 : _GEN_2646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2648 = 9'h170 == _GEN_10152 ? phv_data_368 : _GEN_2647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2649 = 9'h171 == _GEN_10152 ? phv_data_369 : _GEN_2648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2650 = 9'h172 == _GEN_10152 ? phv_data_370 : _GEN_2649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2651 = 9'h173 == _GEN_10152 ? phv_data_371 : _GEN_2650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2652 = 9'h174 == _GEN_10152 ? phv_data_372 : _GEN_2651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2653 = 9'h175 == _GEN_10152 ? phv_data_373 : _GEN_2652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2654 = 9'h176 == _GEN_10152 ? phv_data_374 : _GEN_2653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2655 = 9'h177 == _GEN_10152 ? phv_data_375 : _GEN_2654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2656 = 9'h178 == _GEN_10152 ? phv_data_376 : _GEN_2655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2657 = 9'h179 == _GEN_10152 ? phv_data_377 : _GEN_2656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2658 = 9'h17a == _GEN_10152 ? phv_data_378 : _GEN_2657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2659 = 9'h17b == _GEN_10152 ? phv_data_379 : _GEN_2658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2660 = 9'h17c == _GEN_10152 ? phv_data_380 : _GEN_2659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2661 = 9'h17d == _GEN_10152 ? phv_data_381 : _GEN_2660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2662 = 9'h17e == _GEN_10152 ? phv_data_382 : _GEN_2661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2663 = 9'h17f == _GEN_10152 ? phv_data_383 : _GEN_2662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2664 = 9'h180 == _GEN_10152 ? phv_data_384 : _GEN_2663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2665 = 9'h181 == _GEN_10152 ? phv_data_385 : _GEN_2664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2666 = 9'h182 == _GEN_10152 ? phv_data_386 : _GEN_2665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2667 = 9'h183 == _GEN_10152 ? phv_data_387 : _GEN_2666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2668 = 9'h184 == _GEN_10152 ? phv_data_388 : _GEN_2667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2669 = 9'h185 == _GEN_10152 ? phv_data_389 : _GEN_2668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2670 = 9'h186 == _GEN_10152 ? phv_data_390 : _GEN_2669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2671 = 9'h187 == _GEN_10152 ? phv_data_391 : _GEN_2670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2672 = 9'h188 == _GEN_10152 ? phv_data_392 : _GEN_2671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2673 = 9'h189 == _GEN_10152 ? phv_data_393 : _GEN_2672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2674 = 9'h18a == _GEN_10152 ? phv_data_394 : _GEN_2673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2675 = 9'h18b == _GEN_10152 ? phv_data_395 : _GEN_2674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2676 = 9'h18c == _GEN_10152 ? phv_data_396 : _GEN_2675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2677 = 9'h18d == _GEN_10152 ? phv_data_397 : _GEN_2676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2678 = 9'h18e == _GEN_10152 ? phv_data_398 : _GEN_2677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2679 = 9'h18f == _GEN_10152 ? phv_data_399 : _GEN_2678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2680 = 9'h190 == _GEN_10152 ? phv_data_400 : _GEN_2679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2681 = 9'h191 == _GEN_10152 ? phv_data_401 : _GEN_2680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2682 = 9'h192 == _GEN_10152 ? phv_data_402 : _GEN_2681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2683 = 9'h193 == _GEN_10152 ? phv_data_403 : _GEN_2682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2684 = 9'h194 == _GEN_10152 ? phv_data_404 : _GEN_2683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2685 = 9'h195 == _GEN_10152 ? phv_data_405 : _GEN_2684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2686 = 9'h196 == _GEN_10152 ? phv_data_406 : _GEN_2685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2687 = 9'h197 == _GEN_10152 ? phv_data_407 : _GEN_2686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2688 = 9'h198 == _GEN_10152 ? phv_data_408 : _GEN_2687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2689 = 9'h199 == _GEN_10152 ? phv_data_409 : _GEN_2688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2690 = 9'h19a == _GEN_10152 ? phv_data_410 : _GEN_2689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2691 = 9'h19b == _GEN_10152 ? phv_data_411 : _GEN_2690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2692 = 9'h19c == _GEN_10152 ? phv_data_412 : _GEN_2691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2693 = 9'h19d == _GEN_10152 ? phv_data_413 : _GEN_2692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2694 = 9'h19e == _GEN_10152 ? phv_data_414 : _GEN_2693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2695 = 9'h19f == _GEN_10152 ? phv_data_415 : _GEN_2694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2696 = 9'h1a0 == _GEN_10152 ? phv_data_416 : _GEN_2695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2697 = 9'h1a1 == _GEN_10152 ? phv_data_417 : _GEN_2696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2698 = 9'h1a2 == _GEN_10152 ? phv_data_418 : _GEN_2697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2699 = 9'h1a3 == _GEN_10152 ? phv_data_419 : _GEN_2698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2700 = 9'h1a4 == _GEN_10152 ? phv_data_420 : _GEN_2699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2701 = 9'h1a5 == _GEN_10152 ? phv_data_421 : _GEN_2700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2702 = 9'h1a6 == _GEN_10152 ? phv_data_422 : _GEN_2701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2703 = 9'h1a7 == _GEN_10152 ? phv_data_423 : _GEN_2702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2704 = 9'h1a8 == _GEN_10152 ? phv_data_424 : _GEN_2703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2705 = 9'h1a9 == _GEN_10152 ? phv_data_425 : _GEN_2704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2706 = 9'h1aa == _GEN_10152 ? phv_data_426 : _GEN_2705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2707 = 9'h1ab == _GEN_10152 ? phv_data_427 : _GEN_2706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2708 = 9'h1ac == _GEN_10152 ? phv_data_428 : _GEN_2707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2709 = 9'h1ad == _GEN_10152 ? phv_data_429 : _GEN_2708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2710 = 9'h1ae == _GEN_10152 ? phv_data_430 : _GEN_2709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2711 = 9'h1af == _GEN_10152 ? phv_data_431 : _GEN_2710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2712 = 9'h1b0 == _GEN_10152 ? phv_data_432 : _GEN_2711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2713 = 9'h1b1 == _GEN_10152 ? phv_data_433 : _GEN_2712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2714 = 9'h1b2 == _GEN_10152 ? phv_data_434 : _GEN_2713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2715 = 9'h1b3 == _GEN_10152 ? phv_data_435 : _GEN_2714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2716 = 9'h1b4 == _GEN_10152 ? phv_data_436 : _GEN_2715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2717 = 9'h1b5 == _GEN_10152 ? phv_data_437 : _GEN_2716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2718 = 9'h1b6 == _GEN_10152 ? phv_data_438 : _GEN_2717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2719 = 9'h1b7 == _GEN_10152 ? phv_data_439 : _GEN_2718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2720 = 9'h1b8 == _GEN_10152 ? phv_data_440 : _GEN_2719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2721 = 9'h1b9 == _GEN_10152 ? phv_data_441 : _GEN_2720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2722 = 9'h1ba == _GEN_10152 ? phv_data_442 : _GEN_2721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2723 = 9'h1bb == _GEN_10152 ? phv_data_443 : _GEN_2722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2724 = 9'h1bc == _GEN_10152 ? phv_data_444 : _GEN_2723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2725 = 9'h1bd == _GEN_10152 ? phv_data_445 : _GEN_2724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2726 = 9'h1be == _GEN_10152 ? phv_data_446 : _GEN_2725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2727 = 9'h1bf == _GEN_10152 ? phv_data_447 : _GEN_2726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2728 = 9'h1c0 == _GEN_10152 ? phv_data_448 : _GEN_2727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2729 = 9'h1c1 == _GEN_10152 ? phv_data_449 : _GEN_2728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2730 = 9'h1c2 == _GEN_10152 ? phv_data_450 : _GEN_2729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2731 = 9'h1c3 == _GEN_10152 ? phv_data_451 : _GEN_2730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2732 = 9'h1c4 == _GEN_10152 ? phv_data_452 : _GEN_2731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2733 = 9'h1c5 == _GEN_10152 ? phv_data_453 : _GEN_2732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2734 = 9'h1c6 == _GEN_10152 ? phv_data_454 : _GEN_2733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2735 = 9'h1c7 == _GEN_10152 ? phv_data_455 : _GEN_2734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2736 = 9'h1c8 == _GEN_10152 ? phv_data_456 : _GEN_2735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2737 = 9'h1c9 == _GEN_10152 ? phv_data_457 : _GEN_2736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2738 = 9'h1ca == _GEN_10152 ? phv_data_458 : _GEN_2737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2739 = 9'h1cb == _GEN_10152 ? phv_data_459 : _GEN_2738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2740 = 9'h1cc == _GEN_10152 ? phv_data_460 : _GEN_2739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2741 = 9'h1cd == _GEN_10152 ? phv_data_461 : _GEN_2740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2742 = 9'h1ce == _GEN_10152 ? phv_data_462 : _GEN_2741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2743 = 9'h1cf == _GEN_10152 ? phv_data_463 : _GEN_2742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2744 = 9'h1d0 == _GEN_10152 ? phv_data_464 : _GEN_2743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2745 = 9'h1d1 == _GEN_10152 ? phv_data_465 : _GEN_2744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2746 = 9'h1d2 == _GEN_10152 ? phv_data_466 : _GEN_2745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2747 = 9'h1d3 == _GEN_10152 ? phv_data_467 : _GEN_2746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2748 = 9'h1d4 == _GEN_10152 ? phv_data_468 : _GEN_2747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2749 = 9'h1d5 == _GEN_10152 ? phv_data_469 : _GEN_2748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2750 = 9'h1d6 == _GEN_10152 ? phv_data_470 : _GEN_2749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2751 = 9'h1d7 == _GEN_10152 ? phv_data_471 : _GEN_2750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2752 = 9'h1d8 == _GEN_10152 ? phv_data_472 : _GEN_2751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2753 = 9'h1d9 == _GEN_10152 ? phv_data_473 : _GEN_2752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2754 = 9'h1da == _GEN_10152 ? phv_data_474 : _GEN_2753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2755 = 9'h1db == _GEN_10152 ? phv_data_475 : _GEN_2754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2756 = 9'h1dc == _GEN_10152 ? phv_data_476 : _GEN_2755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2757 = 9'h1dd == _GEN_10152 ? phv_data_477 : _GEN_2756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2758 = 9'h1de == _GEN_10152 ? phv_data_478 : _GEN_2757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2759 = 9'h1df == _GEN_10152 ? phv_data_479 : _GEN_2758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2760 = 9'h1e0 == _GEN_10152 ? phv_data_480 : _GEN_2759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2761 = 9'h1e1 == _GEN_10152 ? phv_data_481 : _GEN_2760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2762 = 9'h1e2 == _GEN_10152 ? phv_data_482 : _GEN_2761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2763 = 9'h1e3 == _GEN_10152 ? phv_data_483 : _GEN_2762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2764 = 9'h1e4 == _GEN_10152 ? phv_data_484 : _GEN_2763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2765 = 9'h1e5 == _GEN_10152 ? phv_data_485 : _GEN_2764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2766 = 9'h1e6 == _GEN_10152 ? phv_data_486 : _GEN_2765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2767 = 9'h1e7 == _GEN_10152 ? phv_data_487 : _GEN_2766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2768 = 9'h1e8 == _GEN_10152 ? phv_data_488 : _GEN_2767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2769 = 9'h1e9 == _GEN_10152 ? phv_data_489 : _GEN_2768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2770 = 9'h1ea == _GEN_10152 ? phv_data_490 : _GEN_2769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2771 = 9'h1eb == _GEN_10152 ? phv_data_491 : _GEN_2770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2772 = 9'h1ec == _GEN_10152 ? phv_data_492 : _GEN_2771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2773 = 9'h1ed == _GEN_10152 ? phv_data_493 : _GEN_2772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2774 = 9'h1ee == _GEN_10152 ? phv_data_494 : _GEN_2773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2775 = 9'h1ef == _GEN_10152 ? phv_data_495 : _GEN_2774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2776 = 9'h1f0 == _GEN_10152 ? phv_data_496 : _GEN_2775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2777 = 9'h1f1 == _GEN_10152 ? phv_data_497 : _GEN_2776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2778 = 9'h1f2 == _GEN_10152 ? phv_data_498 : _GEN_2777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2779 = 9'h1f3 == _GEN_10152 ? phv_data_499 : _GEN_2778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2780 = 9'h1f4 == _GEN_10152 ? phv_data_500 : _GEN_2779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2781 = 9'h1f5 == _GEN_10152 ? phv_data_501 : _GEN_2780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2782 = 9'h1f6 == _GEN_10152 ? phv_data_502 : _GEN_2781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2783 = 9'h1f7 == _GEN_10152 ? phv_data_503 : _GEN_2782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2784 = 9'h1f8 == _GEN_10152 ? phv_data_504 : _GEN_2783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2785 = 9'h1f9 == _GEN_10152 ? phv_data_505 : _GEN_2784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2786 = 9'h1fa == _GEN_10152 ? phv_data_506 : _GEN_2785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2787 = 9'h1fb == _GEN_10152 ? phv_data_507 : _GEN_2786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2788 = 9'h1fc == _GEN_10152 ? phv_data_508 : _GEN_2787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2789 = 9'h1fd == _GEN_10152 ? phv_data_509 : _GEN_2788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2790 = 9'h1fe == _GEN_10152 ? phv_data_510 : _GEN_2789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_3 = 9'h1ff == _GEN_10152 ? phv_data_511 : _GEN_2790; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_10 = ending_1 == 2'h0; // @[executor.scala 199:88]
  wire  mask_1_3 = 2'h0 >= offset_1[1:0] & (2'h0 < ending_1 | ending_1 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_5 = {total_offset_hi_1,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_2793 = 8'h1 == total_offset_5 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2794 = 8'h2 == total_offset_5 ? phv_data_2 : _GEN_2793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2795 = 8'h3 == total_offset_5 ? phv_data_3 : _GEN_2794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2796 = 8'h4 == total_offset_5 ? phv_data_4 : _GEN_2795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2797 = 8'h5 == total_offset_5 ? phv_data_5 : _GEN_2796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2798 = 8'h6 == total_offset_5 ? phv_data_6 : _GEN_2797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2799 = 8'h7 == total_offset_5 ? phv_data_7 : _GEN_2798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2800 = 8'h8 == total_offset_5 ? phv_data_8 : _GEN_2799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2801 = 8'h9 == total_offset_5 ? phv_data_9 : _GEN_2800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2802 = 8'ha == total_offset_5 ? phv_data_10 : _GEN_2801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2803 = 8'hb == total_offset_5 ? phv_data_11 : _GEN_2802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2804 = 8'hc == total_offset_5 ? phv_data_12 : _GEN_2803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2805 = 8'hd == total_offset_5 ? phv_data_13 : _GEN_2804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2806 = 8'he == total_offset_5 ? phv_data_14 : _GEN_2805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2807 = 8'hf == total_offset_5 ? phv_data_15 : _GEN_2806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2808 = 8'h10 == total_offset_5 ? phv_data_16 : _GEN_2807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2809 = 8'h11 == total_offset_5 ? phv_data_17 : _GEN_2808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2810 = 8'h12 == total_offset_5 ? phv_data_18 : _GEN_2809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2811 = 8'h13 == total_offset_5 ? phv_data_19 : _GEN_2810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2812 = 8'h14 == total_offset_5 ? phv_data_20 : _GEN_2811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2813 = 8'h15 == total_offset_5 ? phv_data_21 : _GEN_2812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2814 = 8'h16 == total_offset_5 ? phv_data_22 : _GEN_2813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2815 = 8'h17 == total_offset_5 ? phv_data_23 : _GEN_2814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2816 = 8'h18 == total_offset_5 ? phv_data_24 : _GEN_2815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2817 = 8'h19 == total_offset_5 ? phv_data_25 : _GEN_2816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2818 = 8'h1a == total_offset_5 ? phv_data_26 : _GEN_2817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2819 = 8'h1b == total_offset_5 ? phv_data_27 : _GEN_2818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2820 = 8'h1c == total_offset_5 ? phv_data_28 : _GEN_2819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2821 = 8'h1d == total_offset_5 ? phv_data_29 : _GEN_2820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2822 = 8'h1e == total_offset_5 ? phv_data_30 : _GEN_2821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2823 = 8'h1f == total_offset_5 ? phv_data_31 : _GEN_2822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2824 = 8'h20 == total_offset_5 ? phv_data_32 : _GEN_2823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2825 = 8'h21 == total_offset_5 ? phv_data_33 : _GEN_2824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2826 = 8'h22 == total_offset_5 ? phv_data_34 : _GEN_2825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2827 = 8'h23 == total_offset_5 ? phv_data_35 : _GEN_2826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2828 = 8'h24 == total_offset_5 ? phv_data_36 : _GEN_2827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2829 = 8'h25 == total_offset_5 ? phv_data_37 : _GEN_2828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2830 = 8'h26 == total_offset_5 ? phv_data_38 : _GEN_2829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2831 = 8'h27 == total_offset_5 ? phv_data_39 : _GEN_2830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2832 = 8'h28 == total_offset_5 ? phv_data_40 : _GEN_2831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2833 = 8'h29 == total_offset_5 ? phv_data_41 : _GEN_2832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2834 = 8'h2a == total_offset_5 ? phv_data_42 : _GEN_2833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2835 = 8'h2b == total_offset_5 ? phv_data_43 : _GEN_2834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2836 = 8'h2c == total_offset_5 ? phv_data_44 : _GEN_2835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2837 = 8'h2d == total_offset_5 ? phv_data_45 : _GEN_2836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2838 = 8'h2e == total_offset_5 ? phv_data_46 : _GEN_2837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2839 = 8'h2f == total_offset_5 ? phv_data_47 : _GEN_2838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2840 = 8'h30 == total_offset_5 ? phv_data_48 : _GEN_2839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2841 = 8'h31 == total_offset_5 ? phv_data_49 : _GEN_2840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2842 = 8'h32 == total_offset_5 ? phv_data_50 : _GEN_2841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2843 = 8'h33 == total_offset_5 ? phv_data_51 : _GEN_2842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2844 = 8'h34 == total_offset_5 ? phv_data_52 : _GEN_2843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2845 = 8'h35 == total_offset_5 ? phv_data_53 : _GEN_2844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2846 = 8'h36 == total_offset_5 ? phv_data_54 : _GEN_2845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2847 = 8'h37 == total_offset_5 ? phv_data_55 : _GEN_2846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2848 = 8'h38 == total_offset_5 ? phv_data_56 : _GEN_2847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2849 = 8'h39 == total_offset_5 ? phv_data_57 : _GEN_2848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2850 = 8'h3a == total_offset_5 ? phv_data_58 : _GEN_2849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2851 = 8'h3b == total_offset_5 ? phv_data_59 : _GEN_2850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2852 = 8'h3c == total_offset_5 ? phv_data_60 : _GEN_2851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2853 = 8'h3d == total_offset_5 ? phv_data_61 : _GEN_2852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2854 = 8'h3e == total_offset_5 ? phv_data_62 : _GEN_2853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2855 = 8'h3f == total_offset_5 ? phv_data_63 : _GEN_2854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2856 = 8'h40 == total_offset_5 ? phv_data_64 : _GEN_2855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2857 = 8'h41 == total_offset_5 ? phv_data_65 : _GEN_2856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2858 = 8'h42 == total_offset_5 ? phv_data_66 : _GEN_2857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2859 = 8'h43 == total_offset_5 ? phv_data_67 : _GEN_2858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2860 = 8'h44 == total_offset_5 ? phv_data_68 : _GEN_2859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2861 = 8'h45 == total_offset_5 ? phv_data_69 : _GEN_2860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2862 = 8'h46 == total_offset_5 ? phv_data_70 : _GEN_2861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2863 = 8'h47 == total_offset_5 ? phv_data_71 : _GEN_2862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2864 = 8'h48 == total_offset_5 ? phv_data_72 : _GEN_2863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2865 = 8'h49 == total_offset_5 ? phv_data_73 : _GEN_2864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2866 = 8'h4a == total_offset_5 ? phv_data_74 : _GEN_2865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2867 = 8'h4b == total_offset_5 ? phv_data_75 : _GEN_2866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2868 = 8'h4c == total_offset_5 ? phv_data_76 : _GEN_2867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2869 = 8'h4d == total_offset_5 ? phv_data_77 : _GEN_2868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2870 = 8'h4e == total_offset_5 ? phv_data_78 : _GEN_2869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2871 = 8'h4f == total_offset_5 ? phv_data_79 : _GEN_2870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2872 = 8'h50 == total_offset_5 ? phv_data_80 : _GEN_2871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2873 = 8'h51 == total_offset_5 ? phv_data_81 : _GEN_2872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2874 = 8'h52 == total_offset_5 ? phv_data_82 : _GEN_2873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2875 = 8'h53 == total_offset_5 ? phv_data_83 : _GEN_2874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2876 = 8'h54 == total_offset_5 ? phv_data_84 : _GEN_2875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2877 = 8'h55 == total_offset_5 ? phv_data_85 : _GEN_2876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2878 = 8'h56 == total_offset_5 ? phv_data_86 : _GEN_2877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2879 = 8'h57 == total_offset_5 ? phv_data_87 : _GEN_2878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2880 = 8'h58 == total_offset_5 ? phv_data_88 : _GEN_2879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2881 = 8'h59 == total_offset_5 ? phv_data_89 : _GEN_2880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2882 = 8'h5a == total_offset_5 ? phv_data_90 : _GEN_2881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2883 = 8'h5b == total_offset_5 ? phv_data_91 : _GEN_2882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2884 = 8'h5c == total_offset_5 ? phv_data_92 : _GEN_2883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2885 = 8'h5d == total_offset_5 ? phv_data_93 : _GEN_2884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2886 = 8'h5e == total_offset_5 ? phv_data_94 : _GEN_2885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2887 = 8'h5f == total_offset_5 ? phv_data_95 : _GEN_2886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2888 = 8'h60 == total_offset_5 ? phv_data_96 : _GEN_2887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2889 = 8'h61 == total_offset_5 ? phv_data_97 : _GEN_2888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2890 = 8'h62 == total_offset_5 ? phv_data_98 : _GEN_2889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2891 = 8'h63 == total_offset_5 ? phv_data_99 : _GEN_2890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2892 = 8'h64 == total_offset_5 ? phv_data_100 : _GEN_2891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2893 = 8'h65 == total_offset_5 ? phv_data_101 : _GEN_2892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2894 = 8'h66 == total_offset_5 ? phv_data_102 : _GEN_2893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2895 = 8'h67 == total_offset_5 ? phv_data_103 : _GEN_2894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2896 = 8'h68 == total_offset_5 ? phv_data_104 : _GEN_2895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2897 = 8'h69 == total_offset_5 ? phv_data_105 : _GEN_2896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2898 = 8'h6a == total_offset_5 ? phv_data_106 : _GEN_2897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2899 = 8'h6b == total_offset_5 ? phv_data_107 : _GEN_2898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2900 = 8'h6c == total_offset_5 ? phv_data_108 : _GEN_2899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2901 = 8'h6d == total_offset_5 ? phv_data_109 : _GEN_2900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2902 = 8'h6e == total_offset_5 ? phv_data_110 : _GEN_2901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2903 = 8'h6f == total_offset_5 ? phv_data_111 : _GEN_2902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2904 = 8'h70 == total_offset_5 ? phv_data_112 : _GEN_2903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2905 = 8'h71 == total_offset_5 ? phv_data_113 : _GEN_2904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2906 = 8'h72 == total_offset_5 ? phv_data_114 : _GEN_2905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2907 = 8'h73 == total_offset_5 ? phv_data_115 : _GEN_2906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2908 = 8'h74 == total_offset_5 ? phv_data_116 : _GEN_2907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2909 = 8'h75 == total_offset_5 ? phv_data_117 : _GEN_2908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2910 = 8'h76 == total_offset_5 ? phv_data_118 : _GEN_2909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2911 = 8'h77 == total_offset_5 ? phv_data_119 : _GEN_2910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2912 = 8'h78 == total_offset_5 ? phv_data_120 : _GEN_2911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2913 = 8'h79 == total_offset_5 ? phv_data_121 : _GEN_2912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2914 = 8'h7a == total_offset_5 ? phv_data_122 : _GEN_2913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2915 = 8'h7b == total_offset_5 ? phv_data_123 : _GEN_2914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2916 = 8'h7c == total_offset_5 ? phv_data_124 : _GEN_2915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2917 = 8'h7d == total_offset_5 ? phv_data_125 : _GEN_2916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2918 = 8'h7e == total_offset_5 ? phv_data_126 : _GEN_2917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2919 = 8'h7f == total_offset_5 ? phv_data_127 : _GEN_2918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2920 = 8'h80 == total_offset_5 ? phv_data_128 : _GEN_2919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2921 = 8'h81 == total_offset_5 ? phv_data_129 : _GEN_2920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2922 = 8'h82 == total_offset_5 ? phv_data_130 : _GEN_2921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2923 = 8'h83 == total_offset_5 ? phv_data_131 : _GEN_2922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2924 = 8'h84 == total_offset_5 ? phv_data_132 : _GEN_2923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2925 = 8'h85 == total_offset_5 ? phv_data_133 : _GEN_2924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2926 = 8'h86 == total_offset_5 ? phv_data_134 : _GEN_2925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2927 = 8'h87 == total_offset_5 ? phv_data_135 : _GEN_2926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2928 = 8'h88 == total_offset_5 ? phv_data_136 : _GEN_2927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2929 = 8'h89 == total_offset_5 ? phv_data_137 : _GEN_2928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2930 = 8'h8a == total_offset_5 ? phv_data_138 : _GEN_2929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2931 = 8'h8b == total_offset_5 ? phv_data_139 : _GEN_2930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2932 = 8'h8c == total_offset_5 ? phv_data_140 : _GEN_2931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2933 = 8'h8d == total_offset_5 ? phv_data_141 : _GEN_2932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2934 = 8'h8e == total_offset_5 ? phv_data_142 : _GEN_2933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2935 = 8'h8f == total_offset_5 ? phv_data_143 : _GEN_2934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2936 = 8'h90 == total_offset_5 ? phv_data_144 : _GEN_2935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2937 = 8'h91 == total_offset_5 ? phv_data_145 : _GEN_2936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2938 = 8'h92 == total_offset_5 ? phv_data_146 : _GEN_2937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2939 = 8'h93 == total_offset_5 ? phv_data_147 : _GEN_2938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2940 = 8'h94 == total_offset_5 ? phv_data_148 : _GEN_2939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2941 = 8'h95 == total_offset_5 ? phv_data_149 : _GEN_2940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2942 = 8'h96 == total_offset_5 ? phv_data_150 : _GEN_2941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2943 = 8'h97 == total_offset_5 ? phv_data_151 : _GEN_2942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2944 = 8'h98 == total_offset_5 ? phv_data_152 : _GEN_2943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2945 = 8'h99 == total_offset_5 ? phv_data_153 : _GEN_2944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2946 = 8'h9a == total_offset_5 ? phv_data_154 : _GEN_2945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2947 = 8'h9b == total_offset_5 ? phv_data_155 : _GEN_2946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2948 = 8'h9c == total_offset_5 ? phv_data_156 : _GEN_2947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2949 = 8'h9d == total_offset_5 ? phv_data_157 : _GEN_2948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2950 = 8'h9e == total_offset_5 ? phv_data_158 : _GEN_2949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2951 = 8'h9f == total_offset_5 ? phv_data_159 : _GEN_2950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2952 = 8'ha0 == total_offset_5 ? phv_data_160 : _GEN_2951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2953 = 8'ha1 == total_offset_5 ? phv_data_161 : _GEN_2952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2954 = 8'ha2 == total_offset_5 ? phv_data_162 : _GEN_2953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2955 = 8'ha3 == total_offset_5 ? phv_data_163 : _GEN_2954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2956 = 8'ha4 == total_offset_5 ? phv_data_164 : _GEN_2955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2957 = 8'ha5 == total_offset_5 ? phv_data_165 : _GEN_2956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2958 = 8'ha6 == total_offset_5 ? phv_data_166 : _GEN_2957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2959 = 8'ha7 == total_offset_5 ? phv_data_167 : _GEN_2958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2960 = 8'ha8 == total_offset_5 ? phv_data_168 : _GEN_2959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2961 = 8'ha9 == total_offset_5 ? phv_data_169 : _GEN_2960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2962 = 8'haa == total_offset_5 ? phv_data_170 : _GEN_2961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2963 = 8'hab == total_offset_5 ? phv_data_171 : _GEN_2962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2964 = 8'hac == total_offset_5 ? phv_data_172 : _GEN_2963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2965 = 8'had == total_offset_5 ? phv_data_173 : _GEN_2964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2966 = 8'hae == total_offset_5 ? phv_data_174 : _GEN_2965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2967 = 8'haf == total_offset_5 ? phv_data_175 : _GEN_2966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2968 = 8'hb0 == total_offset_5 ? phv_data_176 : _GEN_2967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2969 = 8'hb1 == total_offset_5 ? phv_data_177 : _GEN_2968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2970 = 8'hb2 == total_offset_5 ? phv_data_178 : _GEN_2969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2971 = 8'hb3 == total_offset_5 ? phv_data_179 : _GEN_2970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2972 = 8'hb4 == total_offset_5 ? phv_data_180 : _GEN_2971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2973 = 8'hb5 == total_offset_5 ? phv_data_181 : _GEN_2972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2974 = 8'hb6 == total_offset_5 ? phv_data_182 : _GEN_2973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2975 = 8'hb7 == total_offset_5 ? phv_data_183 : _GEN_2974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2976 = 8'hb8 == total_offset_5 ? phv_data_184 : _GEN_2975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2977 = 8'hb9 == total_offset_5 ? phv_data_185 : _GEN_2976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2978 = 8'hba == total_offset_5 ? phv_data_186 : _GEN_2977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2979 = 8'hbb == total_offset_5 ? phv_data_187 : _GEN_2978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2980 = 8'hbc == total_offset_5 ? phv_data_188 : _GEN_2979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2981 = 8'hbd == total_offset_5 ? phv_data_189 : _GEN_2980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2982 = 8'hbe == total_offset_5 ? phv_data_190 : _GEN_2981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2983 = 8'hbf == total_offset_5 ? phv_data_191 : _GEN_2982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2984 = 8'hc0 == total_offset_5 ? phv_data_192 : _GEN_2983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2985 = 8'hc1 == total_offset_5 ? phv_data_193 : _GEN_2984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2986 = 8'hc2 == total_offset_5 ? phv_data_194 : _GEN_2985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2987 = 8'hc3 == total_offset_5 ? phv_data_195 : _GEN_2986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2988 = 8'hc4 == total_offset_5 ? phv_data_196 : _GEN_2987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2989 = 8'hc5 == total_offset_5 ? phv_data_197 : _GEN_2988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2990 = 8'hc6 == total_offset_5 ? phv_data_198 : _GEN_2989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2991 = 8'hc7 == total_offset_5 ? phv_data_199 : _GEN_2990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2992 = 8'hc8 == total_offset_5 ? phv_data_200 : _GEN_2991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2993 = 8'hc9 == total_offset_5 ? phv_data_201 : _GEN_2992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2994 = 8'hca == total_offset_5 ? phv_data_202 : _GEN_2993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2995 = 8'hcb == total_offset_5 ? phv_data_203 : _GEN_2994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2996 = 8'hcc == total_offset_5 ? phv_data_204 : _GEN_2995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2997 = 8'hcd == total_offset_5 ? phv_data_205 : _GEN_2996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2998 = 8'hce == total_offset_5 ? phv_data_206 : _GEN_2997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_2999 = 8'hcf == total_offset_5 ? phv_data_207 : _GEN_2998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3000 = 8'hd0 == total_offset_5 ? phv_data_208 : _GEN_2999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3001 = 8'hd1 == total_offset_5 ? phv_data_209 : _GEN_3000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3002 = 8'hd2 == total_offset_5 ? phv_data_210 : _GEN_3001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3003 = 8'hd3 == total_offset_5 ? phv_data_211 : _GEN_3002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3004 = 8'hd4 == total_offset_5 ? phv_data_212 : _GEN_3003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3005 = 8'hd5 == total_offset_5 ? phv_data_213 : _GEN_3004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3006 = 8'hd6 == total_offset_5 ? phv_data_214 : _GEN_3005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3007 = 8'hd7 == total_offset_5 ? phv_data_215 : _GEN_3006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3008 = 8'hd8 == total_offset_5 ? phv_data_216 : _GEN_3007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3009 = 8'hd9 == total_offset_5 ? phv_data_217 : _GEN_3008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3010 = 8'hda == total_offset_5 ? phv_data_218 : _GEN_3009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3011 = 8'hdb == total_offset_5 ? phv_data_219 : _GEN_3010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3012 = 8'hdc == total_offset_5 ? phv_data_220 : _GEN_3011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3013 = 8'hdd == total_offset_5 ? phv_data_221 : _GEN_3012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3014 = 8'hde == total_offset_5 ? phv_data_222 : _GEN_3013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3015 = 8'hdf == total_offset_5 ? phv_data_223 : _GEN_3014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3016 = 8'he0 == total_offset_5 ? phv_data_224 : _GEN_3015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3017 = 8'he1 == total_offset_5 ? phv_data_225 : _GEN_3016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3018 = 8'he2 == total_offset_5 ? phv_data_226 : _GEN_3017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3019 = 8'he3 == total_offset_5 ? phv_data_227 : _GEN_3018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3020 = 8'he4 == total_offset_5 ? phv_data_228 : _GEN_3019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3021 = 8'he5 == total_offset_5 ? phv_data_229 : _GEN_3020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3022 = 8'he6 == total_offset_5 ? phv_data_230 : _GEN_3021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3023 = 8'he7 == total_offset_5 ? phv_data_231 : _GEN_3022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3024 = 8'he8 == total_offset_5 ? phv_data_232 : _GEN_3023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3025 = 8'he9 == total_offset_5 ? phv_data_233 : _GEN_3024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3026 = 8'hea == total_offset_5 ? phv_data_234 : _GEN_3025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3027 = 8'heb == total_offset_5 ? phv_data_235 : _GEN_3026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3028 = 8'hec == total_offset_5 ? phv_data_236 : _GEN_3027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3029 = 8'hed == total_offset_5 ? phv_data_237 : _GEN_3028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3030 = 8'hee == total_offset_5 ? phv_data_238 : _GEN_3029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3031 = 8'hef == total_offset_5 ? phv_data_239 : _GEN_3030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3032 = 8'hf0 == total_offset_5 ? phv_data_240 : _GEN_3031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3033 = 8'hf1 == total_offset_5 ? phv_data_241 : _GEN_3032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3034 = 8'hf2 == total_offset_5 ? phv_data_242 : _GEN_3033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3035 = 8'hf3 == total_offset_5 ? phv_data_243 : _GEN_3034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3036 = 8'hf4 == total_offset_5 ? phv_data_244 : _GEN_3035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3037 = 8'hf5 == total_offset_5 ? phv_data_245 : _GEN_3036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3038 = 8'hf6 == total_offset_5 ? phv_data_246 : _GEN_3037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3039 = 8'hf7 == total_offset_5 ? phv_data_247 : _GEN_3038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3040 = 8'hf8 == total_offset_5 ? phv_data_248 : _GEN_3039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3041 = 8'hf9 == total_offset_5 ? phv_data_249 : _GEN_3040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3042 = 8'hfa == total_offset_5 ? phv_data_250 : _GEN_3041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3043 = 8'hfb == total_offset_5 ? phv_data_251 : _GEN_3042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3044 = 8'hfc == total_offset_5 ? phv_data_252 : _GEN_3043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3045 = 8'hfd == total_offset_5 ? phv_data_253 : _GEN_3044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3046 = 8'hfe == total_offset_5 ? phv_data_254 : _GEN_3045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3047 = 8'hff == total_offset_5 ? phv_data_255 : _GEN_3046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_10408 = {{1'd0}, total_offset_5}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3048 = 9'h100 == _GEN_10408 ? phv_data_256 : _GEN_3047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3049 = 9'h101 == _GEN_10408 ? phv_data_257 : _GEN_3048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3050 = 9'h102 == _GEN_10408 ? phv_data_258 : _GEN_3049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3051 = 9'h103 == _GEN_10408 ? phv_data_259 : _GEN_3050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3052 = 9'h104 == _GEN_10408 ? phv_data_260 : _GEN_3051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3053 = 9'h105 == _GEN_10408 ? phv_data_261 : _GEN_3052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3054 = 9'h106 == _GEN_10408 ? phv_data_262 : _GEN_3053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3055 = 9'h107 == _GEN_10408 ? phv_data_263 : _GEN_3054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3056 = 9'h108 == _GEN_10408 ? phv_data_264 : _GEN_3055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3057 = 9'h109 == _GEN_10408 ? phv_data_265 : _GEN_3056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3058 = 9'h10a == _GEN_10408 ? phv_data_266 : _GEN_3057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3059 = 9'h10b == _GEN_10408 ? phv_data_267 : _GEN_3058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3060 = 9'h10c == _GEN_10408 ? phv_data_268 : _GEN_3059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3061 = 9'h10d == _GEN_10408 ? phv_data_269 : _GEN_3060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3062 = 9'h10e == _GEN_10408 ? phv_data_270 : _GEN_3061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3063 = 9'h10f == _GEN_10408 ? phv_data_271 : _GEN_3062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3064 = 9'h110 == _GEN_10408 ? phv_data_272 : _GEN_3063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3065 = 9'h111 == _GEN_10408 ? phv_data_273 : _GEN_3064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3066 = 9'h112 == _GEN_10408 ? phv_data_274 : _GEN_3065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3067 = 9'h113 == _GEN_10408 ? phv_data_275 : _GEN_3066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3068 = 9'h114 == _GEN_10408 ? phv_data_276 : _GEN_3067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3069 = 9'h115 == _GEN_10408 ? phv_data_277 : _GEN_3068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3070 = 9'h116 == _GEN_10408 ? phv_data_278 : _GEN_3069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3071 = 9'h117 == _GEN_10408 ? phv_data_279 : _GEN_3070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3072 = 9'h118 == _GEN_10408 ? phv_data_280 : _GEN_3071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3073 = 9'h119 == _GEN_10408 ? phv_data_281 : _GEN_3072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3074 = 9'h11a == _GEN_10408 ? phv_data_282 : _GEN_3073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3075 = 9'h11b == _GEN_10408 ? phv_data_283 : _GEN_3074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3076 = 9'h11c == _GEN_10408 ? phv_data_284 : _GEN_3075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3077 = 9'h11d == _GEN_10408 ? phv_data_285 : _GEN_3076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3078 = 9'h11e == _GEN_10408 ? phv_data_286 : _GEN_3077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3079 = 9'h11f == _GEN_10408 ? phv_data_287 : _GEN_3078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3080 = 9'h120 == _GEN_10408 ? phv_data_288 : _GEN_3079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3081 = 9'h121 == _GEN_10408 ? phv_data_289 : _GEN_3080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3082 = 9'h122 == _GEN_10408 ? phv_data_290 : _GEN_3081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3083 = 9'h123 == _GEN_10408 ? phv_data_291 : _GEN_3082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3084 = 9'h124 == _GEN_10408 ? phv_data_292 : _GEN_3083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3085 = 9'h125 == _GEN_10408 ? phv_data_293 : _GEN_3084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3086 = 9'h126 == _GEN_10408 ? phv_data_294 : _GEN_3085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3087 = 9'h127 == _GEN_10408 ? phv_data_295 : _GEN_3086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3088 = 9'h128 == _GEN_10408 ? phv_data_296 : _GEN_3087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3089 = 9'h129 == _GEN_10408 ? phv_data_297 : _GEN_3088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3090 = 9'h12a == _GEN_10408 ? phv_data_298 : _GEN_3089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3091 = 9'h12b == _GEN_10408 ? phv_data_299 : _GEN_3090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3092 = 9'h12c == _GEN_10408 ? phv_data_300 : _GEN_3091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3093 = 9'h12d == _GEN_10408 ? phv_data_301 : _GEN_3092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3094 = 9'h12e == _GEN_10408 ? phv_data_302 : _GEN_3093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3095 = 9'h12f == _GEN_10408 ? phv_data_303 : _GEN_3094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3096 = 9'h130 == _GEN_10408 ? phv_data_304 : _GEN_3095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3097 = 9'h131 == _GEN_10408 ? phv_data_305 : _GEN_3096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3098 = 9'h132 == _GEN_10408 ? phv_data_306 : _GEN_3097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3099 = 9'h133 == _GEN_10408 ? phv_data_307 : _GEN_3098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3100 = 9'h134 == _GEN_10408 ? phv_data_308 : _GEN_3099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3101 = 9'h135 == _GEN_10408 ? phv_data_309 : _GEN_3100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3102 = 9'h136 == _GEN_10408 ? phv_data_310 : _GEN_3101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3103 = 9'h137 == _GEN_10408 ? phv_data_311 : _GEN_3102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3104 = 9'h138 == _GEN_10408 ? phv_data_312 : _GEN_3103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3105 = 9'h139 == _GEN_10408 ? phv_data_313 : _GEN_3104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3106 = 9'h13a == _GEN_10408 ? phv_data_314 : _GEN_3105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3107 = 9'h13b == _GEN_10408 ? phv_data_315 : _GEN_3106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3108 = 9'h13c == _GEN_10408 ? phv_data_316 : _GEN_3107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3109 = 9'h13d == _GEN_10408 ? phv_data_317 : _GEN_3108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3110 = 9'h13e == _GEN_10408 ? phv_data_318 : _GEN_3109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3111 = 9'h13f == _GEN_10408 ? phv_data_319 : _GEN_3110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3112 = 9'h140 == _GEN_10408 ? phv_data_320 : _GEN_3111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3113 = 9'h141 == _GEN_10408 ? phv_data_321 : _GEN_3112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3114 = 9'h142 == _GEN_10408 ? phv_data_322 : _GEN_3113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3115 = 9'h143 == _GEN_10408 ? phv_data_323 : _GEN_3114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3116 = 9'h144 == _GEN_10408 ? phv_data_324 : _GEN_3115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3117 = 9'h145 == _GEN_10408 ? phv_data_325 : _GEN_3116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3118 = 9'h146 == _GEN_10408 ? phv_data_326 : _GEN_3117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3119 = 9'h147 == _GEN_10408 ? phv_data_327 : _GEN_3118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3120 = 9'h148 == _GEN_10408 ? phv_data_328 : _GEN_3119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3121 = 9'h149 == _GEN_10408 ? phv_data_329 : _GEN_3120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3122 = 9'h14a == _GEN_10408 ? phv_data_330 : _GEN_3121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3123 = 9'h14b == _GEN_10408 ? phv_data_331 : _GEN_3122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3124 = 9'h14c == _GEN_10408 ? phv_data_332 : _GEN_3123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3125 = 9'h14d == _GEN_10408 ? phv_data_333 : _GEN_3124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3126 = 9'h14e == _GEN_10408 ? phv_data_334 : _GEN_3125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3127 = 9'h14f == _GEN_10408 ? phv_data_335 : _GEN_3126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3128 = 9'h150 == _GEN_10408 ? phv_data_336 : _GEN_3127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3129 = 9'h151 == _GEN_10408 ? phv_data_337 : _GEN_3128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3130 = 9'h152 == _GEN_10408 ? phv_data_338 : _GEN_3129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3131 = 9'h153 == _GEN_10408 ? phv_data_339 : _GEN_3130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3132 = 9'h154 == _GEN_10408 ? phv_data_340 : _GEN_3131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3133 = 9'h155 == _GEN_10408 ? phv_data_341 : _GEN_3132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3134 = 9'h156 == _GEN_10408 ? phv_data_342 : _GEN_3133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3135 = 9'h157 == _GEN_10408 ? phv_data_343 : _GEN_3134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3136 = 9'h158 == _GEN_10408 ? phv_data_344 : _GEN_3135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3137 = 9'h159 == _GEN_10408 ? phv_data_345 : _GEN_3136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3138 = 9'h15a == _GEN_10408 ? phv_data_346 : _GEN_3137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3139 = 9'h15b == _GEN_10408 ? phv_data_347 : _GEN_3138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3140 = 9'h15c == _GEN_10408 ? phv_data_348 : _GEN_3139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3141 = 9'h15d == _GEN_10408 ? phv_data_349 : _GEN_3140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3142 = 9'h15e == _GEN_10408 ? phv_data_350 : _GEN_3141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3143 = 9'h15f == _GEN_10408 ? phv_data_351 : _GEN_3142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3144 = 9'h160 == _GEN_10408 ? phv_data_352 : _GEN_3143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3145 = 9'h161 == _GEN_10408 ? phv_data_353 : _GEN_3144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3146 = 9'h162 == _GEN_10408 ? phv_data_354 : _GEN_3145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3147 = 9'h163 == _GEN_10408 ? phv_data_355 : _GEN_3146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3148 = 9'h164 == _GEN_10408 ? phv_data_356 : _GEN_3147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3149 = 9'h165 == _GEN_10408 ? phv_data_357 : _GEN_3148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3150 = 9'h166 == _GEN_10408 ? phv_data_358 : _GEN_3149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3151 = 9'h167 == _GEN_10408 ? phv_data_359 : _GEN_3150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3152 = 9'h168 == _GEN_10408 ? phv_data_360 : _GEN_3151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3153 = 9'h169 == _GEN_10408 ? phv_data_361 : _GEN_3152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3154 = 9'h16a == _GEN_10408 ? phv_data_362 : _GEN_3153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3155 = 9'h16b == _GEN_10408 ? phv_data_363 : _GEN_3154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3156 = 9'h16c == _GEN_10408 ? phv_data_364 : _GEN_3155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3157 = 9'h16d == _GEN_10408 ? phv_data_365 : _GEN_3156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3158 = 9'h16e == _GEN_10408 ? phv_data_366 : _GEN_3157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3159 = 9'h16f == _GEN_10408 ? phv_data_367 : _GEN_3158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3160 = 9'h170 == _GEN_10408 ? phv_data_368 : _GEN_3159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3161 = 9'h171 == _GEN_10408 ? phv_data_369 : _GEN_3160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3162 = 9'h172 == _GEN_10408 ? phv_data_370 : _GEN_3161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3163 = 9'h173 == _GEN_10408 ? phv_data_371 : _GEN_3162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3164 = 9'h174 == _GEN_10408 ? phv_data_372 : _GEN_3163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3165 = 9'h175 == _GEN_10408 ? phv_data_373 : _GEN_3164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3166 = 9'h176 == _GEN_10408 ? phv_data_374 : _GEN_3165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3167 = 9'h177 == _GEN_10408 ? phv_data_375 : _GEN_3166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3168 = 9'h178 == _GEN_10408 ? phv_data_376 : _GEN_3167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3169 = 9'h179 == _GEN_10408 ? phv_data_377 : _GEN_3168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3170 = 9'h17a == _GEN_10408 ? phv_data_378 : _GEN_3169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3171 = 9'h17b == _GEN_10408 ? phv_data_379 : _GEN_3170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3172 = 9'h17c == _GEN_10408 ? phv_data_380 : _GEN_3171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3173 = 9'h17d == _GEN_10408 ? phv_data_381 : _GEN_3172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3174 = 9'h17e == _GEN_10408 ? phv_data_382 : _GEN_3173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3175 = 9'h17f == _GEN_10408 ? phv_data_383 : _GEN_3174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3176 = 9'h180 == _GEN_10408 ? phv_data_384 : _GEN_3175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3177 = 9'h181 == _GEN_10408 ? phv_data_385 : _GEN_3176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3178 = 9'h182 == _GEN_10408 ? phv_data_386 : _GEN_3177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3179 = 9'h183 == _GEN_10408 ? phv_data_387 : _GEN_3178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3180 = 9'h184 == _GEN_10408 ? phv_data_388 : _GEN_3179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3181 = 9'h185 == _GEN_10408 ? phv_data_389 : _GEN_3180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3182 = 9'h186 == _GEN_10408 ? phv_data_390 : _GEN_3181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3183 = 9'h187 == _GEN_10408 ? phv_data_391 : _GEN_3182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3184 = 9'h188 == _GEN_10408 ? phv_data_392 : _GEN_3183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3185 = 9'h189 == _GEN_10408 ? phv_data_393 : _GEN_3184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3186 = 9'h18a == _GEN_10408 ? phv_data_394 : _GEN_3185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3187 = 9'h18b == _GEN_10408 ? phv_data_395 : _GEN_3186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3188 = 9'h18c == _GEN_10408 ? phv_data_396 : _GEN_3187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3189 = 9'h18d == _GEN_10408 ? phv_data_397 : _GEN_3188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3190 = 9'h18e == _GEN_10408 ? phv_data_398 : _GEN_3189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3191 = 9'h18f == _GEN_10408 ? phv_data_399 : _GEN_3190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3192 = 9'h190 == _GEN_10408 ? phv_data_400 : _GEN_3191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3193 = 9'h191 == _GEN_10408 ? phv_data_401 : _GEN_3192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3194 = 9'h192 == _GEN_10408 ? phv_data_402 : _GEN_3193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3195 = 9'h193 == _GEN_10408 ? phv_data_403 : _GEN_3194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3196 = 9'h194 == _GEN_10408 ? phv_data_404 : _GEN_3195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3197 = 9'h195 == _GEN_10408 ? phv_data_405 : _GEN_3196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3198 = 9'h196 == _GEN_10408 ? phv_data_406 : _GEN_3197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3199 = 9'h197 == _GEN_10408 ? phv_data_407 : _GEN_3198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3200 = 9'h198 == _GEN_10408 ? phv_data_408 : _GEN_3199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3201 = 9'h199 == _GEN_10408 ? phv_data_409 : _GEN_3200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3202 = 9'h19a == _GEN_10408 ? phv_data_410 : _GEN_3201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3203 = 9'h19b == _GEN_10408 ? phv_data_411 : _GEN_3202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3204 = 9'h19c == _GEN_10408 ? phv_data_412 : _GEN_3203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3205 = 9'h19d == _GEN_10408 ? phv_data_413 : _GEN_3204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3206 = 9'h19e == _GEN_10408 ? phv_data_414 : _GEN_3205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3207 = 9'h19f == _GEN_10408 ? phv_data_415 : _GEN_3206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3208 = 9'h1a0 == _GEN_10408 ? phv_data_416 : _GEN_3207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3209 = 9'h1a1 == _GEN_10408 ? phv_data_417 : _GEN_3208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3210 = 9'h1a2 == _GEN_10408 ? phv_data_418 : _GEN_3209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3211 = 9'h1a3 == _GEN_10408 ? phv_data_419 : _GEN_3210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3212 = 9'h1a4 == _GEN_10408 ? phv_data_420 : _GEN_3211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3213 = 9'h1a5 == _GEN_10408 ? phv_data_421 : _GEN_3212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3214 = 9'h1a6 == _GEN_10408 ? phv_data_422 : _GEN_3213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3215 = 9'h1a7 == _GEN_10408 ? phv_data_423 : _GEN_3214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3216 = 9'h1a8 == _GEN_10408 ? phv_data_424 : _GEN_3215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3217 = 9'h1a9 == _GEN_10408 ? phv_data_425 : _GEN_3216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3218 = 9'h1aa == _GEN_10408 ? phv_data_426 : _GEN_3217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3219 = 9'h1ab == _GEN_10408 ? phv_data_427 : _GEN_3218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3220 = 9'h1ac == _GEN_10408 ? phv_data_428 : _GEN_3219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3221 = 9'h1ad == _GEN_10408 ? phv_data_429 : _GEN_3220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3222 = 9'h1ae == _GEN_10408 ? phv_data_430 : _GEN_3221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3223 = 9'h1af == _GEN_10408 ? phv_data_431 : _GEN_3222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3224 = 9'h1b0 == _GEN_10408 ? phv_data_432 : _GEN_3223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3225 = 9'h1b1 == _GEN_10408 ? phv_data_433 : _GEN_3224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3226 = 9'h1b2 == _GEN_10408 ? phv_data_434 : _GEN_3225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3227 = 9'h1b3 == _GEN_10408 ? phv_data_435 : _GEN_3226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3228 = 9'h1b4 == _GEN_10408 ? phv_data_436 : _GEN_3227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3229 = 9'h1b5 == _GEN_10408 ? phv_data_437 : _GEN_3228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3230 = 9'h1b6 == _GEN_10408 ? phv_data_438 : _GEN_3229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3231 = 9'h1b7 == _GEN_10408 ? phv_data_439 : _GEN_3230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3232 = 9'h1b8 == _GEN_10408 ? phv_data_440 : _GEN_3231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3233 = 9'h1b9 == _GEN_10408 ? phv_data_441 : _GEN_3232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3234 = 9'h1ba == _GEN_10408 ? phv_data_442 : _GEN_3233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3235 = 9'h1bb == _GEN_10408 ? phv_data_443 : _GEN_3234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3236 = 9'h1bc == _GEN_10408 ? phv_data_444 : _GEN_3235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3237 = 9'h1bd == _GEN_10408 ? phv_data_445 : _GEN_3236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3238 = 9'h1be == _GEN_10408 ? phv_data_446 : _GEN_3237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3239 = 9'h1bf == _GEN_10408 ? phv_data_447 : _GEN_3238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3240 = 9'h1c0 == _GEN_10408 ? phv_data_448 : _GEN_3239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3241 = 9'h1c1 == _GEN_10408 ? phv_data_449 : _GEN_3240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3242 = 9'h1c2 == _GEN_10408 ? phv_data_450 : _GEN_3241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3243 = 9'h1c3 == _GEN_10408 ? phv_data_451 : _GEN_3242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3244 = 9'h1c4 == _GEN_10408 ? phv_data_452 : _GEN_3243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3245 = 9'h1c5 == _GEN_10408 ? phv_data_453 : _GEN_3244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3246 = 9'h1c6 == _GEN_10408 ? phv_data_454 : _GEN_3245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3247 = 9'h1c7 == _GEN_10408 ? phv_data_455 : _GEN_3246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3248 = 9'h1c8 == _GEN_10408 ? phv_data_456 : _GEN_3247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3249 = 9'h1c9 == _GEN_10408 ? phv_data_457 : _GEN_3248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3250 = 9'h1ca == _GEN_10408 ? phv_data_458 : _GEN_3249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3251 = 9'h1cb == _GEN_10408 ? phv_data_459 : _GEN_3250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3252 = 9'h1cc == _GEN_10408 ? phv_data_460 : _GEN_3251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3253 = 9'h1cd == _GEN_10408 ? phv_data_461 : _GEN_3252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3254 = 9'h1ce == _GEN_10408 ? phv_data_462 : _GEN_3253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3255 = 9'h1cf == _GEN_10408 ? phv_data_463 : _GEN_3254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3256 = 9'h1d0 == _GEN_10408 ? phv_data_464 : _GEN_3255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3257 = 9'h1d1 == _GEN_10408 ? phv_data_465 : _GEN_3256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3258 = 9'h1d2 == _GEN_10408 ? phv_data_466 : _GEN_3257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3259 = 9'h1d3 == _GEN_10408 ? phv_data_467 : _GEN_3258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3260 = 9'h1d4 == _GEN_10408 ? phv_data_468 : _GEN_3259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3261 = 9'h1d5 == _GEN_10408 ? phv_data_469 : _GEN_3260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3262 = 9'h1d6 == _GEN_10408 ? phv_data_470 : _GEN_3261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3263 = 9'h1d7 == _GEN_10408 ? phv_data_471 : _GEN_3262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3264 = 9'h1d8 == _GEN_10408 ? phv_data_472 : _GEN_3263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3265 = 9'h1d9 == _GEN_10408 ? phv_data_473 : _GEN_3264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3266 = 9'h1da == _GEN_10408 ? phv_data_474 : _GEN_3265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3267 = 9'h1db == _GEN_10408 ? phv_data_475 : _GEN_3266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3268 = 9'h1dc == _GEN_10408 ? phv_data_476 : _GEN_3267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3269 = 9'h1dd == _GEN_10408 ? phv_data_477 : _GEN_3268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3270 = 9'h1de == _GEN_10408 ? phv_data_478 : _GEN_3269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3271 = 9'h1df == _GEN_10408 ? phv_data_479 : _GEN_3270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3272 = 9'h1e0 == _GEN_10408 ? phv_data_480 : _GEN_3271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3273 = 9'h1e1 == _GEN_10408 ? phv_data_481 : _GEN_3272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3274 = 9'h1e2 == _GEN_10408 ? phv_data_482 : _GEN_3273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3275 = 9'h1e3 == _GEN_10408 ? phv_data_483 : _GEN_3274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3276 = 9'h1e4 == _GEN_10408 ? phv_data_484 : _GEN_3275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3277 = 9'h1e5 == _GEN_10408 ? phv_data_485 : _GEN_3276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3278 = 9'h1e6 == _GEN_10408 ? phv_data_486 : _GEN_3277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3279 = 9'h1e7 == _GEN_10408 ? phv_data_487 : _GEN_3278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3280 = 9'h1e8 == _GEN_10408 ? phv_data_488 : _GEN_3279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3281 = 9'h1e9 == _GEN_10408 ? phv_data_489 : _GEN_3280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3282 = 9'h1ea == _GEN_10408 ? phv_data_490 : _GEN_3281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3283 = 9'h1eb == _GEN_10408 ? phv_data_491 : _GEN_3282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3284 = 9'h1ec == _GEN_10408 ? phv_data_492 : _GEN_3283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3285 = 9'h1ed == _GEN_10408 ? phv_data_493 : _GEN_3284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3286 = 9'h1ee == _GEN_10408 ? phv_data_494 : _GEN_3285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3287 = 9'h1ef == _GEN_10408 ? phv_data_495 : _GEN_3286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3288 = 9'h1f0 == _GEN_10408 ? phv_data_496 : _GEN_3287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3289 = 9'h1f1 == _GEN_10408 ? phv_data_497 : _GEN_3288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3290 = 9'h1f2 == _GEN_10408 ? phv_data_498 : _GEN_3289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3291 = 9'h1f3 == _GEN_10408 ? phv_data_499 : _GEN_3290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3292 = 9'h1f4 == _GEN_10408 ? phv_data_500 : _GEN_3291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3293 = 9'h1f5 == _GEN_10408 ? phv_data_501 : _GEN_3292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3294 = 9'h1f6 == _GEN_10408 ? phv_data_502 : _GEN_3293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3295 = 9'h1f7 == _GEN_10408 ? phv_data_503 : _GEN_3294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3296 = 9'h1f8 == _GEN_10408 ? phv_data_504 : _GEN_3295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3297 = 9'h1f9 == _GEN_10408 ? phv_data_505 : _GEN_3296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3298 = 9'h1fa == _GEN_10408 ? phv_data_506 : _GEN_3297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3299 = 9'h1fb == _GEN_10408 ? phv_data_507 : _GEN_3298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3300 = 9'h1fc == _GEN_10408 ? phv_data_508 : _GEN_3299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3301 = 9'h1fd == _GEN_10408 ? phv_data_509 : _GEN_3300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3302 = 9'h1fe == _GEN_10408 ? phv_data_510 : _GEN_3301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_2 = 9'h1ff == _GEN_10408 ? phv_data_511 : _GEN_3302; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_1_2 = 2'h1 >= offset_1[1:0] & (2'h1 < ending_1 | ending_1 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_6 = {total_offset_hi_1,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_3305 = 8'h1 == total_offset_6 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3306 = 8'h2 == total_offset_6 ? phv_data_2 : _GEN_3305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3307 = 8'h3 == total_offset_6 ? phv_data_3 : _GEN_3306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3308 = 8'h4 == total_offset_6 ? phv_data_4 : _GEN_3307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3309 = 8'h5 == total_offset_6 ? phv_data_5 : _GEN_3308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3310 = 8'h6 == total_offset_6 ? phv_data_6 : _GEN_3309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3311 = 8'h7 == total_offset_6 ? phv_data_7 : _GEN_3310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3312 = 8'h8 == total_offset_6 ? phv_data_8 : _GEN_3311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3313 = 8'h9 == total_offset_6 ? phv_data_9 : _GEN_3312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3314 = 8'ha == total_offset_6 ? phv_data_10 : _GEN_3313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3315 = 8'hb == total_offset_6 ? phv_data_11 : _GEN_3314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3316 = 8'hc == total_offset_6 ? phv_data_12 : _GEN_3315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3317 = 8'hd == total_offset_6 ? phv_data_13 : _GEN_3316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3318 = 8'he == total_offset_6 ? phv_data_14 : _GEN_3317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3319 = 8'hf == total_offset_6 ? phv_data_15 : _GEN_3318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3320 = 8'h10 == total_offset_6 ? phv_data_16 : _GEN_3319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3321 = 8'h11 == total_offset_6 ? phv_data_17 : _GEN_3320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3322 = 8'h12 == total_offset_6 ? phv_data_18 : _GEN_3321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3323 = 8'h13 == total_offset_6 ? phv_data_19 : _GEN_3322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3324 = 8'h14 == total_offset_6 ? phv_data_20 : _GEN_3323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3325 = 8'h15 == total_offset_6 ? phv_data_21 : _GEN_3324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3326 = 8'h16 == total_offset_6 ? phv_data_22 : _GEN_3325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3327 = 8'h17 == total_offset_6 ? phv_data_23 : _GEN_3326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3328 = 8'h18 == total_offset_6 ? phv_data_24 : _GEN_3327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3329 = 8'h19 == total_offset_6 ? phv_data_25 : _GEN_3328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3330 = 8'h1a == total_offset_6 ? phv_data_26 : _GEN_3329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3331 = 8'h1b == total_offset_6 ? phv_data_27 : _GEN_3330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3332 = 8'h1c == total_offset_6 ? phv_data_28 : _GEN_3331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3333 = 8'h1d == total_offset_6 ? phv_data_29 : _GEN_3332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3334 = 8'h1e == total_offset_6 ? phv_data_30 : _GEN_3333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3335 = 8'h1f == total_offset_6 ? phv_data_31 : _GEN_3334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3336 = 8'h20 == total_offset_6 ? phv_data_32 : _GEN_3335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3337 = 8'h21 == total_offset_6 ? phv_data_33 : _GEN_3336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3338 = 8'h22 == total_offset_6 ? phv_data_34 : _GEN_3337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3339 = 8'h23 == total_offset_6 ? phv_data_35 : _GEN_3338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3340 = 8'h24 == total_offset_6 ? phv_data_36 : _GEN_3339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3341 = 8'h25 == total_offset_6 ? phv_data_37 : _GEN_3340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3342 = 8'h26 == total_offset_6 ? phv_data_38 : _GEN_3341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3343 = 8'h27 == total_offset_6 ? phv_data_39 : _GEN_3342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3344 = 8'h28 == total_offset_6 ? phv_data_40 : _GEN_3343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3345 = 8'h29 == total_offset_6 ? phv_data_41 : _GEN_3344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3346 = 8'h2a == total_offset_6 ? phv_data_42 : _GEN_3345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3347 = 8'h2b == total_offset_6 ? phv_data_43 : _GEN_3346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3348 = 8'h2c == total_offset_6 ? phv_data_44 : _GEN_3347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3349 = 8'h2d == total_offset_6 ? phv_data_45 : _GEN_3348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3350 = 8'h2e == total_offset_6 ? phv_data_46 : _GEN_3349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3351 = 8'h2f == total_offset_6 ? phv_data_47 : _GEN_3350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3352 = 8'h30 == total_offset_6 ? phv_data_48 : _GEN_3351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3353 = 8'h31 == total_offset_6 ? phv_data_49 : _GEN_3352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3354 = 8'h32 == total_offset_6 ? phv_data_50 : _GEN_3353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3355 = 8'h33 == total_offset_6 ? phv_data_51 : _GEN_3354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3356 = 8'h34 == total_offset_6 ? phv_data_52 : _GEN_3355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3357 = 8'h35 == total_offset_6 ? phv_data_53 : _GEN_3356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3358 = 8'h36 == total_offset_6 ? phv_data_54 : _GEN_3357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3359 = 8'h37 == total_offset_6 ? phv_data_55 : _GEN_3358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3360 = 8'h38 == total_offset_6 ? phv_data_56 : _GEN_3359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3361 = 8'h39 == total_offset_6 ? phv_data_57 : _GEN_3360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3362 = 8'h3a == total_offset_6 ? phv_data_58 : _GEN_3361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3363 = 8'h3b == total_offset_6 ? phv_data_59 : _GEN_3362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3364 = 8'h3c == total_offset_6 ? phv_data_60 : _GEN_3363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3365 = 8'h3d == total_offset_6 ? phv_data_61 : _GEN_3364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3366 = 8'h3e == total_offset_6 ? phv_data_62 : _GEN_3365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3367 = 8'h3f == total_offset_6 ? phv_data_63 : _GEN_3366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3368 = 8'h40 == total_offset_6 ? phv_data_64 : _GEN_3367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3369 = 8'h41 == total_offset_6 ? phv_data_65 : _GEN_3368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3370 = 8'h42 == total_offset_6 ? phv_data_66 : _GEN_3369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3371 = 8'h43 == total_offset_6 ? phv_data_67 : _GEN_3370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3372 = 8'h44 == total_offset_6 ? phv_data_68 : _GEN_3371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3373 = 8'h45 == total_offset_6 ? phv_data_69 : _GEN_3372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3374 = 8'h46 == total_offset_6 ? phv_data_70 : _GEN_3373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3375 = 8'h47 == total_offset_6 ? phv_data_71 : _GEN_3374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3376 = 8'h48 == total_offset_6 ? phv_data_72 : _GEN_3375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3377 = 8'h49 == total_offset_6 ? phv_data_73 : _GEN_3376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3378 = 8'h4a == total_offset_6 ? phv_data_74 : _GEN_3377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3379 = 8'h4b == total_offset_6 ? phv_data_75 : _GEN_3378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3380 = 8'h4c == total_offset_6 ? phv_data_76 : _GEN_3379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3381 = 8'h4d == total_offset_6 ? phv_data_77 : _GEN_3380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3382 = 8'h4e == total_offset_6 ? phv_data_78 : _GEN_3381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3383 = 8'h4f == total_offset_6 ? phv_data_79 : _GEN_3382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3384 = 8'h50 == total_offset_6 ? phv_data_80 : _GEN_3383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3385 = 8'h51 == total_offset_6 ? phv_data_81 : _GEN_3384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3386 = 8'h52 == total_offset_6 ? phv_data_82 : _GEN_3385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3387 = 8'h53 == total_offset_6 ? phv_data_83 : _GEN_3386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3388 = 8'h54 == total_offset_6 ? phv_data_84 : _GEN_3387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3389 = 8'h55 == total_offset_6 ? phv_data_85 : _GEN_3388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3390 = 8'h56 == total_offset_6 ? phv_data_86 : _GEN_3389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3391 = 8'h57 == total_offset_6 ? phv_data_87 : _GEN_3390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3392 = 8'h58 == total_offset_6 ? phv_data_88 : _GEN_3391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3393 = 8'h59 == total_offset_6 ? phv_data_89 : _GEN_3392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3394 = 8'h5a == total_offset_6 ? phv_data_90 : _GEN_3393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3395 = 8'h5b == total_offset_6 ? phv_data_91 : _GEN_3394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3396 = 8'h5c == total_offset_6 ? phv_data_92 : _GEN_3395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3397 = 8'h5d == total_offset_6 ? phv_data_93 : _GEN_3396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3398 = 8'h5e == total_offset_6 ? phv_data_94 : _GEN_3397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3399 = 8'h5f == total_offset_6 ? phv_data_95 : _GEN_3398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3400 = 8'h60 == total_offset_6 ? phv_data_96 : _GEN_3399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3401 = 8'h61 == total_offset_6 ? phv_data_97 : _GEN_3400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3402 = 8'h62 == total_offset_6 ? phv_data_98 : _GEN_3401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3403 = 8'h63 == total_offset_6 ? phv_data_99 : _GEN_3402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3404 = 8'h64 == total_offset_6 ? phv_data_100 : _GEN_3403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3405 = 8'h65 == total_offset_6 ? phv_data_101 : _GEN_3404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3406 = 8'h66 == total_offset_6 ? phv_data_102 : _GEN_3405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3407 = 8'h67 == total_offset_6 ? phv_data_103 : _GEN_3406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3408 = 8'h68 == total_offset_6 ? phv_data_104 : _GEN_3407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3409 = 8'h69 == total_offset_6 ? phv_data_105 : _GEN_3408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3410 = 8'h6a == total_offset_6 ? phv_data_106 : _GEN_3409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3411 = 8'h6b == total_offset_6 ? phv_data_107 : _GEN_3410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3412 = 8'h6c == total_offset_6 ? phv_data_108 : _GEN_3411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3413 = 8'h6d == total_offset_6 ? phv_data_109 : _GEN_3412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3414 = 8'h6e == total_offset_6 ? phv_data_110 : _GEN_3413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3415 = 8'h6f == total_offset_6 ? phv_data_111 : _GEN_3414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3416 = 8'h70 == total_offset_6 ? phv_data_112 : _GEN_3415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3417 = 8'h71 == total_offset_6 ? phv_data_113 : _GEN_3416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3418 = 8'h72 == total_offset_6 ? phv_data_114 : _GEN_3417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3419 = 8'h73 == total_offset_6 ? phv_data_115 : _GEN_3418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3420 = 8'h74 == total_offset_6 ? phv_data_116 : _GEN_3419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3421 = 8'h75 == total_offset_6 ? phv_data_117 : _GEN_3420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3422 = 8'h76 == total_offset_6 ? phv_data_118 : _GEN_3421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3423 = 8'h77 == total_offset_6 ? phv_data_119 : _GEN_3422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3424 = 8'h78 == total_offset_6 ? phv_data_120 : _GEN_3423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3425 = 8'h79 == total_offset_6 ? phv_data_121 : _GEN_3424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3426 = 8'h7a == total_offset_6 ? phv_data_122 : _GEN_3425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3427 = 8'h7b == total_offset_6 ? phv_data_123 : _GEN_3426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3428 = 8'h7c == total_offset_6 ? phv_data_124 : _GEN_3427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3429 = 8'h7d == total_offset_6 ? phv_data_125 : _GEN_3428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3430 = 8'h7e == total_offset_6 ? phv_data_126 : _GEN_3429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3431 = 8'h7f == total_offset_6 ? phv_data_127 : _GEN_3430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3432 = 8'h80 == total_offset_6 ? phv_data_128 : _GEN_3431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3433 = 8'h81 == total_offset_6 ? phv_data_129 : _GEN_3432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3434 = 8'h82 == total_offset_6 ? phv_data_130 : _GEN_3433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3435 = 8'h83 == total_offset_6 ? phv_data_131 : _GEN_3434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3436 = 8'h84 == total_offset_6 ? phv_data_132 : _GEN_3435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3437 = 8'h85 == total_offset_6 ? phv_data_133 : _GEN_3436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3438 = 8'h86 == total_offset_6 ? phv_data_134 : _GEN_3437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3439 = 8'h87 == total_offset_6 ? phv_data_135 : _GEN_3438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3440 = 8'h88 == total_offset_6 ? phv_data_136 : _GEN_3439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3441 = 8'h89 == total_offset_6 ? phv_data_137 : _GEN_3440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3442 = 8'h8a == total_offset_6 ? phv_data_138 : _GEN_3441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3443 = 8'h8b == total_offset_6 ? phv_data_139 : _GEN_3442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3444 = 8'h8c == total_offset_6 ? phv_data_140 : _GEN_3443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3445 = 8'h8d == total_offset_6 ? phv_data_141 : _GEN_3444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3446 = 8'h8e == total_offset_6 ? phv_data_142 : _GEN_3445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3447 = 8'h8f == total_offset_6 ? phv_data_143 : _GEN_3446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3448 = 8'h90 == total_offset_6 ? phv_data_144 : _GEN_3447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3449 = 8'h91 == total_offset_6 ? phv_data_145 : _GEN_3448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3450 = 8'h92 == total_offset_6 ? phv_data_146 : _GEN_3449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3451 = 8'h93 == total_offset_6 ? phv_data_147 : _GEN_3450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3452 = 8'h94 == total_offset_6 ? phv_data_148 : _GEN_3451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3453 = 8'h95 == total_offset_6 ? phv_data_149 : _GEN_3452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3454 = 8'h96 == total_offset_6 ? phv_data_150 : _GEN_3453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3455 = 8'h97 == total_offset_6 ? phv_data_151 : _GEN_3454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3456 = 8'h98 == total_offset_6 ? phv_data_152 : _GEN_3455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3457 = 8'h99 == total_offset_6 ? phv_data_153 : _GEN_3456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3458 = 8'h9a == total_offset_6 ? phv_data_154 : _GEN_3457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3459 = 8'h9b == total_offset_6 ? phv_data_155 : _GEN_3458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3460 = 8'h9c == total_offset_6 ? phv_data_156 : _GEN_3459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3461 = 8'h9d == total_offset_6 ? phv_data_157 : _GEN_3460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3462 = 8'h9e == total_offset_6 ? phv_data_158 : _GEN_3461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3463 = 8'h9f == total_offset_6 ? phv_data_159 : _GEN_3462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3464 = 8'ha0 == total_offset_6 ? phv_data_160 : _GEN_3463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3465 = 8'ha1 == total_offset_6 ? phv_data_161 : _GEN_3464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3466 = 8'ha2 == total_offset_6 ? phv_data_162 : _GEN_3465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3467 = 8'ha3 == total_offset_6 ? phv_data_163 : _GEN_3466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3468 = 8'ha4 == total_offset_6 ? phv_data_164 : _GEN_3467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3469 = 8'ha5 == total_offset_6 ? phv_data_165 : _GEN_3468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3470 = 8'ha6 == total_offset_6 ? phv_data_166 : _GEN_3469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3471 = 8'ha7 == total_offset_6 ? phv_data_167 : _GEN_3470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3472 = 8'ha8 == total_offset_6 ? phv_data_168 : _GEN_3471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3473 = 8'ha9 == total_offset_6 ? phv_data_169 : _GEN_3472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3474 = 8'haa == total_offset_6 ? phv_data_170 : _GEN_3473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3475 = 8'hab == total_offset_6 ? phv_data_171 : _GEN_3474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3476 = 8'hac == total_offset_6 ? phv_data_172 : _GEN_3475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3477 = 8'had == total_offset_6 ? phv_data_173 : _GEN_3476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3478 = 8'hae == total_offset_6 ? phv_data_174 : _GEN_3477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3479 = 8'haf == total_offset_6 ? phv_data_175 : _GEN_3478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3480 = 8'hb0 == total_offset_6 ? phv_data_176 : _GEN_3479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3481 = 8'hb1 == total_offset_6 ? phv_data_177 : _GEN_3480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3482 = 8'hb2 == total_offset_6 ? phv_data_178 : _GEN_3481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3483 = 8'hb3 == total_offset_6 ? phv_data_179 : _GEN_3482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3484 = 8'hb4 == total_offset_6 ? phv_data_180 : _GEN_3483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3485 = 8'hb5 == total_offset_6 ? phv_data_181 : _GEN_3484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3486 = 8'hb6 == total_offset_6 ? phv_data_182 : _GEN_3485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3487 = 8'hb7 == total_offset_6 ? phv_data_183 : _GEN_3486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3488 = 8'hb8 == total_offset_6 ? phv_data_184 : _GEN_3487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3489 = 8'hb9 == total_offset_6 ? phv_data_185 : _GEN_3488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3490 = 8'hba == total_offset_6 ? phv_data_186 : _GEN_3489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3491 = 8'hbb == total_offset_6 ? phv_data_187 : _GEN_3490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3492 = 8'hbc == total_offset_6 ? phv_data_188 : _GEN_3491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3493 = 8'hbd == total_offset_6 ? phv_data_189 : _GEN_3492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3494 = 8'hbe == total_offset_6 ? phv_data_190 : _GEN_3493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3495 = 8'hbf == total_offset_6 ? phv_data_191 : _GEN_3494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3496 = 8'hc0 == total_offset_6 ? phv_data_192 : _GEN_3495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3497 = 8'hc1 == total_offset_6 ? phv_data_193 : _GEN_3496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3498 = 8'hc2 == total_offset_6 ? phv_data_194 : _GEN_3497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3499 = 8'hc3 == total_offset_6 ? phv_data_195 : _GEN_3498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3500 = 8'hc4 == total_offset_6 ? phv_data_196 : _GEN_3499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3501 = 8'hc5 == total_offset_6 ? phv_data_197 : _GEN_3500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3502 = 8'hc6 == total_offset_6 ? phv_data_198 : _GEN_3501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3503 = 8'hc7 == total_offset_6 ? phv_data_199 : _GEN_3502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3504 = 8'hc8 == total_offset_6 ? phv_data_200 : _GEN_3503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3505 = 8'hc9 == total_offset_6 ? phv_data_201 : _GEN_3504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3506 = 8'hca == total_offset_6 ? phv_data_202 : _GEN_3505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3507 = 8'hcb == total_offset_6 ? phv_data_203 : _GEN_3506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3508 = 8'hcc == total_offset_6 ? phv_data_204 : _GEN_3507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3509 = 8'hcd == total_offset_6 ? phv_data_205 : _GEN_3508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3510 = 8'hce == total_offset_6 ? phv_data_206 : _GEN_3509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3511 = 8'hcf == total_offset_6 ? phv_data_207 : _GEN_3510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3512 = 8'hd0 == total_offset_6 ? phv_data_208 : _GEN_3511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3513 = 8'hd1 == total_offset_6 ? phv_data_209 : _GEN_3512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3514 = 8'hd2 == total_offset_6 ? phv_data_210 : _GEN_3513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3515 = 8'hd3 == total_offset_6 ? phv_data_211 : _GEN_3514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3516 = 8'hd4 == total_offset_6 ? phv_data_212 : _GEN_3515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3517 = 8'hd5 == total_offset_6 ? phv_data_213 : _GEN_3516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3518 = 8'hd6 == total_offset_6 ? phv_data_214 : _GEN_3517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3519 = 8'hd7 == total_offset_6 ? phv_data_215 : _GEN_3518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3520 = 8'hd8 == total_offset_6 ? phv_data_216 : _GEN_3519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3521 = 8'hd9 == total_offset_6 ? phv_data_217 : _GEN_3520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3522 = 8'hda == total_offset_6 ? phv_data_218 : _GEN_3521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3523 = 8'hdb == total_offset_6 ? phv_data_219 : _GEN_3522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3524 = 8'hdc == total_offset_6 ? phv_data_220 : _GEN_3523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3525 = 8'hdd == total_offset_6 ? phv_data_221 : _GEN_3524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3526 = 8'hde == total_offset_6 ? phv_data_222 : _GEN_3525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3527 = 8'hdf == total_offset_6 ? phv_data_223 : _GEN_3526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3528 = 8'he0 == total_offset_6 ? phv_data_224 : _GEN_3527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3529 = 8'he1 == total_offset_6 ? phv_data_225 : _GEN_3528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3530 = 8'he2 == total_offset_6 ? phv_data_226 : _GEN_3529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3531 = 8'he3 == total_offset_6 ? phv_data_227 : _GEN_3530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3532 = 8'he4 == total_offset_6 ? phv_data_228 : _GEN_3531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3533 = 8'he5 == total_offset_6 ? phv_data_229 : _GEN_3532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3534 = 8'he6 == total_offset_6 ? phv_data_230 : _GEN_3533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3535 = 8'he7 == total_offset_6 ? phv_data_231 : _GEN_3534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3536 = 8'he8 == total_offset_6 ? phv_data_232 : _GEN_3535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3537 = 8'he9 == total_offset_6 ? phv_data_233 : _GEN_3536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3538 = 8'hea == total_offset_6 ? phv_data_234 : _GEN_3537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3539 = 8'heb == total_offset_6 ? phv_data_235 : _GEN_3538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3540 = 8'hec == total_offset_6 ? phv_data_236 : _GEN_3539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3541 = 8'hed == total_offset_6 ? phv_data_237 : _GEN_3540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3542 = 8'hee == total_offset_6 ? phv_data_238 : _GEN_3541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3543 = 8'hef == total_offset_6 ? phv_data_239 : _GEN_3542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3544 = 8'hf0 == total_offset_6 ? phv_data_240 : _GEN_3543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3545 = 8'hf1 == total_offset_6 ? phv_data_241 : _GEN_3544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3546 = 8'hf2 == total_offset_6 ? phv_data_242 : _GEN_3545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3547 = 8'hf3 == total_offset_6 ? phv_data_243 : _GEN_3546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3548 = 8'hf4 == total_offset_6 ? phv_data_244 : _GEN_3547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3549 = 8'hf5 == total_offset_6 ? phv_data_245 : _GEN_3548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3550 = 8'hf6 == total_offset_6 ? phv_data_246 : _GEN_3549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3551 = 8'hf7 == total_offset_6 ? phv_data_247 : _GEN_3550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3552 = 8'hf8 == total_offset_6 ? phv_data_248 : _GEN_3551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3553 = 8'hf9 == total_offset_6 ? phv_data_249 : _GEN_3552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3554 = 8'hfa == total_offset_6 ? phv_data_250 : _GEN_3553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3555 = 8'hfb == total_offset_6 ? phv_data_251 : _GEN_3554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3556 = 8'hfc == total_offset_6 ? phv_data_252 : _GEN_3555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3557 = 8'hfd == total_offset_6 ? phv_data_253 : _GEN_3556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3558 = 8'hfe == total_offset_6 ? phv_data_254 : _GEN_3557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3559 = 8'hff == total_offset_6 ? phv_data_255 : _GEN_3558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_10664 = {{1'd0}, total_offset_6}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3560 = 9'h100 == _GEN_10664 ? phv_data_256 : _GEN_3559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3561 = 9'h101 == _GEN_10664 ? phv_data_257 : _GEN_3560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3562 = 9'h102 == _GEN_10664 ? phv_data_258 : _GEN_3561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3563 = 9'h103 == _GEN_10664 ? phv_data_259 : _GEN_3562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3564 = 9'h104 == _GEN_10664 ? phv_data_260 : _GEN_3563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3565 = 9'h105 == _GEN_10664 ? phv_data_261 : _GEN_3564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3566 = 9'h106 == _GEN_10664 ? phv_data_262 : _GEN_3565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3567 = 9'h107 == _GEN_10664 ? phv_data_263 : _GEN_3566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3568 = 9'h108 == _GEN_10664 ? phv_data_264 : _GEN_3567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3569 = 9'h109 == _GEN_10664 ? phv_data_265 : _GEN_3568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3570 = 9'h10a == _GEN_10664 ? phv_data_266 : _GEN_3569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3571 = 9'h10b == _GEN_10664 ? phv_data_267 : _GEN_3570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3572 = 9'h10c == _GEN_10664 ? phv_data_268 : _GEN_3571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3573 = 9'h10d == _GEN_10664 ? phv_data_269 : _GEN_3572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3574 = 9'h10e == _GEN_10664 ? phv_data_270 : _GEN_3573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3575 = 9'h10f == _GEN_10664 ? phv_data_271 : _GEN_3574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3576 = 9'h110 == _GEN_10664 ? phv_data_272 : _GEN_3575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3577 = 9'h111 == _GEN_10664 ? phv_data_273 : _GEN_3576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3578 = 9'h112 == _GEN_10664 ? phv_data_274 : _GEN_3577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3579 = 9'h113 == _GEN_10664 ? phv_data_275 : _GEN_3578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3580 = 9'h114 == _GEN_10664 ? phv_data_276 : _GEN_3579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3581 = 9'h115 == _GEN_10664 ? phv_data_277 : _GEN_3580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3582 = 9'h116 == _GEN_10664 ? phv_data_278 : _GEN_3581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3583 = 9'h117 == _GEN_10664 ? phv_data_279 : _GEN_3582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3584 = 9'h118 == _GEN_10664 ? phv_data_280 : _GEN_3583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3585 = 9'h119 == _GEN_10664 ? phv_data_281 : _GEN_3584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3586 = 9'h11a == _GEN_10664 ? phv_data_282 : _GEN_3585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3587 = 9'h11b == _GEN_10664 ? phv_data_283 : _GEN_3586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3588 = 9'h11c == _GEN_10664 ? phv_data_284 : _GEN_3587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3589 = 9'h11d == _GEN_10664 ? phv_data_285 : _GEN_3588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3590 = 9'h11e == _GEN_10664 ? phv_data_286 : _GEN_3589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3591 = 9'h11f == _GEN_10664 ? phv_data_287 : _GEN_3590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3592 = 9'h120 == _GEN_10664 ? phv_data_288 : _GEN_3591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3593 = 9'h121 == _GEN_10664 ? phv_data_289 : _GEN_3592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3594 = 9'h122 == _GEN_10664 ? phv_data_290 : _GEN_3593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3595 = 9'h123 == _GEN_10664 ? phv_data_291 : _GEN_3594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3596 = 9'h124 == _GEN_10664 ? phv_data_292 : _GEN_3595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3597 = 9'h125 == _GEN_10664 ? phv_data_293 : _GEN_3596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3598 = 9'h126 == _GEN_10664 ? phv_data_294 : _GEN_3597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3599 = 9'h127 == _GEN_10664 ? phv_data_295 : _GEN_3598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3600 = 9'h128 == _GEN_10664 ? phv_data_296 : _GEN_3599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3601 = 9'h129 == _GEN_10664 ? phv_data_297 : _GEN_3600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3602 = 9'h12a == _GEN_10664 ? phv_data_298 : _GEN_3601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3603 = 9'h12b == _GEN_10664 ? phv_data_299 : _GEN_3602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3604 = 9'h12c == _GEN_10664 ? phv_data_300 : _GEN_3603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3605 = 9'h12d == _GEN_10664 ? phv_data_301 : _GEN_3604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3606 = 9'h12e == _GEN_10664 ? phv_data_302 : _GEN_3605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3607 = 9'h12f == _GEN_10664 ? phv_data_303 : _GEN_3606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3608 = 9'h130 == _GEN_10664 ? phv_data_304 : _GEN_3607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3609 = 9'h131 == _GEN_10664 ? phv_data_305 : _GEN_3608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3610 = 9'h132 == _GEN_10664 ? phv_data_306 : _GEN_3609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3611 = 9'h133 == _GEN_10664 ? phv_data_307 : _GEN_3610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3612 = 9'h134 == _GEN_10664 ? phv_data_308 : _GEN_3611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3613 = 9'h135 == _GEN_10664 ? phv_data_309 : _GEN_3612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3614 = 9'h136 == _GEN_10664 ? phv_data_310 : _GEN_3613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3615 = 9'h137 == _GEN_10664 ? phv_data_311 : _GEN_3614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3616 = 9'h138 == _GEN_10664 ? phv_data_312 : _GEN_3615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3617 = 9'h139 == _GEN_10664 ? phv_data_313 : _GEN_3616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3618 = 9'h13a == _GEN_10664 ? phv_data_314 : _GEN_3617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3619 = 9'h13b == _GEN_10664 ? phv_data_315 : _GEN_3618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3620 = 9'h13c == _GEN_10664 ? phv_data_316 : _GEN_3619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3621 = 9'h13d == _GEN_10664 ? phv_data_317 : _GEN_3620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3622 = 9'h13e == _GEN_10664 ? phv_data_318 : _GEN_3621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3623 = 9'h13f == _GEN_10664 ? phv_data_319 : _GEN_3622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3624 = 9'h140 == _GEN_10664 ? phv_data_320 : _GEN_3623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3625 = 9'h141 == _GEN_10664 ? phv_data_321 : _GEN_3624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3626 = 9'h142 == _GEN_10664 ? phv_data_322 : _GEN_3625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3627 = 9'h143 == _GEN_10664 ? phv_data_323 : _GEN_3626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3628 = 9'h144 == _GEN_10664 ? phv_data_324 : _GEN_3627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3629 = 9'h145 == _GEN_10664 ? phv_data_325 : _GEN_3628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3630 = 9'h146 == _GEN_10664 ? phv_data_326 : _GEN_3629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3631 = 9'h147 == _GEN_10664 ? phv_data_327 : _GEN_3630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3632 = 9'h148 == _GEN_10664 ? phv_data_328 : _GEN_3631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3633 = 9'h149 == _GEN_10664 ? phv_data_329 : _GEN_3632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3634 = 9'h14a == _GEN_10664 ? phv_data_330 : _GEN_3633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3635 = 9'h14b == _GEN_10664 ? phv_data_331 : _GEN_3634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3636 = 9'h14c == _GEN_10664 ? phv_data_332 : _GEN_3635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3637 = 9'h14d == _GEN_10664 ? phv_data_333 : _GEN_3636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3638 = 9'h14e == _GEN_10664 ? phv_data_334 : _GEN_3637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3639 = 9'h14f == _GEN_10664 ? phv_data_335 : _GEN_3638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3640 = 9'h150 == _GEN_10664 ? phv_data_336 : _GEN_3639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3641 = 9'h151 == _GEN_10664 ? phv_data_337 : _GEN_3640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3642 = 9'h152 == _GEN_10664 ? phv_data_338 : _GEN_3641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3643 = 9'h153 == _GEN_10664 ? phv_data_339 : _GEN_3642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3644 = 9'h154 == _GEN_10664 ? phv_data_340 : _GEN_3643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3645 = 9'h155 == _GEN_10664 ? phv_data_341 : _GEN_3644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3646 = 9'h156 == _GEN_10664 ? phv_data_342 : _GEN_3645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3647 = 9'h157 == _GEN_10664 ? phv_data_343 : _GEN_3646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3648 = 9'h158 == _GEN_10664 ? phv_data_344 : _GEN_3647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3649 = 9'h159 == _GEN_10664 ? phv_data_345 : _GEN_3648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3650 = 9'h15a == _GEN_10664 ? phv_data_346 : _GEN_3649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3651 = 9'h15b == _GEN_10664 ? phv_data_347 : _GEN_3650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3652 = 9'h15c == _GEN_10664 ? phv_data_348 : _GEN_3651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3653 = 9'h15d == _GEN_10664 ? phv_data_349 : _GEN_3652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3654 = 9'h15e == _GEN_10664 ? phv_data_350 : _GEN_3653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3655 = 9'h15f == _GEN_10664 ? phv_data_351 : _GEN_3654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3656 = 9'h160 == _GEN_10664 ? phv_data_352 : _GEN_3655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3657 = 9'h161 == _GEN_10664 ? phv_data_353 : _GEN_3656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3658 = 9'h162 == _GEN_10664 ? phv_data_354 : _GEN_3657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3659 = 9'h163 == _GEN_10664 ? phv_data_355 : _GEN_3658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3660 = 9'h164 == _GEN_10664 ? phv_data_356 : _GEN_3659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3661 = 9'h165 == _GEN_10664 ? phv_data_357 : _GEN_3660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3662 = 9'h166 == _GEN_10664 ? phv_data_358 : _GEN_3661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3663 = 9'h167 == _GEN_10664 ? phv_data_359 : _GEN_3662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3664 = 9'h168 == _GEN_10664 ? phv_data_360 : _GEN_3663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3665 = 9'h169 == _GEN_10664 ? phv_data_361 : _GEN_3664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3666 = 9'h16a == _GEN_10664 ? phv_data_362 : _GEN_3665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3667 = 9'h16b == _GEN_10664 ? phv_data_363 : _GEN_3666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3668 = 9'h16c == _GEN_10664 ? phv_data_364 : _GEN_3667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3669 = 9'h16d == _GEN_10664 ? phv_data_365 : _GEN_3668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3670 = 9'h16e == _GEN_10664 ? phv_data_366 : _GEN_3669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3671 = 9'h16f == _GEN_10664 ? phv_data_367 : _GEN_3670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3672 = 9'h170 == _GEN_10664 ? phv_data_368 : _GEN_3671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3673 = 9'h171 == _GEN_10664 ? phv_data_369 : _GEN_3672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3674 = 9'h172 == _GEN_10664 ? phv_data_370 : _GEN_3673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3675 = 9'h173 == _GEN_10664 ? phv_data_371 : _GEN_3674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3676 = 9'h174 == _GEN_10664 ? phv_data_372 : _GEN_3675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3677 = 9'h175 == _GEN_10664 ? phv_data_373 : _GEN_3676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3678 = 9'h176 == _GEN_10664 ? phv_data_374 : _GEN_3677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3679 = 9'h177 == _GEN_10664 ? phv_data_375 : _GEN_3678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3680 = 9'h178 == _GEN_10664 ? phv_data_376 : _GEN_3679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3681 = 9'h179 == _GEN_10664 ? phv_data_377 : _GEN_3680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3682 = 9'h17a == _GEN_10664 ? phv_data_378 : _GEN_3681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3683 = 9'h17b == _GEN_10664 ? phv_data_379 : _GEN_3682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3684 = 9'h17c == _GEN_10664 ? phv_data_380 : _GEN_3683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3685 = 9'h17d == _GEN_10664 ? phv_data_381 : _GEN_3684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3686 = 9'h17e == _GEN_10664 ? phv_data_382 : _GEN_3685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3687 = 9'h17f == _GEN_10664 ? phv_data_383 : _GEN_3686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3688 = 9'h180 == _GEN_10664 ? phv_data_384 : _GEN_3687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3689 = 9'h181 == _GEN_10664 ? phv_data_385 : _GEN_3688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3690 = 9'h182 == _GEN_10664 ? phv_data_386 : _GEN_3689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3691 = 9'h183 == _GEN_10664 ? phv_data_387 : _GEN_3690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3692 = 9'h184 == _GEN_10664 ? phv_data_388 : _GEN_3691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3693 = 9'h185 == _GEN_10664 ? phv_data_389 : _GEN_3692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3694 = 9'h186 == _GEN_10664 ? phv_data_390 : _GEN_3693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3695 = 9'h187 == _GEN_10664 ? phv_data_391 : _GEN_3694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3696 = 9'h188 == _GEN_10664 ? phv_data_392 : _GEN_3695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3697 = 9'h189 == _GEN_10664 ? phv_data_393 : _GEN_3696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3698 = 9'h18a == _GEN_10664 ? phv_data_394 : _GEN_3697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3699 = 9'h18b == _GEN_10664 ? phv_data_395 : _GEN_3698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3700 = 9'h18c == _GEN_10664 ? phv_data_396 : _GEN_3699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3701 = 9'h18d == _GEN_10664 ? phv_data_397 : _GEN_3700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3702 = 9'h18e == _GEN_10664 ? phv_data_398 : _GEN_3701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3703 = 9'h18f == _GEN_10664 ? phv_data_399 : _GEN_3702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3704 = 9'h190 == _GEN_10664 ? phv_data_400 : _GEN_3703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3705 = 9'h191 == _GEN_10664 ? phv_data_401 : _GEN_3704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3706 = 9'h192 == _GEN_10664 ? phv_data_402 : _GEN_3705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3707 = 9'h193 == _GEN_10664 ? phv_data_403 : _GEN_3706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3708 = 9'h194 == _GEN_10664 ? phv_data_404 : _GEN_3707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3709 = 9'h195 == _GEN_10664 ? phv_data_405 : _GEN_3708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3710 = 9'h196 == _GEN_10664 ? phv_data_406 : _GEN_3709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3711 = 9'h197 == _GEN_10664 ? phv_data_407 : _GEN_3710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3712 = 9'h198 == _GEN_10664 ? phv_data_408 : _GEN_3711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3713 = 9'h199 == _GEN_10664 ? phv_data_409 : _GEN_3712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3714 = 9'h19a == _GEN_10664 ? phv_data_410 : _GEN_3713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3715 = 9'h19b == _GEN_10664 ? phv_data_411 : _GEN_3714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3716 = 9'h19c == _GEN_10664 ? phv_data_412 : _GEN_3715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3717 = 9'h19d == _GEN_10664 ? phv_data_413 : _GEN_3716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3718 = 9'h19e == _GEN_10664 ? phv_data_414 : _GEN_3717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3719 = 9'h19f == _GEN_10664 ? phv_data_415 : _GEN_3718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3720 = 9'h1a0 == _GEN_10664 ? phv_data_416 : _GEN_3719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3721 = 9'h1a1 == _GEN_10664 ? phv_data_417 : _GEN_3720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3722 = 9'h1a2 == _GEN_10664 ? phv_data_418 : _GEN_3721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3723 = 9'h1a3 == _GEN_10664 ? phv_data_419 : _GEN_3722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3724 = 9'h1a4 == _GEN_10664 ? phv_data_420 : _GEN_3723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3725 = 9'h1a5 == _GEN_10664 ? phv_data_421 : _GEN_3724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3726 = 9'h1a6 == _GEN_10664 ? phv_data_422 : _GEN_3725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3727 = 9'h1a7 == _GEN_10664 ? phv_data_423 : _GEN_3726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3728 = 9'h1a8 == _GEN_10664 ? phv_data_424 : _GEN_3727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3729 = 9'h1a9 == _GEN_10664 ? phv_data_425 : _GEN_3728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3730 = 9'h1aa == _GEN_10664 ? phv_data_426 : _GEN_3729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3731 = 9'h1ab == _GEN_10664 ? phv_data_427 : _GEN_3730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3732 = 9'h1ac == _GEN_10664 ? phv_data_428 : _GEN_3731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3733 = 9'h1ad == _GEN_10664 ? phv_data_429 : _GEN_3732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3734 = 9'h1ae == _GEN_10664 ? phv_data_430 : _GEN_3733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3735 = 9'h1af == _GEN_10664 ? phv_data_431 : _GEN_3734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3736 = 9'h1b0 == _GEN_10664 ? phv_data_432 : _GEN_3735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3737 = 9'h1b1 == _GEN_10664 ? phv_data_433 : _GEN_3736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3738 = 9'h1b2 == _GEN_10664 ? phv_data_434 : _GEN_3737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3739 = 9'h1b3 == _GEN_10664 ? phv_data_435 : _GEN_3738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3740 = 9'h1b4 == _GEN_10664 ? phv_data_436 : _GEN_3739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3741 = 9'h1b5 == _GEN_10664 ? phv_data_437 : _GEN_3740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3742 = 9'h1b6 == _GEN_10664 ? phv_data_438 : _GEN_3741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3743 = 9'h1b7 == _GEN_10664 ? phv_data_439 : _GEN_3742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3744 = 9'h1b8 == _GEN_10664 ? phv_data_440 : _GEN_3743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3745 = 9'h1b9 == _GEN_10664 ? phv_data_441 : _GEN_3744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3746 = 9'h1ba == _GEN_10664 ? phv_data_442 : _GEN_3745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3747 = 9'h1bb == _GEN_10664 ? phv_data_443 : _GEN_3746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3748 = 9'h1bc == _GEN_10664 ? phv_data_444 : _GEN_3747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3749 = 9'h1bd == _GEN_10664 ? phv_data_445 : _GEN_3748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3750 = 9'h1be == _GEN_10664 ? phv_data_446 : _GEN_3749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3751 = 9'h1bf == _GEN_10664 ? phv_data_447 : _GEN_3750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3752 = 9'h1c0 == _GEN_10664 ? phv_data_448 : _GEN_3751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3753 = 9'h1c1 == _GEN_10664 ? phv_data_449 : _GEN_3752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3754 = 9'h1c2 == _GEN_10664 ? phv_data_450 : _GEN_3753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3755 = 9'h1c3 == _GEN_10664 ? phv_data_451 : _GEN_3754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3756 = 9'h1c4 == _GEN_10664 ? phv_data_452 : _GEN_3755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3757 = 9'h1c5 == _GEN_10664 ? phv_data_453 : _GEN_3756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3758 = 9'h1c6 == _GEN_10664 ? phv_data_454 : _GEN_3757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3759 = 9'h1c7 == _GEN_10664 ? phv_data_455 : _GEN_3758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3760 = 9'h1c8 == _GEN_10664 ? phv_data_456 : _GEN_3759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3761 = 9'h1c9 == _GEN_10664 ? phv_data_457 : _GEN_3760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3762 = 9'h1ca == _GEN_10664 ? phv_data_458 : _GEN_3761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3763 = 9'h1cb == _GEN_10664 ? phv_data_459 : _GEN_3762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3764 = 9'h1cc == _GEN_10664 ? phv_data_460 : _GEN_3763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3765 = 9'h1cd == _GEN_10664 ? phv_data_461 : _GEN_3764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3766 = 9'h1ce == _GEN_10664 ? phv_data_462 : _GEN_3765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3767 = 9'h1cf == _GEN_10664 ? phv_data_463 : _GEN_3766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3768 = 9'h1d0 == _GEN_10664 ? phv_data_464 : _GEN_3767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3769 = 9'h1d1 == _GEN_10664 ? phv_data_465 : _GEN_3768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3770 = 9'h1d2 == _GEN_10664 ? phv_data_466 : _GEN_3769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3771 = 9'h1d3 == _GEN_10664 ? phv_data_467 : _GEN_3770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3772 = 9'h1d4 == _GEN_10664 ? phv_data_468 : _GEN_3771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3773 = 9'h1d5 == _GEN_10664 ? phv_data_469 : _GEN_3772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3774 = 9'h1d6 == _GEN_10664 ? phv_data_470 : _GEN_3773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3775 = 9'h1d7 == _GEN_10664 ? phv_data_471 : _GEN_3774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3776 = 9'h1d8 == _GEN_10664 ? phv_data_472 : _GEN_3775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3777 = 9'h1d9 == _GEN_10664 ? phv_data_473 : _GEN_3776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3778 = 9'h1da == _GEN_10664 ? phv_data_474 : _GEN_3777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3779 = 9'h1db == _GEN_10664 ? phv_data_475 : _GEN_3778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3780 = 9'h1dc == _GEN_10664 ? phv_data_476 : _GEN_3779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3781 = 9'h1dd == _GEN_10664 ? phv_data_477 : _GEN_3780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3782 = 9'h1de == _GEN_10664 ? phv_data_478 : _GEN_3781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3783 = 9'h1df == _GEN_10664 ? phv_data_479 : _GEN_3782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3784 = 9'h1e0 == _GEN_10664 ? phv_data_480 : _GEN_3783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3785 = 9'h1e1 == _GEN_10664 ? phv_data_481 : _GEN_3784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3786 = 9'h1e2 == _GEN_10664 ? phv_data_482 : _GEN_3785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3787 = 9'h1e3 == _GEN_10664 ? phv_data_483 : _GEN_3786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3788 = 9'h1e4 == _GEN_10664 ? phv_data_484 : _GEN_3787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3789 = 9'h1e5 == _GEN_10664 ? phv_data_485 : _GEN_3788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3790 = 9'h1e6 == _GEN_10664 ? phv_data_486 : _GEN_3789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3791 = 9'h1e7 == _GEN_10664 ? phv_data_487 : _GEN_3790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3792 = 9'h1e8 == _GEN_10664 ? phv_data_488 : _GEN_3791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3793 = 9'h1e9 == _GEN_10664 ? phv_data_489 : _GEN_3792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3794 = 9'h1ea == _GEN_10664 ? phv_data_490 : _GEN_3793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3795 = 9'h1eb == _GEN_10664 ? phv_data_491 : _GEN_3794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3796 = 9'h1ec == _GEN_10664 ? phv_data_492 : _GEN_3795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3797 = 9'h1ed == _GEN_10664 ? phv_data_493 : _GEN_3796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3798 = 9'h1ee == _GEN_10664 ? phv_data_494 : _GEN_3797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3799 = 9'h1ef == _GEN_10664 ? phv_data_495 : _GEN_3798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3800 = 9'h1f0 == _GEN_10664 ? phv_data_496 : _GEN_3799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3801 = 9'h1f1 == _GEN_10664 ? phv_data_497 : _GEN_3800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3802 = 9'h1f2 == _GEN_10664 ? phv_data_498 : _GEN_3801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3803 = 9'h1f3 == _GEN_10664 ? phv_data_499 : _GEN_3802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3804 = 9'h1f4 == _GEN_10664 ? phv_data_500 : _GEN_3803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3805 = 9'h1f5 == _GEN_10664 ? phv_data_501 : _GEN_3804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3806 = 9'h1f6 == _GEN_10664 ? phv_data_502 : _GEN_3805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3807 = 9'h1f7 == _GEN_10664 ? phv_data_503 : _GEN_3806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3808 = 9'h1f8 == _GEN_10664 ? phv_data_504 : _GEN_3807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3809 = 9'h1f9 == _GEN_10664 ? phv_data_505 : _GEN_3808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3810 = 9'h1fa == _GEN_10664 ? phv_data_506 : _GEN_3809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3811 = 9'h1fb == _GEN_10664 ? phv_data_507 : _GEN_3810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3812 = 9'h1fc == _GEN_10664 ? phv_data_508 : _GEN_3811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3813 = 9'h1fd == _GEN_10664 ? phv_data_509 : _GEN_3812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3814 = 9'h1fe == _GEN_10664 ? phv_data_510 : _GEN_3813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_1 = 9'h1ff == _GEN_10664 ? phv_data_511 : _GEN_3814; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_1_1 = 2'h2 >= offset_1[1:0] & (2'h2 < ending_1 | ending_1 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_7 = {total_offset_hi_1,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_3817 = 8'h1 == total_offset_7 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3818 = 8'h2 == total_offset_7 ? phv_data_2 : _GEN_3817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3819 = 8'h3 == total_offset_7 ? phv_data_3 : _GEN_3818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3820 = 8'h4 == total_offset_7 ? phv_data_4 : _GEN_3819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3821 = 8'h5 == total_offset_7 ? phv_data_5 : _GEN_3820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3822 = 8'h6 == total_offset_7 ? phv_data_6 : _GEN_3821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3823 = 8'h7 == total_offset_7 ? phv_data_7 : _GEN_3822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3824 = 8'h8 == total_offset_7 ? phv_data_8 : _GEN_3823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3825 = 8'h9 == total_offset_7 ? phv_data_9 : _GEN_3824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3826 = 8'ha == total_offset_7 ? phv_data_10 : _GEN_3825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3827 = 8'hb == total_offset_7 ? phv_data_11 : _GEN_3826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3828 = 8'hc == total_offset_7 ? phv_data_12 : _GEN_3827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3829 = 8'hd == total_offset_7 ? phv_data_13 : _GEN_3828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3830 = 8'he == total_offset_7 ? phv_data_14 : _GEN_3829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3831 = 8'hf == total_offset_7 ? phv_data_15 : _GEN_3830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3832 = 8'h10 == total_offset_7 ? phv_data_16 : _GEN_3831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3833 = 8'h11 == total_offset_7 ? phv_data_17 : _GEN_3832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3834 = 8'h12 == total_offset_7 ? phv_data_18 : _GEN_3833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3835 = 8'h13 == total_offset_7 ? phv_data_19 : _GEN_3834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3836 = 8'h14 == total_offset_7 ? phv_data_20 : _GEN_3835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3837 = 8'h15 == total_offset_7 ? phv_data_21 : _GEN_3836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3838 = 8'h16 == total_offset_7 ? phv_data_22 : _GEN_3837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3839 = 8'h17 == total_offset_7 ? phv_data_23 : _GEN_3838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3840 = 8'h18 == total_offset_7 ? phv_data_24 : _GEN_3839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3841 = 8'h19 == total_offset_7 ? phv_data_25 : _GEN_3840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3842 = 8'h1a == total_offset_7 ? phv_data_26 : _GEN_3841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3843 = 8'h1b == total_offset_7 ? phv_data_27 : _GEN_3842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3844 = 8'h1c == total_offset_7 ? phv_data_28 : _GEN_3843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3845 = 8'h1d == total_offset_7 ? phv_data_29 : _GEN_3844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3846 = 8'h1e == total_offset_7 ? phv_data_30 : _GEN_3845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3847 = 8'h1f == total_offset_7 ? phv_data_31 : _GEN_3846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3848 = 8'h20 == total_offset_7 ? phv_data_32 : _GEN_3847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3849 = 8'h21 == total_offset_7 ? phv_data_33 : _GEN_3848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3850 = 8'h22 == total_offset_7 ? phv_data_34 : _GEN_3849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3851 = 8'h23 == total_offset_7 ? phv_data_35 : _GEN_3850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3852 = 8'h24 == total_offset_7 ? phv_data_36 : _GEN_3851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3853 = 8'h25 == total_offset_7 ? phv_data_37 : _GEN_3852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3854 = 8'h26 == total_offset_7 ? phv_data_38 : _GEN_3853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3855 = 8'h27 == total_offset_7 ? phv_data_39 : _GEN_3854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3856 = 8'h28 == total_offset_7 ? phv_data_40 : _GEN_3855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3857 = 8'h29 == total_offset_7 ? phv_data_41 : _GEN_3856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3858 = 8'h2a == total_offset_7 ? phv_data_42 : _GEN_3857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3859 = 8'h2b == total_offset_7 ? phv_data_43 : _GEN_3858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3860 = 8'h2c == total_offset_7 ? phv_data_44 : _GEN_3859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3861 = 8'h2d == total_offset_7 ? phv_data_45 : _GEN_3860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3862 = 8'h2e == total_offset_7 ? phv_data_46 : _GEN_3861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3863 = 8'h2f == total_offset_7 ? phv_data_47 : _GEN_3862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3864 = 8'h30 == total_offset_7 ? phv_data_48 : _GEN_3863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3865 = 8'h31 == total_offset_7 ? phv_data_49 : _GEN_3864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3866 = 8'h32 == total_offset_7 ? phv_data_50 : _GEN_3865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3867 = 8'h33 == total_offset_7 ? phv_data_51 : _GEN_3866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3868 = 8'h34 == total_offset_7 ? phv_data_52 : _GEN_3867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3869 = 8'h35 == total_offset_7 ? phv_data_53 : _GEN_3868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3870 = 8'h36 == total_offset_7 ? phv_data_54 : _GEN_3869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3871 = 8'h37 == total_offset_7 ? phv_data_55 : _GEN_3870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3872 = 8'h38 == total_offset_7 ? phv_data_56 : _GEN_3871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3873 = 8'h39 == total_offset_7 ? phv_data_57 : _GEN_3872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3874 = 8'h3a == total_offset_7 ? phv_data_58 : _GEN_3873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3875 = 8'h3b == total_offset_7 ? phv_data_59 : _GEN_3874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3876 = 8'h3c == total_offset_7 ? phv_data_60 : _GEN_3875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3877 = 8'h3d == total_offset_7 ? phv_data_61 : _GEN_3876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3878 = 8'h3e == total_offset_7 ? phv_data_62 : _GEN_3877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3879 = 8'h3f == total_offset_7 ? phv_data_63 : _GEN_3878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3880 = 8'h40 == total_offset_7 ? phv_data_64 : _GEN_3879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3881 = 8'h41 == total_offset_7 ? phv_data_65 : _GEN_3880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3882 = 8'h42 == total_offset_7 ? phv_data_66 : _GEN_3881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3883 = 8'h43 == total_offset_7 ? phv_data_67 : _GEN_3882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3884 = 8'h44 == total_offset_7 ? phv_data_68 : _GEN_3883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3885 = 8'h45 == total_offset_7 ? phv_data_69 : _GEN_3884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3886 = 8'h46 == total_offset_7 ? phv_data_70 : _GEN_3885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3887 = 8'h47 == total_offset_7 ? phv_data_71 : _GEN_3886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3888 = 8'h48 == total_offset_7 ? phv_data_72 : _GEN_3887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3889 = 8'h49 == total_offset_7 ? phv_data_73 : _GEN_3888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3890 = 8'h4a == total_offset_7 ? phv_data_74 : _GEN_3889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3891 = 8'h4b == total_offset_7 ? phv_data_75 : _GEN_3890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3892 = 8'h4c == total_offset_7 ? phv_data_76 : _GEN_3891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3893 = 8'h4d == total_offset_7 ? phv_data_77 : _GEN_3892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3894 = 8'h4e == total_offset_7 ? phv_data_78 : _GEN_3893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3895 = 8'h4f == total_offset_7 ? phv_data_79 : _GEN_3894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3896 = 8'h50 == total_offset_7 ? phv_data_80 : _GEN_3895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3897 = 8'h51 == total_offset_7 ? phv_data_81 : _GEN_3896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3898 = 8'h52 == total_offset_7 ? phv_data_82 : _GEN_3897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3899 = 8'h53 == total_offset_7 ? phv_data_83 : _GEN_3898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3900 = 8'h54 == total_offset_7 ? phv_data_84 : _GEN_3899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3901 = 8'h55 == total_offset_7 ? phv_data_85 : _GEN_3900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3902 = 8'h56 == total_offset_7 ? phv_data_86 : _GEN_3901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3903 = 8'h57 == total_offset_7 ? phv_data_87 : _GEN_3902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3904 = 8'h58 == total_offset_7 ? phv_data_88 : _GEN_3903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3905 = 8'h59 == total_offset_7 ? phv_data_89 : _GEN_3904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3906 = 8'h5a == total_offset_7 ? phv_data_90 : _GEN_3905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3907 = 8'h5b == total_offset_7 ? phv_data_91 : _GEN_3906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3908 = 8'h5c == total_offset_7 ? phv_data_92 : _GEN_3907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3909 = 8'h5d == total_offset_7 ? phv_data_93 : _GEN_3908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3910 = 8'h5e == total_offset_7 ? phv_data_94 : _GEN_3909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3911 = 8'h5f == total_offset_7 ? phv_data_95 : _GEN_3910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3912 = 8'h60 == total_offset_7 ? phv_data_96 : _GEN_3911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3913 = 8'h61 == total_offset_7 ? phv_data_97 : _GEN_3912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3914 = 8'h62 == total_offset_7 ? phv_data_98 : _GEN_3913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3915 = 8'h63 == total_offset_7 ? phv_data_99 : _GEN_3914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3916 = 8'h64 == total_offset_7 ? phv_data_100 : _GEN_3915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3917 = 8'h65 == total_offset_7 ? phv_data_101 : _GEN_3916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3918 = 8'h66 == total_offset_7 ? phv_data_102 : _GEN_3917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3919 = 8'h67 == total_offset_7 ? phv_data_103 : _GEN_3918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3920 = 8'h68 == total_offset_7 ? phv_data_104 : _GEN_3919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3921 = 8'h69 == total_offset_7 ? phv_data_105 : _GEN_3920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3922 = 8'h6a == total_offset_7 ? phv_data_106 : _GEN_3921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3923 = 8'h6b == total_offset_7 ? phv_data_107 : _GEN_3922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3924 = 8'h6c == total_offset_7 ? phv_data_108 : _GEN_3923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3925 = 8'h6d == total_offset_7 ? phv_data_109 : _GEN_3924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3926 = 8'h6e == total_offset_7 ? phv_data_110 : _GEN_3925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3927 = 8'h6f == total_offset_7 ? phv_data_111 : _GEN_3926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3928 = 8'h70 == total_offset_7 ? phv_data_112 : _GEN_3927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3929 = 8'h71 == total_offset_7 ? phv_data_113 : _GEN_3928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3930 = 8'h72 == total_offset_7 ? phv_data_114 : _GEN_3929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3931 = 8'h73 == total_offset_7 ? phv_data_115 : _GEN_3930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3932 = 8'h74 == total_offset_7 ? phv_data_116 : _GEN_3931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3933 = 8'h75 == total_offset_7 ? phv_data_117 : _GEN_3932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3934 = 8'h76 == total_offset_7 ? phv_data_118 : _GEN_3933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3935 = 8'h77 == total_offset_7 ? phv_data_119 : _GEN_3934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3936 = 8'h78 == total_offset_7 ? phv_data_120 : _GEN_3935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3937 = 8'h79 == total_offset_7 ? phv_data_121 : _GEN_3936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3938 = 8'h7a == total_offset_7 ? phv_data_122 : _GEN_3937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3939 = 8'h7b == total_offset_7 ? phv_data_123 : _GEN_3938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3940 = 8'h7c == total_offset_7 ? phv_data_124 : _GEN_3939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3941 = 8'h7d == total_offset_7 ? phv_data_125 : _GEN_3940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3942 = 8'h7e == total_offset_7 ? phv_data_126 : _GEN_3941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3943 = 8'h7f == total_offset_7 ? phv_data_127 : _GEN_3942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3944 = 8'h80 == total_offset_7 ? phv_data_128 : _GEN_3943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3945 = 8'h81 == total_offset_7 ? phv_data_129 : _GEN_3944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3946 = 8'h82 == total_offset_7 ? phv_data_130 : _GEN_3945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3947 = 8'h83 == total_offset_7 ? phv_data_131 : _GEN_3946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3948 = 8'h84 == total_offset_7 ? phv_data_132 : _GEN_3947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3949 = 8'h85 == total_offset_7 ? phv_data_133 : _GEN_3948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3950 = 8'h86 == total_offset_7 ? phv_data_134 : _GEN_3949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3951 = 8'h87 == total_offset_7 ? phv_data_135 : _GEN_3950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3952 = 8'h88 == total_offset_7 ? phv_data_136 : _GEN_3951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3953 = 8'h89 == total_offset_7 ? phv_data_137 : _GEN_3952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3954 = 8'h8a == total_offset_7 ? phv_data_138 : _GEN_3953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3955 = 8'h8b == total_offset_7 ? phv_data_139 : _GEN_3954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3956 = 8'h8c == total_offset_7 ? phv_data_140 : _GEN_3955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3957 = 8'h8d == total_offset_7 ? phv_data_141 : _GEN_3956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3958 = 8'h8e == total_offset_7 ? phv_data_142 : _GEN_3957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3959 = 8'h8f == total_offset_7 ? phv_data_143 : _GEN_3958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3960 = 8'h90 == total_offset_7 ? phv_data_144 : _GEN_3959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3961 = 8'h91 == total_offset_7 ? phv_data_145 : _GEN_3960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3962 = 8'h92 == total_offset_7 ? phv_data_146 : _GEN_3961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3963 = 8'h93 == total_offset_7 ? phv_data_147 : _GEN_3962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3964 = 8'h94 == total_offset_7 ? phv_data_148 : _GEN_3963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3965 = 8'h95 == total_offset_7 ? phv_data_149 : _GEN_3964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3966 = 8'h96 == total_offset_7 ? phv_data_150 : _GEN_3965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3967 = 8'h97 == total_offset_7 ? phv_data_151 : _GEN_3966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3968 = 8'h98 == total_offset_7 ? phv_data_152 : _GEN_3967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3969 = 8'h99 == total_offset_7 ? phv_data_153 : _GEN_3968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3970 = 8'h9a == total_offset_7 ? phv_data_154 : _GEN_3969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3971 = 8'h9b == total_offset_7 ? phv_data_155 : _GEN_3970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3972 = 8'h9c == total_offset_7 ? phv_data_156 : _GEN_3971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3973 = 8'h9d == total_offset_7 ? phv_data_157 : _GEN_3972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3974 = 8'h9e == total_offset_7 ? phv_data_158 : _GEN_3973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3975 = 8'h9f == total_offset_7 ? phv_data_159 : _GEN_3974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3976 = 8'ha0 == total_offset_7 ? phv_data_160 : _GEN_3975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3977 = 8'ha1 == total_offset_7 ? phv_data_161 : _GEN_3976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3978 = 8'ha2 == total_offset_7 ? phv_data_162 : _GEN_3977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3979 = 8'ha3 == total_offset_7 ? phv_data_163 : _GEN_3978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3980 = 8'ha4 == total_offset_7 ? phv_data_164 : _GEN_3979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3981 = 8'ha5 == total_offset_7 ? phv_data_165 : _GEN_3980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3982 = 8'ha6 == total_offset_7 ? phv_data_166 : _GEN_3981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3983 = 8'ha7 == total_offset_7 ? phv_data_167 : _GEN_3982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3984 = 8'ha8 == total_offset_7 ? phv_data_168 : _GEN_3983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3985 = 8'ha9 == total_offset_7 ? phv_data_169 : _GEN_3984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3986 = 8'haa == total_offset_7 ? phv_data_170 : _GEN_3985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3987 = 8'hab == total_offset_7 ? phv_data_171 : _GEN_3986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3988 = 8'hac == total_offset_7 ? phv_data_172 : _GEN_3987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3989 = 8'had == total_offset_7 ? phv_data_173 : _GEN_3988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3990 = 8'hae == total_offset_7 ? phv_data_174 : _GEN_3989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3991 = 8'haf == total_offset_7 ? phv_data_175 : _GEN_3990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3992 = 8'hb0 == total_offset_7 ? phv_data_176 : _GEN_3991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3993 = 8'hb1 == total_offset_7 ? phv_data_177 : _GEN_3992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3994 = 8'hb2 == total_offset_7 ? phv_data_178 : _GEN_3993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3995 = 8'hb3 == total_offset_7 ? phv_data_179 : _GEN_3994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3996 = 8'hb4 == total_offset_7 ? phv_data_180 : _GEN_3995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3997 = 8'hb5 == total_offset_7 ? phv_data_181 : _GEN_3996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3998 = 8'hb6 == total_offset_7 ? phv_data_182 : _GEN_3997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_3999 = 8'hb7 == total_offset_7 ? phv_data_183 : _GEN_3998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4000 = 8'hb8 == total_offset_7 ? phv_data_184 : _GEN_3999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4001 = 8'hb9 == total_offset_7 ? phv_data_185 : _GEN_4000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4002 = 8'hba == total_offset_7 ? phv_data_186 : _GEN_4001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4003 = 8'hbb == total_offset_7 ? phv_data_187 : _GEN_4002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4004 = 8'hbc == total_offset_7 ? phv_data_188 : _GEN_4003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4005 = 8'hbd == total_offset_7 ? phv_data_189 : _GEN_4004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4006 = 8'hbe == total_offset_7 ? phv_data_190 : _GEN_4005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4007 = 8'hbf == total_offset_7 ? phv_data_191 : _GEN_4006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4008 = 8'hc0 == total_offset_7 ? phv_data_192 : _GEN_4007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4009 = 8'hc1 == total_offset_7 ? phv_data_193 : _GEN_4008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4010 = 8'hc2 == total_offset_7 ? phv_data_194 : _GEN_4009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4011 = 8'hc3 == total_offset_7 ? phv_data_195 : _GEN_4010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4012 = 8'hc4 == total_offset_7 ? phv_data_196 : _GEN_4011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4013 = 8'hc5 == total_offset_7 ? phv_data_197 : _GEN_4012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4014 = 8'hc6 == total_offset_7 ? phv_data_198 : _GEN_4013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4015 = 8'hc7 == total_offset_7 ? phv_data_199 : _GEN_4014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4016 = 8'hc8 == total_offset_7 ? phv_data_200 : _GEN_4015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4017 = 8'hc9 == total_offset_7 ? phv_data_201 : _GEN_4016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4018 = 8'hca == total_offset_7 ? phv_data_202 : _GEN_4017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4019 = 8'hcb == total_offset_7 ? phv_data_203 : _GEN_4018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4020 = 8'hcc == total_offset_7 ? phv_data_204 : _GEN_4019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4021 = 8'hcd == total_offset_7 ? phv_data_205 : _GEN_4020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4022 = 8'hce == total_offset_7 ? phv_data_206 : _GEN_4021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4023 = 8'hcf == total_offset_7 ? phv_data_207 : _GEN_4022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4024 = 8'hd0 == total_offset_7 ? phv_data_208 : _GEN_4023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4025 = 8'hd1 == total_offset_7 ? phv_data_209 : _GEN_4024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4026 = 8'hd2 == total_offset_7 ? phv_data_210 : _GEN_4025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4027 = 8'hd3 == total_offset_7 ? phv_data_211 : _GEN_4026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4028 = 8'hd4 == total_offset_7 ? phv_data_212 : _GEN_4027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4029 = 8'hd5 == total_offset_7 ? phv_data_213 : _GEN_4028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4030 = 8'hd6 == total_offset_7 ? phv_data_214 : _GEN_4029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4031 = 8'hd7 == total_offset_7 ? phv_data_215 : _GEN_4030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4032 = 8'hd8 == total_offset_7 ? phv_data_216 : _GEN_4031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4033 = 8'hd9 == total_offset_7 ? phv_data_217 : _GEN_4032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4034 = 8'hda == total_offset_7 ? phv_data_218 : _GEN_4033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4035 = 8'hdb == total_offset_7 ? phv_data_219 : _GEN_4034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4036 = 8'hdc == total_offset_7 ? phv_data_220 : _GEN_4035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4037 = 8'hdd == total_offset_7 ? phv_data_221 : _GEN_4036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4038 = 8'hde == total_offset_7 ? phv_data_222 : _GEN_4037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4039 = 8'hdf == total_offset_7 ? phv_data_223 : _GEN_4038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4040 = 8'he0 == total_offset_7 ? phv_data_224 : _GEN_4039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4041 = 8'he1 == total_offset_7 ? phv_data_225 : _GEN_4040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4042 = 8'he2 == total_offset_7 ? phv_data_226 : _GEN_4041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4043 = 8'he3 == total_offset_7 ? phv_data_227 : _GEN_4042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4044 = 8'he4 == total_offset_7 ? phv_data_228 : _GEN_4043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4045 = 8'he5 == total_offset_7 ? phv_data_229 : _GEN_4044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4046 = 8'he6 == total_offset_7 ? phv_data_230 : _GEN_4045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4047 = 8'he7 == total_offset_7 ? phv_data_231 : _GEN_4046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4048 = 8'he8 == total_offset_7 ? phv_data_232 : _GEN_4047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4049 = 8'he9 == total_offset_7 ? phv_data_233 : _GEN_4048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4050 = 8'hea == total_offset_7 ? phv_data_234 : _GEN_4049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4051 = 8'heb == total_offset_7 ? phv_data_235 : _GEN_4050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4052 = 8'hec == total_offset_7 ? phv_data_236 : _GEN_4051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4053 = 8'hed == total_offset_7 ? phv_data_237 : _GEN_4052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4054 = 8'hee == total_offset_7 ? phv_data_238 : _GEN_4053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4055 = 8'hef == total_offset_7 ? phv_data_239 : _GEN_4054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4056 = 8'hf0 == total_offset_7 ? phv_data_240 : _GEN_4055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4057 = 8'hf1 == total_offset_7 ? phv_data_241 : _GEN_4056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4058 = 8'hf2 == total_offset_7 ? phv_data_242 : _GEN_4057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4059 = 8'hf3 == total_offset_7 ? phv_data_243 : _GEN_4058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4060 = 8'hf4 == total_offset_7 ? phv_data_244 : _GEN_4059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4061 = 8'hf5 == total_offset_7 ? phv_data_245 : _GEN_4060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4062 = 8'hf6 == total_offset_7 ? phv_data_246 : _GEN_4061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4063 = 8'hf7 == total_offset_7 ? phv_data_247 : _GEN_4062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4064 = 8'hf8 == total_offset_7 ? phv_data_248 : _GEN_4063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4065 = 8'hf9 == total_offset_7 ? phv_data_249 : _GEN_4064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4066 = 8'hfa == total_offset_7 ? phv_data_250 : _GEN_4065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4067 = 8'hfb == total_offset_7 ? phv_data_251 : _GEN_4066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4068 = 8'hfc == total_offset_7 ? phv_data_252 : _GEN_4067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4069 = 8'hfd == total_offset_7 ? phv_data_253 : _GEN_4068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4070 = 8'hfe == total_offset_7 ? phv_data_254 : _GEN_4069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4071 = 8'hff == total_offset_7 ? phv_data_255 : _GEN_4070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_10920 = {{1'd0}, total_offset_7}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4072 = 9'h100 == _GEN_10920 ? phv_data_256 : _GEN_4071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4073 = 9'h101 == _GEN_10920 ? phv_data_257 : _GEN_4072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4074 = 9'h102 == _GEN_10920 ? phv_data_258 : _GEN_4073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4075 = 9'h103 == _GEN_10920 ? phv_data_259 : _GEN_4074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4076 = 9'h104 == _GEN_10920 ? phv_data_260 : _GEN_4075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4077 = 9'h105 == _GEN_10920 ? phv_data_261 : _GEN_4076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4078 = 9'h106 == _GEN_10920 ? phv_data_262 : _GEN_4077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4079 = 9'h107 == _GEN_10920 ? phv_data_263 : _GEN_4078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4080 = 9'h108 == _GEN_10920 ? phv_data_264 : _GEN_4079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4081 = 9'h109 == _GEN_10920 ? phv_data_265 : _GEN_4080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4082 = 9'h10a == _GEN_10920 ? phv_data_266 : _GEN_4081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4083 = 9'h10b == _GEN_10920 ? phv_data_267 : _GEN_4082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4084 = 9'h10c == _GEN_10920 ? phv_data_268 : _GEN_4083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4085 = 9'h10d == _GEN_10920 ? phv_data_269 : _GEN_4084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4086 = 9'h10e == _GEN_10920 ? phv_data_270 : _GEN_4085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4087 = 9'h10f == _GEN_10920 ? phv_data_271 : _GEN_4086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4088 = 9'h110 == _GEN_10920 ? phv_data_272 : _GEN_4087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4089 = 9'h111 == _GEN_10920 ? phv_data_273 : _GEN_4088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4090 = 9'h112 == _GEN_10920 ? phv_data_274 : _GEN_4089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4091 = 9'h113 == _GEN_10920 ? phv_data_275 : _GEN_4090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4092 = 9'h114 == _GEN_10920 ? phv_data_276 : _GEN_4091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4093 = 9'h115 == _GEN_10920 ? phv_data_277 : _GEN_4092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4094 = 9'h116 == _GEN_10920 ? phv_data_278 : _GEN_4093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4095 = 9'h117 == _GEN_10920 ? phv_data_279 : _GEN_4094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4096 = 9'h118 == _GEN_10920 ? phv_data_280 : _GEN_4095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4097 = 9'h119 == _GEN_10920 ? phv_data_281 : _GEN_4096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4098 = 9'h11a == _GEN_10920 ? phv_data_282 : _GEN_4097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4099 = 9'h11b == _GEN_10920 ? phv_data_283 : _GEN_4098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4100 = 9'h11c == _GEN_10920 ? phv_data_284 : _GEN_4099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4101 = 9'h11d == _GEN_10920 ? phv_data_285 : _GEN_4100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4102 = 9'h11e == _GEN_10920 ? phv_data_286 : _GEN_4101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4103 = 9'h11f == _GEN_10920 ? phv_data_287 : _GEN_4102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4104 = 9'h120 == _GEN_10920 ? phv_data_288 : _GEN_4103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4105 = 9'h121 == _GEN_10920 ? phv_data_289 : _GEN_4104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4106 = 9'h122 == _GEN_10920 ? phv_data_290 : _GEN_4105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4107 = 9'h123 == _GEN_10920 ? phv_data_291 : _GEN_4106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4108 = 9'h124 == _GEN_10920 ? phv_data_292 : _GEN_4107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4109 = 9'h125 == _GEN_10920 ? phv_data_293 : _GEN_4108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4110 = 9'h126 == _GEN_10920 ? phv_data_294 : _GEN_4109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4111 = 9'h127 == _GEN_10920 ? phv_data_295 : _GEN_4110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4112 = 9'h128 == _GEN_10920 ? phv_data_296 : _GEN_4111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4113 = 9'h129 == _GEN_10920 ? phv_data_297 : _GEN_4112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4114 = 9'h12a == _GEN_10920 ? phv_data_298 : _GEN_4113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4115 = 9'h12b == _GEN_10920 ? phv_data_299 : _GEN_4114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4116 = 9'h12c == _GEN_10920 ? phv_data_300 : _GEN_4115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4117 = 9'h12d == _GEN_10920 ? phv_data_301 : _GEN_4116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4118 = 9'h12e == _GEN_10920 ? phv_data_302 : _GEN_4117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4119 = 9'h12f == _GEN_10920 ? phv_data_303 : _GEN_4118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4120 = 9'h130 == _GEN_10920 ? phv_data_304 : _GEN_4119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4121 = 9'h131 == _GEN_10920 ? phv_data_305 : _GEN_4120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4122 = 9'h132 == _GEN_10920 ? phv_data_306 : _GEN_4121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4123 = 9'h133 == _GEN_10920 ? phv_data_307 : _GEN_4122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4124 = 9'h134 == _GEN_10920 ? phv_data_308 : _GEN_4123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4125 = 9'h135 == _GEN_10920 ? phv_data_309 : _GEN_4124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4126 = 9'h136 == _GEN_10920 ? phv_data_310 : _GEN_4125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4127 = 9'h137 == _GEN_10920 ? phv_data_311 : _GEN_4126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4128 = 9'h138 == _GEN_10920 ? phv_data_312 : _GEN_4127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4129 = 9'h139 == _GEN_10920 ? phv_data_313 : _GEN_4128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4130 = 9'h13a == _GEN_10920 ? phv_data_314 : _GEN_4129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4131 = 9'h13b == _GEN_10920 ? phv_data_315 : _GEN_4130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4132 = 9'h13c == _GEN_10920 ? phv_data_316 : _GEN_4131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4133 = 9'h13d == _GEN_10920 ? phv_data_317 : _GEN_4132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4134 = 9'h13e == _GEN_10920 ? phv_data_318 : _GEN_4133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4135 = 9'h13f == _GEN_10920 ? phv_data_319 : _GEN_4134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4136 = 9'h140 == _GEN_10920 ? phv_data_320 : _GEN_4135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4137 = 9'h141 == _GEN_10920 ? phv_data_321 : _GEN_4136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4138 = 9'h142 == _GEN_10920 ? phv_data_322 : _GEN_4137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4139 = 9'h143 == _GEN_10920 ? phv_data_323 : _GEN_4138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4140 = 9'h144 == _GEN_10920 ? phv_data_324 : _GEN_4139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4141 = 9'h145 == _GEN_10920 ? phv_data_325 : _GEN_4140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4142 = 9'h146 == _GEN_10920 ? phv_data_326 : _GEN_4141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4143 = 9'h147 == _GEN_10920 ? phv_data_327 : _GEN_4142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4144 = 9'h148 == _GEN_10920 ? phv_data_328 : _GEN_4143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4145 = 9'h149 == _GEN_10920 ? phv_data_329 : _GEN_4144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4146 = 9'h14a == _GEN_10920 ? phv_data_330 : _GEN_4145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4147 = 9'h14b == _GEN_10920 ? phv_data_331 : _GEN_4146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4148 = 9'h14c == _GEN_10920 ? phv_data_332 : _GEN_4147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4149 = 9'h14d == _GEN_10920 ? phv_data_333 : _GEN_4148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4150 = 9'h14e == _GEN_10920 ? phv_data_334 : _GEN_4149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4151 = 9'h14f == _GEN_10920 ? phv_data_335 : _GEN_4150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4152 = 9'h150 == _GEN_10920 ? phv_data_336 : _GEN_4151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4153 = 9'h151 == _GEN_10920 ? phv_data_337 : _GEN_4152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4154 = 9'h152 == _GEN_10920 ? phv_data_338 : _GEN_4153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4155 = 9'h153 == _GEN_10920 ? phv_data_339 : _GEN_4154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4156 = 9'h154 == _GEN_10920 ? phv_data_340 : _GEN_4155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4157 = 9'h155 == _GEN_10920 ? phv_data_341 : _GEN_4156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4158 = 9'h156 == _GEN_10920 ? phv_data_342 : _GEN_4157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4159 = 9'h157 == _GEN_10920 ? phv_data_343 : _GEN_4158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4160 = 9'h158 == _GEN_10920 ? phv_data_344 : _GEN_4159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4161 = 9'h159 == _GEN_10920 ? phv_data_345 : _GEN_4160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4162 = 9'h15a == _GEN_10920 ? phv_data_346 : _GEN_4161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4163 = 9'h15b == _GEN_10920 ? phv_data_347 : _GEN_4162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4164 = 9'h15c == _GEN_10920 ? phv_data_348 : _GEN_4163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4165 = 9'h15d == _GEN_10920 ? phv_data_349 : _GEN_4164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4166 = 9'h15e == _GEN_10920 ? phv_data_350 : _GEN_4165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4167 = 9'h15f == _GEN_10920 ? phv_data_351 : _GEN_4166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4168 = 9'h160 == _GEN_10920 ? phv_data_352 : _GEN_4167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4169 = 9'h161 == _GEN_10920 ? phv_data_353 : _GEN_4168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4170 = 9'h162 == _GEN_10920 ? phv_data_354 : _GEN_4169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4171 = 9'h163 == _GEN_10920 ? phv_data_355 : _GEN_4170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4172 = 9'h164 == _GEN_10920 ? phv_data_356 : _GEN_4171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4173 = 9'h165 == _GEN_10920 ? phv_data_357 : _GEN_4172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4174 = 9'h166 == _GEN_10920 ? phv_data_358 : _GEN_4173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4175 = 9'h167 == _GEN_10920 ? phv_data_359 : _GEN_4174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4176 = 9'h168 == _GEN_10920 ? phv_data_360 : _GEN_4175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4177 = 9'h169 == _GEN_10920 ? phv_data_361 : _GEN_4176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4178 = 9'h16a == _GEN_10920 ? phv_data_362 : _GEN_4177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4179 = 9'h16b == _GEN_10920 ? phv_data_363 : _GEN_4178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4180 = 9'h16c == _GEN_10920 ? phv_data_364 : _GEN_4179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4181 = 9'h16d == _GEN_10920 ? phv_data_365 : _GEN_4180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4182 = 9'h16e == _GEN_10920 ? phv_data_366 : _GEN_4181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4183 = 9'h16f == _GEN_10920 ? phv_data_367 : _GEN_4182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4184 = 9'h170 == _GEN_10920 ? phv_data_368 : _GEN_4183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4185 = 9'h171 == _GEN_10920 ? phv_data_369 : _GEN_4184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4186 = 9'h172 == _GEN_10920 ? phv_data_370 : _GEN_4185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4187 = 9'h173 == _GEN_10920 ? phv_data_371 : _GEN_4186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4188 = 9'h174 == _GEN_10920 ? phv_data_372 : _GEN_4187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4189 = 9'h175 == _GEN_10920 ? phv_data_373 : _GEN_4188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4190 = 9'h176 == _GEN_10920 ? phv_data_374 : _GEN_4189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4191 = 9'h177 == _GEN_10920 ? phv_data_375 : _GEN_4190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4192 = 9'h178 == _GEN_10920 ? phv_data_376 : _GEN_4191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4193 = 9'h179 == _GEN_10920 ? phv_data_377 : _GEN_4192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4194 = 9'h17a == _GEN_10920 ? phv_data_378 : _GEN_4193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4195 = 9'h17b == _GEN_10920 ? phv_data_379 : _GEN_4194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4196 = 9'h17c == _GEN_10920 ? phv_data_380 : _GEN_4195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4197 = 9'h17d == _GEN_10920 ? phv_data_381 : _GEN_4196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4198 = 9'h17e == _GEN_10920 ? phv_data_382 : _GEN_4197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4199 = 9'h17f == _GEN_10920 ? phv_data_383 : _GEN_4198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4200 = 9'h180 == _GEN_10920 ? phv_data_384 : _GEN_4199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4201 = 9'h181 == _GEN_10920 ? phv_data_385 : _GEN_4200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4202 = 9'h182 == _GEN_10920 ? phv_data_386 : _GEN_4201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4203 = 9'h183 == _GEN_10920 ? phv_data_387 : _GEN_4202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4204 = 9'h184 == _GEN_10920 ? phv_data_388 : _GEN_4203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4205 = 9'h185 == _GEN_10920 ? phv_data_389 : _GEN_4204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4206 = 9'h186 == _GEN_10920 ? phv_data_390 : _GEN_4205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4207 = 9'h187 == _GEN_10920 ? phv_data_391 : _GEN_4206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4208 = 9'h188 == _GEN_10920 ? phv_data_392 : _GEN_4207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4209 = 9'h189 == _GEN_10920 ? phv_data_393 : _GEN_4208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4210 = 9'h18a == _GEN_10920 ? phv_data_394 : _GEN_4209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4211 = 9'h18b == _GEN_10920 ? phv_data_395 : _GEN_4210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4212 = 9'h18c == _GEN_10920 ? phv_data_396 : _GEN_4211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4213 = 9'h18d == _GEN_10920 ? phv_data_397 : _GEN_4212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4214 = 9'h18e == _GEN_10920 ? phv_data_398 : _GEN_4213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4215 = 9'h18f == _GEN_10920 ? phv_data_399 : _GEN_4214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4216 = 9'h190 == _GEN_10920 ? phv_data_400 : _GEN_4215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4217 = 9'h191 == _GEN_10920 ? phv_data_401 : _GEN_4216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4218 = 9'h192 == _GEN_10920 ? phv_data_402 : _GEN_4217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4219 = 9'h193 == _GEN_10920 ? phv_data_403 : _GEN_4218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4220 = 9'h194 == _GEN_10920 ? phv_data_404 : _GEN_4219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4221 = 9'h195 == _GEN_10920 ? phv_data_405 : _GEN_4220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4222 = 9'h196 == _GEN_10920 ? phv_data_406 : _GEN_4221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4223 = 9'h197 == _GEN_10920 ? phv_data_407 : _GEN_4222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4224 = 9'h198 == _GEN_10920 ? phv_data_408 : _GEN_4223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4225 = 9'h199 == _GEN_10920 ? phv_data_409 : _GEN_4224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4226 = 9'h19a == _GEN_10920 ? phv_data_410 : _GEN_4225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4227 = 9'h19b == _GEN_10920 ? phv_data_411 : _GEN_4226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4228 = 9'h19c == _GEN_10920 ? phv_data_412 : _GEN_4227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4229 = 9'h19d == _GEN_10920 ? phv_data_413 : _GEN_4228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4230 = 9'h19e == _GEN_10920 ? phv_data_414 : _GEN_4229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4231 = 9'h19f == _GEN_10920 ? phv_data_415 : _GEN_4230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4232 = 9'h1a0 == _GEN_10920 ? phv_data_416 : _GEN_4231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4233 = 9'h1a1 == _GEN_10920 ? phv_data_417 : _GEN_4232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4234 = 9'h1a2 == _GEN_10920 ? phv_data_418 : _GEN_4233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4235 = 9'h1a3 == _GEN_10920 ? phv_data_419 : _GEN_4234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4236 = 9'h1a4 == _GEN_10920 ? phv_data_420 : _GEN_4235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4237 = 9'h1a5 == _GEN_10920 ? phv_data_421 : _GEN_4236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4238 = 9'h1a6 == _GEN_10920 ? phv_data_422 : _GEN_4237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4239 = 9'h1a7 == _GEN_10920 ? phv_data_423 : _GEN_4238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4240 = 9'h1a8 == _GEN_10920 ? phv_data_424 : _GEN_4239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4241 = 9'h1a9 == _GEN_10920 ? phv_data_425 : _GEN_4240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4242 = 9'h1aa == _GEN_10920 ? phv_data_426 : _GEN_4241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4243 = 9'h1ab == _GEN_10920 ? phv_data_427 : _GEN_4242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4244 = 9'h1ac == _GEN_10920 ? phv_data_428 : _GEN_4243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4245 = 9'h1ad == _GEN_10920 ? phv_data_429 : _GEN_4244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4246 = 9'h1ae == _GEN_10920 ? phv_data_430 : _GEN_4245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4247 = 9'h1af == _GEN_10920 ? phv_data_431 : _GEN_4246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4248 = 9'h1b0 == _GEN_10920 ? phv_data_432 : _GEN_4247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4249 = 9'h1b1 == _GEN_10920 ? phv_data_433 : _GEN_4248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4250 = 9'h1b2 == _GEN_10920 ? phv_data_434 : _GEN_4249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4251 = 9'h1b3 == _GEN_10920 ? phv_data_435 : _GEN_4250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4252 = 9'h1b4 == _GEN_10920 ? phv_data_436 : _GEN_4251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4253 = 9'h1b5 == _GEN_10920 ? phv_data_437 : _GEN_4252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4254 = 9'h1b6 == _GEN_10920 ? phv_data_438 : _GEN_4253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4255 = 9'h1b7 == _GEN_10920 ? phv_data_439 : _GEN_4254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4256 = 9'h1b8 == _GEN_10920 ? phv_data_440 : _GEN_4255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4257 = 9'h1b9 == _GEN_10920 ? phv_data_441 : _GEN_4256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4258 = 9'h1ba == _GEN_10920 ? phv_data_442 : _GEN_4257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4259 = 9'h1bb == _GEN_10920 ? phv_data_443 : _GEN_4258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4260 = 9'h1bc == _GEN_10920 ? phv_data_444 : _GEN_4259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4261 = 9'h1bd == _GEN_10920 ? phv_data_445 : _GEN_4260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4262 = 9'h1be == _GEN_10920 ? phv_data_446 : _GEN_4261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4263 = 9'h1bf == _GEN_10920 ? phv_data_447 : _GEN_4262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4264 = 9'h1c0 == _GEN_10920 ? phv_data_448 : _GEN_4263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4265 = 9'h1c1 == _GEN_10920 ? phv_data_449 : _GEN_4264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4266 = 9'h1c2 == _GEN_10920 ? phv_data_450 : _GEN_4265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4267 = 9'h1c3 == _GEN_10920 ? phv_data_451 : _GEN_4266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4268 = 9'h1c4 == _GEN_10920 ? phv_data_452 : _GEN_4267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4269 = 9'h1c5 == _GEN_10920 ? phv_data_453 : _GEN_4268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4270 = 9'h1c6 == _GEN_10920 ? phv_data_454 : _GEN_4269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4271 = 9'h1c7 == _GEN_10920 ? phv_data_455 : _GEN_4270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4272 = 9'h1c8 == _GEN_10920 ? phv_data_456 : _GEN_4271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4273 = 9'h1c9 == _GEN_10920 ? phv_data_457 : _GEN_4272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4274 = 9'h1ca == _GEN_10920 ? phv_data_458 : _GEN_4273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4275 = 9'h1cb == _GEN_10920 ? phv_data_459 : _GEN_4274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4276 = 9'h1cc == _GEN_10920 ? phv_data_460 : _GEN_4275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4277 = 9'h1cd == _GEN_10920 ? phv_data_461 : _GEN_4276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4278 = 9'h1ce == _GEN_10920 ? phv_data_462 : _GEN_4277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4279 = 9'h1cf == _GEN_10920 ? phv_data_463 : _GEN_4278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4280 = 9'h1d0 == _GEN_10920 ? phv_data_464 : _GEN_4279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4281 = 9'h1d1 == _GEN_10920 ? phv_data_465 : _GEN_4280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4282 = 9'h1d2 == _GEN_10920 ? phv_data_466 : _GEN_4281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4283 = 9'h1d3 == _GEN_10920 ? phv_data_467 : _GEN_4282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4284 = 9'h1d4 == _GEN_10920 ? phv_data_468 : _GEN_4283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4285 = 9'h1d5 == _GEN_10920 ? phv_data_469 : _GEN_4284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4286 = 9'h1d6 == _GEN_10920 ? phv_data_470 : _GEN_4285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4287 = 9'h1d7 == _GEN_10920 ? phv_data_471 : _GEN_4286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4288 = 9'h1d8 == _GEN_10920 ? phv_data_472 : _GEN_4287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4289 = 9'h1d9 == _GEN_10920 ? phv_data_473 : _GEN_4288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4290 = 9'h1da == _GEN_10920 ? phv_data_474 : _GEN_4289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4291 = 9'h1db == _GEN_10920 ? phv_data_475 : _GEN_4290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4292 = 9'h1dc == _GEN_10920 ? phv_data_476 : _GEN_4291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4293 = 9'h1dd == _GEN_10920 ? phv_data_477 : _GEN_4292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4294 = 9'h1de == _GEN_10920 ? phv_data_478 : _GEN_4293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4295 = 9'h1df == _GEN_10920 ? phv_data_479 : _GEN_4294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4296 = 9'h1e0 == _GEN_10920 ? phv_data_480 : _GEN_4295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4297 = 9'h1e1 == _GEN_10920 ? phv_data_481 : _GEN_4296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4298 = 9'h1e2 == _GEN_10920 ? phv_data_482 : _GEN_4297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4299 = 9'h1e3 == _GEN_10920 ? phv_data_483 : _GEN_4298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4300 = 9'h1e4 == _GEN_10920 ? phv_data_484 : _GEN_4299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4301 = 9'h1e5 == _GEN_10920 ? phv_data_485 : _GEN_4300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4302 = 9'h1e6 == _GEN_10920 ? phv_data_486 : _GEN_4301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4303 = 9'h1e7 == _GEN_10920 ? phv_data_487 : _GEN_4302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4304 = 9'h1e8 == _GEN_10920 ? phv_data_488 : _GEN_4303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4305 = 9'h1e9 == _GEN_10920 ? phv_data_489 : _GEN_4304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4306 = 9'h1ea == _GEN_10920 ? phv_data_490 : _GEN_4305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4307 = 9'h1eb == _GEN_10920 ? phv_data_491 : _GEN_4306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4308 = 9'h1ec == _GEN_10920 ? phv_data_492 : _GEN_4307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4309 = 9'h1ed == _GEN_10920 ? phv_data_493 : _GEN_4308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4310 = 9'h1ee == _GEN_10920 ? phv_data_494 : _GEN_4309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4311 = 9'h1ef == _GEN_10920 ? phv_data_495 : _GEN_4310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4312 = 9'h1f0 == _GEN_10920 ? phv_data_496 : _GEN_4311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4313 = 9'h1f1 == _GEN_10920 ? phv_data_497 : _GEN_4312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4314 = 9'h1f2 == _GEN_10920 ? phv_data_498 : _GEN_4313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4315 = 9'h1f3 == _GEN_10920 ? phv_data_499 : _GEN_4314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4316 = 9'h1f4 == _GEN_10920 ? phv_data_500 : _GEN_4315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4317 = 9'h1f5 == _GEN_10920 ? phv_data_501 : _GEN_4316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4318 = 9'h1f6 == _GEN_10920 ? phv_data_502 : _GEN_4317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4319 = 9'h1f7 == _GEN_10920 ? phv_data_503 : _GEN_4318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4320 = 9'h1f8 == _GEN_10920 ? phv_data_504 : _GEN_4319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4321 = 9'h1f9 == _GEN_10920 ? phv_data_505 : _GEN_4320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4322 = 9'h1fa == _GEN_10920 ? phv_data_506 : _GEN_4321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4323 = 9'h1fb == _GEN_10920 ? phv_data_507 : _GEN_4322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4324 = 9'h1fc == _GEN_10920 ? phv_data_508 : _GEN_4323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4325 = 9'h1fd == _GEN_10920 ? phv_data_509 : _GEN_4324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4326 = 9'h1fe == _GEN_10920 ? phv_data_510 : _GEN_4325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_1_0 = 9'h1ff == _GEN_10920 ? phv_data_511 : _GEN_4326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_1_T = {bytes_1_0,bytes_1_1,bytes_1_2,bytes_1_3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_1_T = {_mask_3_T_10,mask_1_1,mask_1_2,mask_1_3}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_1 = io_field_out_1_lo[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_1 = io_field_out_1_lo[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _local_offset_T_57 = {{1'd0}, args_offset_1}; // @[executor.scala 222:61]
  wire [2:0] local_offset_28 = _local_offset_T_57[2:0]; // @[executor.scala 222:61]
  wire [7:0] _GEN_4329 = 3'h1 == local_offset_28 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4330 = 3'h2 == local_offset_28 ? args_2 : _GEN_4329; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4331 = 3'h3 == local_offset_28 ? args_3 : _GEN_4330; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4332 = 3'h4 == local_offset_28 ? args_4 : _GEN_4331; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4333 = 3'h5 == local_offset_28 ? args_5 : _GEN_4332; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4334 = 3'h6 == local_offset_28 ? args_6 : _GEN_4333; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4335 = 3'h1 == args_length_1 ? _GEN_4334 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [2:0] local_offset_29 = 3'h1 + args_offset_1; // @[executor.scala 222:61]
  wire [7:0] _GEN_4337 = 3'h1 == local_offset_29 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4338 = 3'h2 == local_offset_29 ? args_2 : _GEN_4337; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4339 = 3'h3 == local_offset_29 ? args_3 : _GEN_4338; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4340 = 3'h4 == local_offset_29 ? args_4 : _GEN_4339; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4341 = 3'h5 == local_offset_29 ? args_5 : _GEN_4340; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4342 = 3'h6 == local_offset_29 ? args_6 : _GEN_4341; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4343 = 3'h2 == args_length_1 ? _GEN_4342 : _GEN_4335; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_30 = 3'h2 + args_offset_1; // @[executor.scala 222:61]
  wire [7:0] _GEN_4345 = 3'h1 == local_offset_30 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4346 = 3'h2 == local_offset_30 ? args_2 : _GEN_4345; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4347 = 3'h3 == local_offset_30 ? args_3 : _GEN_4346; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4348 = 3'h4 == local_offset_30 ? args_4 : _GEN_4347; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4349 = 3'h5 == local_offset_30 ? args_5 : _GEN_4348; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4350 = 3'h6 == local_offset_30 ? args_6 : _GEN_4349; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4351 = 3'h3 == args_length_1 ? _GEN_4350 : _GEN_4343; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_31 = 3'h3 + args_offset_1; // @[executor.scala 222:61]
  wire [7:0] _GEN_4353 = 3'h1 == local_offset_31 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4354 = 3'h2 == local_offset_31 ? args_2 : _GEN_4353; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4355 = 3'h3 == local_offset_31 ? args_3 : _GEN_4354; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4356 = 3'h4 == local_offset_31 ? args_4 : _GEN_4355; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4357 = 3'h5 == local_offset_31 ? args_5 : _GEN_4356; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4358 = 3'h6 == local_offset_31 ? args_6 : _GEN_4357; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4359 = 3'h4 == args_length_1 ? _GEN_4358 : _GEN_4351; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_32 = 3'h4 + args_offset_1; // @[executor.scala 222:61]
  wire [7:0] _GEN_4361 = 3'h1 == local_offset_32 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4362 = 3'h2 == local_offset_32 ? args_2 : _GEN_4361; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4363 = 3'h3 == local_offset_32 ? args_3 : _GEN_4362; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4364 = 3'h4 == local_offset_32 ? args_4 : _GEN_4363; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4365 = 3'h5 == local_offset_32 ? args_5 : _GEN_4364; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4366 = 3'h6 == local_offset_32 ? args_6 : _GEN_4365; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4367 = 3'h5 == args_length_1 ? _GEN_4366 : _GEN_4359; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_33 = 3'h5 + args_offset_1; // @[executor.scala 222:61]
  wire [7:0] _GEN_4369 = 3'h1 == local_offset_33 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4370 = 3'h2 == local_offset_33 ? args_2 : _GEN_4369; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4371 = 3'h3 == local_offset_33 ? args_3 : _GEN_4370; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4372 = 3'h4 == local_offset_33 ? args_4 : _GEN_4371; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4373 = 3'h5 == local_offset_33 ? args_5 : _GEN_4372; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4374 = 3'h6 == local_offset_33 ? args_6 : _GEN_4373; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4375 = 3'h6 == args_length_1 ? _GEN_4374 : _GEN_4367; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_34 = 3'h6 + args_offset_1; // @[executor.scala 222:61]
  wire [7:0] _GEN_4377 = 3'h1 == local_offset_34 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4378 = 3'h2 == local_offset_34 ? args_2 : _GEN_4377; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4379 = 3'h3 == local_offset_34 ? args_3 : _GEN_4378; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4380 = 3'h4 == local_offset_34 ? args_4 : _GEN_4379; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4381 = 3'h5 == local_offset_34 ? args_5 : _GEN_4380; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_4382 = 3'h6 == local_offset_34 ? args_6 : _GEN_4381; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] field_bytes_3_0 = 3'h7 == args_length_1 ? _GEN_4382 : _GEN_4375; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4391 = 3'h2 == args_length_1 ? _GEN_4334 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_4399 = 3'h3 == args_length_1 ? _GEN_4342 : _GEN_4391; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4407 = 3'h4 == args_length_1 ? _GEN_4350 : _GEN_4399; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4415 = 3'h5 == args_length_1 ? _GEN_4358 : _GEN_4407; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4423 = 3'h6 == args_length_1 ? _GEN_4366 : _GEN_4415; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4431 = 3'h7 == args_length_1 ? _GEN_4374 : _GEN_4423; // @[executor.scala 223:66 executor.scala 224:52]
  wire [3:0] _GEN_11176 = {{1'd0}, args_length_1}; // @[executor.scala 223:49]
  wire [7:0] field_bytes_3_1 = 4'h8 == _GEN_11176 ? _GEN_4382 : _GEN_4431; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4447 = 3'h3 == args_length_1 ? _GEN_4334 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_4455 = 3'h4 == args_length_1 ? _GEN_4342 : _GEN_4447; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4463 = 3'h5 == args_length_1 ? _GEN_4350 : _GEN_4455; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4471 = 3'h6 == args_length_1 ? _GEN_4358 : _GEN_4463; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4479 = 3'h7 == args_length_1 ? _GEN_4366 : _GEN_4471; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4487 = 4'h8 == _GEN_11176 ? _GEN_4374 : _GEN_4479; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_3_2 = 4'h9 == _GEN_11176 ? _GEN_4382 : _GEN_4487; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4503 = 3'h4 == args_length_1 ? _GEN_4334 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_4511 = 3'h5 == args_length_1 ? _GEN_4342 : _GEN_4503; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4519 = 3'h6 == args_length_1 ? _GEN_4350 : _GEN_4511; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4527 = 3'h7 == args_length_1 ? _GEN_4358 : _GEN_4519; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4535 = 4'h8 == _GEN_11176 ? _GEN_4366 : _GEN_4527; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_4543 = 4'h9 == _GEN_11176 ? _GEN_4374 : _GEN_4535; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_3_3 = 4'ha == _GEN_11176 ? _GEN_4382 : _GEN_4543; // @[executor.scala 223:66 executor.scala 224:52]
  wire [31:0] _io_field_out_1_T_1 = {field_bytes_3_0,field_bytes_3_1,field_bytes_3_2,field_bytes_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_4552 = 4'ha == opcode_1 ? _io_field_out_1_T_1 : 32'h0; // @[executor.scala 207:55 executor.scala 228:41 executor.scala 172:29]
  wire [17:0] io_field_out_1_hi_4 = io_field_out_1_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_1_T_4 = {io_field_out_1_hi_4,io_field_out_1_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_4553 = 4'hb == opcode_1 ? _io_field_out_1_T_4 : _GEN_4552; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_4554 = from_header_1 ? bias_1 : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_4555 = from_header_1 ? _io_field_out_1_T : _GEN_4553; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_4556 = from_header_1 ? _io_mask_out_1_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  wire [3:0] opcode_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_2_lo = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire  from_header_2 = length_2 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi_2 = offset_2[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_5 = offset_2 + length_2; // @[executor.scala 193:46]
  wire [1:0] ending_2 = _ending_T_5[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_11182 = {{2'd0}, ending_2}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_5 = 4'h4 - _GEN_11182; // @[executor.scala 194:45]
  wire [1:0] bias_2 = _bias_T_5[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset_8 = {total_offset_hi_2,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_4561 = 8'h1 == total_offset_8 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4562 = 8'h2 == total_offset_8 ? phv_data_2 : _GEN_4561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4563 = 8'h3 == total_offset_8 ? phv_data_3 : _GEN_4562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4564 = 8'h4 == total_offset_8 ? phv_data_4 : _GEN_4563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4565 = 8'h5 == total_offset_8 ? phv_data_5 : _GEN_4564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4566 = 8'h6 == total_offset_8 ? phv_data_6 : _GEN_4565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4567 = 8'h7 == total_offset_8 ? phv_data_7 : _GEN_4566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4568 = 8'h8 == total_offset_8 ? phv_data_8 : _GEN_4567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4569 = 8'h9 == total_offset_8 ? phv_data_9 : _GEN_4568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4570 = 8'ha == total_offset_8 ? phv_data_10 : _GEN_4569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4571 = 8'hb == total_offset_8 ? phv_data_11 : _GEN_4570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4572 = 8'hc == total_offset_8 ? phv_data_12 : _GEN_4571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4573 = 8'hd == total_offset_8 ? phv_data_13 : _GEN_4572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4574 = 8'he == total_offset_8 ? phv_data_14 : _GEN_4573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4575 = 8'hf == total_offset_8 ? phv_data_15 : _GEN_4574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4576 = 8'h10 == total_offset_8 ? phv_data_16 : _GEN_4575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4577 = 8'h11 == total_offset_8 ? phv_data_17 : _GEN_4576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4578 = 8'h12 == total_offset_8 ? phv_data_18 : _GEN_4577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4579 = 8'h13 == total_offset_8 ? phv_data_19 : _GEN_4578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4580 = 8'h14 == total_offset_8 ? phv_data_20 : _GEN_4579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4581 = 8'h15 == total_offset_8 ? phv_data_21 : _GEN_4580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4582 = 8'h16 == total_offset_8 ? phv_data_22 : _GEN_4581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4583 = 8'h17 == total_offset_8 ? phv_data_23 : _GEN_4582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4584 = 8'h18 == total_offset_8 ? phv_data_24 : _GEN_4583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4585 = 8'h19 == total_offset_8 ? phv_data_25 : _GEN_4584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4586 = 8'h1a == total_offset_8 ? phv_data_26 : _GEN_4585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4587 = 8'h1b == total_offset_8 ? phv_data_27 : _GEN_4586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4588 = 8'h1c == total_offset_8 ? phv_data_28 : _GEN_4587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4589 = 8'h1d == total_offset_8 ? phv_data_29 : _GEN_4588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4590 = 8'h1e == total_offset_8 ? phv_data_30 : _GEN_4589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4591 = 8'h1f == total_offset_8 ? phv_data_31 : _GEN_4590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4592 = 8'h20 == total_offset_8 ? phv_data_32 : _GEN_4591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4593 = 8'h21 == total_offset_8 ? phv_data_33 : _GEN_4592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4594 = 8'h22 == total_offset_8 ? phv_data_34 : _GEN_4593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4595 = 8'h23 == total_offset_8 ? phv_data_35 : _GEN_4594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4596 = 8'h24 == total_offset_8 ? phv_data_36 : _GEN_4595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4597 = 8'h25 == total_offset_8 ? phv_data_37 : _GEN_4596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4598 = 8'h26 == total_offset_8 ? phv_data_38 : _GEN_4597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4599 = 8'h27 == total_offset_8 ? phv_data_39 : _GEN_4598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4600 = 8'h28 == total_offset_8 ? phv_data_40 : _GEN_4599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4601 = 8'h29 == total_offset_8 ? phv_data_41 : _GEN_4600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4602 = 8'h2a == total_offset_8 ? phv_data_42 : _GEN_4601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4603 = 8'h2b == total_offset_8 ? phv_data_43 : _GEN_4602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4604 = 8'h2c == total_offset_8 ? phv_data_44 : _GEN_4603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4605 = 8'h2d == total_offset_8 ? phv_data_45 : _GEN_4604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4606 = 8'h2e == total_offset_8 ? phv_data_46 : _GEN_4605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4607 = 8'h2f == total_offset_8 ? phv_data_47 : _GEN_4606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4608 = 8'h30 == total_offset_8 ? phv_data_48 : _GEN_4607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4609 = 8'h31 == total_offset_8 ? phv_data_49 : _GEN_4608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4610 = 8'h32 == total_offset_8 ? phv_data_50 : _GEN_4609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4611 = 8'h33 == total_offset_8 ? phv_data_51 : _GEN_4610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4612 = 8'h34 == total_offset_8 ? phv_data_52 : _GEN_4611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4613 = 8'h35 == total_offset_8 ? phv_data_53 : _GEN_4612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4614 = 8'h36 == total_offset_8 ? phv_data_54 : _GEN_4613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4615 = 8'h37 == total_offset_8 ? phv_data_55 : _GEN_4614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4616 = 8'h38 == total_offset_8 ? phv_data_56 : _GEN_4615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4617 = 8'h39 == total_offset_8 ? phv_data_57 : _GEN_4616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4618 = 8'h3a == total_offset_8 ? phv_data_58 : _GEN_4617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4619 = 8'h3b == total_offset_8 ? phv_data_59 : _GEN_4618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4620 = 8'h3c == total_offset_8 ? phv_data_60 : _GEN_4619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4621 = 8'h3d == total_offset_8 ? phv_data_61 : _GEN_4620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4622 = 8'h3e == total_offset_8 ? phv_data_62 : _GEN_4621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4623 = 8'h3f == total_offset_8 ? phv_data_63 : _GEN_4622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4624 = 8'h40 == total_offset_8 ? phv_data_64 : _GEN_4623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4625 = 8'h41 == total_offset_8 ? phv_data_65 : _GEN_4624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4626 = 8'h42 == total_offset_8 ? phv_data_66 : _GEN_4625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4627 = 8'h43 == total_offset_8 ? phv_data_67 : _GEN_4626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4628 = 8'h44 == total_offset_8 ? phv_data_68 : _GEN_4627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4629 = 8'h45 == total_offset_8 ? phv_data_69 : _GEN_4628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4630 = 8'h46 == total_offset_8 ? phv_data_70 : _GEN_4629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4631 = 8'h47 == total_offset_8 ? phv_data_71 : _GEN_4630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4632 = 8'h48 == total_offset_8 ? phv_data_72 : _GEN_4631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4633 = 8'h49 == total_offset_8 ? phv_data_73 : _GEN_4632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4634 = 8'h4a == total_offset_8 ? phv_data_74 : _GEN_4633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4635 = 8'h4b == total_offset_8 ? phv_data_75 : _GEN_4634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4636 = 8'h4c == total_offset_8 ? phv_data_76 : _GEN_4635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4637 = 8'h4d == total_offset_8 ? phv_data_77 : _GEN_4636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4638 = 8'h4e == total_offset_8 ? phv_data_78 : _GEN_4637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4639 = 8'h4f == total_offset_8 ? phv_data_79 : _GEN_4638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4640 = 8'h50 == total_offset_8 ? phv_data_80 : _GEN_4639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4641 = 8'h51 == total_offset_8 ? phv_data_81 : _GEN_4640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4642 = 8'h52 == total_offset_8 ? phv_data_82 : _GEN_4641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4643 = 8'h53 == total_offset_8 ? phv_data_83 : _GEN_4642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4644 = 8'h54 == total_offset_8 ? phv_data_84 : _GEN_4643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4645 = 8'h55 == total_offset_8 ? phv_data_85 : _GEN_4644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4646 = 8'h56 == total_offset_8 ? phv_data_86 : _GEN_4645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4647 = 8'h57 == total_offset_8 ? phv_data_87 : _GEN_4646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4648 = 8'h58 == total_offset_8 ? phv_data_88 : _GEN_4647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4649 = 8'h59 == total_offset_8 ? phv_data_89 : _GEN_4648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4650 = 8'h5a == total_offset_8 ? phv_data_90 : _GEN_4649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4651 = 8'h5b == total_offset_8 ? phv_data_91 : _GEN_4650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4652 = 8'h5c == total_offset_8 ? phv_data_92 : _GEN_4651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4653 = 8'h5d == total_offset_8 ? phv_data_93 : _GEN_4652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4654 = 8'h5e == total_offset_8 ? phv_data_94 : _GEN_4653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4655 = 8'h5f == total_offset_8 ? phv_data_95 : _GEN_4654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4656 = 8'h60 == total_offset_8 ? phv_data_96 : _GEN_4655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4657 = 8'h61 == total_offset_8 ? phv_data_97 : _GEN_4656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4658 = 8'h62 == total_offset_8 ? phv_data_98 : _GEN_4657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4659 = 8'h63 == total_offset_8 ? phv_data_99 : _GEN_4658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4660 = 8'h64 == total_offset_8 ? phv_data_100 : _GEN_4659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4661 = 8'h65 == total_offset_8 ? phv_data_101 : _GEN_4660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4662 = 8'h66 == total_offset_8 ? phv_data_102 : _GEN_4661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4663 = 8'h67 == total_offset_8 ? phv_data_103 : _GEN_4662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4664 = 8'h68 == total_offset_8 ? phv_data_104 : _GEN_4663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4665 = 8'h69 == total_offset_8 ? phv_data_105 : _GEN_4664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4666 = 8'h6a == total_offset_8 ? phv_data_106 : _GEN_4665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4667 = 8'h6b == total_offset_8 ? phv_data_107 : _GEN_4666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4668 = 8'h6c == total_offset_8 ? phv_data_108 : _GEN_4667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4669 = 8'h6d == total_offset_8 ? phv_data_109 : _GEN_4668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4670 = 8'h6e == total_offset_8 ? phv_data_110 : _GEN_4669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4671 = 8'h6f == total_offset_8 ? phv_data_111 : _GEN_4670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4672 = 8'h70 == total_offset_8 ? phv_data_112 : _GEN_4671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4673 = 8'h71 == total_offset_8 ? phv_data_113 : _GEN_4672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4674 = 8'h72 == total_offset_8 ? phv_data_114 : _GEN_4673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4675 = 8'h73 == total_offset_8 ? phv_data_115 : _GEN_4674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4676 = 8'h74 == total_offset_8 ? phv_data_116 : _GEN_4675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4677 = 8'h75 == total_offset_8 ? phv_data_117 : _GEN_4676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4678 = 8'h76 == total_offset_8 ? phv_data_118 : _GEN_4677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4679 = 8'h77 == total_offset_8 ? phv_data_119 : _GEN_4678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4680 = 8'h78 == total_offset_8 ? phv_data_120 : _GEN_4679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4681 = 8'h79 == total_offset_8 ? phv_data_121 : _GEN_4680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4682 = 8'h7a == total_offset_8 ? phv_data_122 : _GEN_4681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4683 = 8'h7b == total_offset_8 ? phv_data_123 : _GEN_4682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4684 = 8'h7c == total_offset_8 ? phv_data_124 : _GEN_4683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4685 = 8'h7d == total_offset_8 ? phv_data_125 : _GEN_4684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4686 = 8'h7e == total_offset_8 ? phv_data_126 : _GEN_4685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4687 = 8'h7f == total_offset_8 ? phv_data_127 : _GEN_4686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4688 = 8'h80 == total_offset_8 ? phv_data_128 : _GEN_4687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4689 = 8'h81 == total_offset_8 ? phv_data_129 : _GEN_4688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4690 = 8'h82 == total_offset_8 ? phv_data_130 : _GEN_4689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4691 = 8'h83 == total_offset_8 ? phv_data_131 : _GEN_4690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4692 = 8'h84 == total_offset_8 ? phv_data_132 : _GEN_4691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4693 = 8'h85 == total_offset_8 ? phv_data_133 : _GEN_4692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4694 = 8'h86 == total_offset_8 ? phv_data_134 : _GEN_4693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4695 = 8'h87 == total_offset_8 ? phv_data_135 : _GEN_4694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4696 = 8'h88 == total_offset_8 ? phv_data_136 : _GEN_4695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4697 = 8'h89 == total_offset_8 ? phv_data_137 : _GEN_4696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4698 = 8'h8a == total_offset_8 ? phv_data_138 : _GEN_4697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4699 = 8'h8b == total_offset_8 ? phv_data_139 : _GEN_4698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4700 = 8'h8c == total_offset_8 ? phv_data_140 : _GEN_4699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4701 = 8'h8d == total_offset_8 ? phv_data_141 : _GEN_4700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4702 = 8'h8e == total_offset_8 ? phv_data_142 : _GEN_4701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4703 = 8'h8f == total_offset_8 ? phv_data_143 : _GEN_4702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4704 = 8'h90 == total_offset_8 ? phv_data_144 : _GEN_4703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4705 = 8'h91 == total_offset_8 ? phv_data_145 : _GEN_4704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4706 = 8'h92 == total_offset_8 ? phv_data_146 : _GEN_4705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4707 = 8'h93 == total_offset_8 ? phv_data_147 : _GEN_4706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4708 = 8'h94 == total_offset_8 ? phv_data_148 : _GEN_4707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4709 = 8'h95 == total_offset_8 ? phv_data_149 : _GEN_4708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4710 = 8'h96 == total_offset_8 ? phv_data_150 : _GEN_4709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4711 = 8'h97 == total_offset_8 ? phv_data_151 : _GEN_4710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4712 = 8'h98 == total_offset_8 ? phv_data_152 : _GEN_4711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4713 = 8'h99 == total_offset_8 ? phv_data_153 : _GEN_4712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4714 = 8'h9a == total_offset_8 ? phv_data_154 : _GEN_4713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4715 = 8'h9b == total_offset_8 ? phv_data_155 : _GEN_4714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4716 = 8'h9c == total_offset_8 ? phv_data_156 : _GEN_4715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4717 = 8'h9d == total_offset_8 ? phv_data_157 : _GEN_4716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4718 = 8'h9e == total_offset_8 ? phv_data_158 : _GEN_4717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4719 = 8'h9f == total_offset_8 ? phv_data_159 : _GEN_4718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4720 = 8'ha0 == total_offset_8 ? phv_data_160 : _GEN_4719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4721 = 8'ha1 == total_offset_8 ? phv_data_161 : _GEN_4720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4722 = 8'ha2 == total_offset_8 ? phv_data_162 : _GEN_4721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4723 = 8'ha3 == total_offset_8 ? phv_data_163 : _GEN_4722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4724 = 8'ha4 == total_offset_8 ? phv_data_164 : _GEN_4723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4725 = 8'ha5 == total_offset_8 ? phv_data_165 : _GEN_4724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4726 = 8'ha6 == total_offset_8 ? phv_data_166 : _GEN_4725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4727 = 8'ha7 == total_offset_8 ? phv_data_167 : _GEN_4726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4728 = 8'ha8 == total_offset_8 ? phv_data_168 : _GEN_4727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4729 = 8'ha9 == total_offset_8 ? phv_data_169 : _GEN_4728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4730 = 8'haa == total_offset_8 ? phv_data_170 : _GEN_4729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4731 = 8'hab == total_offset_8 ? phv_data_171 : _GEN_4730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4732 = 8'hac == total_offset_8 ? phv_data_172 : _GEN_4731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4733 = 8'had == total_offset_8 ? phv_data_173 : _GEN_4732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4734 = 8'hae == total_offset_8 ? phv_data_174 : _GEN_4733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4735 = 8'haf == total_offset_8 ? phv_data_175 : _GEN_4734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4736 = 8'hb0 == total_offset_8 ? phv_data_176 : _GEN_4735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4737 = 8'hb1 == total_offset_8 ? phv_data_177 : _GEN_4736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4738 = 8'hb2 == total_offset_8 ? phv_data_178 : _GEN_4737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4739 = 8'hb3 == total_offset_8 ? phv_data_179 : _GEN_4738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4740 = 8'hb4 == total_offset_8 ? phv_data_180 : _GEN_4739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4741 = 8'hb5 == total_offset_8 ? phv_data_181 : _GEN_4740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4742 = 8'hb6 == total_offset_8 ? phv_data_182 : _GEN_4741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4743 = 8'hb7 == total_offset_8 ? phv_data_183 : _GEN_4742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4744 = 8'hb8 == total_offset_8 ? phv_data_184 : _GEN_4743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4745 = 8'hb9 == total_offset_8 ? phv_data_185 : _GEN_4744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4746 = 8'hba == total_offset_8 ? phv_data_186 : _GEN_4745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4747 = 8'hbb == total_offset_8 ? phv_data_187 : _GEN_4746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4748 = 8'hbc == total_offset_8 ? phv_data_188 : _GEN_4747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4749 = 8'hbd == total_offset_8 ? phv_data_189 : _GEN_4748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4750 = 8'hbe == total_offset_8 ? phv_data_190 : _GEN_4749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4751 = 8'hbf == total_offset_8 ? phv_data_191 : _GEN_4750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4752 = 8'hc0 == total_offset_8 ? phv_data_192 : _GEN_4751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4753 = 8'hc1 == total_offset_8 ? phv_data_193 : _GEN_4752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4754 = 8'hc2 == total_offset_8 ? phv_data_194 : _GEN_4753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4755 = 8'hc3 == total_offset_8 ? phv_data_195 : _GEN_4754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4756 = 8'hc4 == total_offset_8 ? phv_data_196 : _GEN_4755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4757 = 8'hc5 == total_offset_8 ? phv_data_197 : _GEN_4756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4758 = 8'hc6 == total_offset_8 ? phv_data_198 : _GEN_4757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4759 = 8'hc7 == total_offset_8 ? phv_data_199 : _GEN_4758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4760 = 8'hc8 == total_offset_8 ? phv_data_200 : _GEN_4759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4761 = 8'hc9 == total_offset_8 ? phv_data_201 : _GEN_4760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4762 = 8'hca == total_offset_8 ? phv_data_202 : _GEN_4761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4763 = 8'hcb == total_offset_8 ? phv_data_203 : _GEN_4762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4764 = 8'hcc == total_offset_8 ? phv_data_204 : _GEN_4763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4765 = 8'hcd == total_offset_8 ? phv_data_205 : _GEN_4764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4766 = 8'hce == total_offset_8 ? phv_data_206 : _GEN_4765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4767 = 8'hcf == total_offset_8 ? phv_data_207 : _GEN_4766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4768 = 8'hd0 == total_offset_8 ? phv_data_208 : _GEN_4767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4769 = 8'hd1 == total_offset_8 ? phv_data_209 : _GEN_4768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4770 = 8'hd2 == total_offset_8 ? phv_data_210 : _GEN_4769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4771 = 8'hd3 == total_offset_8 ? phv_data_211 : _GEN_4770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4772 = 8'hd4 == total_offset_8 ? phv_data_212 : _GEN_4771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4773 = 8'hd5 == total_offset_8 ? phv_data_213 : _GEN_4772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4774 = 8'hd6 == total_offset_8 ? phv_data_214 : _GEN_4773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4775 = 8'hd7 == total_offset_8 ? phv_data_215 : _GEN_4774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4776 = 8'hd8 == total_offset_8 ? phv_data_216 : _GEN_4775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4777 = 8'hd9 == total_offset_8 ? phv_data_217 : _GEN_4776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4778 = 8'hda == total_offset_8 ? phv_data_218 : _GEN_4777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4779 = 8'hdb == total_offset_8 ? phv_data_219 : _GEN_4778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4780 = 8'hdc == total_offset_8 ? phv_data_220 : _GEN_4779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4781 = 8'hdd == total_offset_8 ? phv_data_221 : _GEN_4780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4782 = 8'hde == total_offset_8 ? phv_data_222 : _GEN_4781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4783 = 8'hdf == total_offset_8 ? phv_data_223 : _GEN_4782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4784 = 8'he0 == total_offset_8 ? phv_data_224 : _GEN_4783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4785 = 8'he1 == total_offset_8 ? phv_data_225 : _GEN_4784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4786 = 8'he2 == total_offset_8 ? phv_data_226 : _GEN_4785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4787 = 8'he3 == total_offset_8 ? phv_data_227 : _GEN_4786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4788 = 8'he4 == total_offset_8 ? phv_data_228 : _GEN_4787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4789 = 8'he5 == total_offset_8 ? phv_data_229 : _GEN_4788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4790 = 8'he6 == total_offset_8 ? phv_data_230 : _GEN_4789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4791 = 8'he7 == total_offset_8 ? phv_data_231 : _GEN_4790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4792 = 8'he8 == total_offset_8 ? phv_data_232 : _GEN_4791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4793 = 8'he9 == total_offset_8 ? phv_data_233 : _GEN_4792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4794 = 8'hea == total_offset_8 ? phv_data_234 : _GEN_4793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4795 = 8'heb == total_offset_8 ? phv_data_235 : _GEN_4794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4796 = 8'hec == total_offset_8 ? phv_data_236 : _GEN_4795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4797 = 8'hed == total_offset_8 ? phv_data_237 : _GEN_4796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4798 = 8'hee == total_offset_8 ? phv_data_238 : _GEN_4797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4799 = 8'hef == total_offset_8 ? phv_data_239 : _GEN_4798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4800 = 8'hf0 == total_offset_8 ? phv_data_240 : _GEN_4799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4801 = 8'hf1 == total_offset_8 ? phv_data_241 : _GEN_4800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4802 = 8'hf2 == total_offset_8 ? phv_data_242 : _GEN_4801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4803 = 8'hf3 == total_offset_8 ? phv_data_243 : _GEN_4802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4804 = 8'hf4 == total_offset_8 ? phv_data_244 : _GEN_4803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4805 = 8'hf5 == total_offset_8 ? phv_data_245 : _GEN_4804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4806 = 8'hf6 == total_offset_8 ? phv_data_246 : _GEN_4805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4807 = 8'hf7 == total_offset_8 ? phv_data_247 : _GEN_4806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4808 = 8'hf8 == total_offset_8 ? phv_data_248 : _GEN_4807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4809 = 8'hf9 == total_offset_8 ? phv_data_249 : _GEN_4808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4810 = 8'hfa == total_offset_8 ? phv_data_250 : _GEN_4809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4811 = 8'hfb == total_offset_8 ? phv_data_251 : _GEN_4810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4812 = 8'hfc == total_offset_8 ? phv_data_252 : _GEN_4811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4813 = 8'hfd == total_offset_8 ? phv_data_253 : _GEN_4812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4814 = 8'hfe == total_offset_8 ? phv_data_254 : _GEN_4813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4815 = 8'hff == total_offset_8 ? phv_data_255 : _GEN_4814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_11183 = {{1'd0}, total_offset_8}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4816 = 9'h100 == _GEN_11183 ? phv_data_256 : _GEN_4815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4817 = 9'h101 == _GEN_11183 ? phv_data_257 : _GEN_4816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4818 = 9'h102 == _GEN_11183 ? phv_data_258 : _GEN_4817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4819 = 9'h103 == _GEN_11183 ? phv_data_259 : _GEN_4818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4820 = 9'h104 == _GEN_11183 ? phv_data_260 : _GEN_4819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4821 = 9'h105 == _GEN_11183 ? phv_data_261 : _GEN_4820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4822 = 9'h106 == _GEN_11183 ? phv_data_262 : _GEN_4821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4823 = 9'h107 == _GEN_11183 ? phv_data_263 : _GEN_4822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4824 = 9'h108 == _GEN_11183 ? phv_data_264 : _GEN_4823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4825 = 9'h109 == _GEN_11183 ? phv_data_265 : _GEN_4824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4826 = 9'h10a == _GEN_11183 ? phv_data_266 : _GEN_4825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4827 = 9'h10b == _GEN_11183 ? phv_data_267 : _GEN_4826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4828 = 9'h10c == _GEN_11183 ? phv_data_268 : _GEN_4827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4829 = 9'h10d == _GEN_11183 ? phv_data_269 : _GEN_4828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4830 = 9'h10e == _GEN_11183 ? phv_data_270 : _GEN_4829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4831 = 9'h10f == _GEN_11183 ? phv_data_271 : _GEN_4830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4832 = 9'h110 == _GEN_11183 ? phv_data_272 : _GEN_4831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4833 = 9'h111 == _GEN_11183 ? phv_data_273 : _GEN_4832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4834 = 9'h112 == _GEN_11183 ? phv_data_274 : _GEN_4833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4835 = 9'h113 == _GEN_11183 ? phv_data_275 : _GEN_4834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4836 = 9'h114 == _GEN_11183 ? phv_data_276 : _GEN_4835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4837 = 9'h115 == _GEN_11183 ? phv_data_277 : _GEN_4836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4838 = 9'h116 == _GEN_11183 ? phv_data_278 : _GEN_4837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4839 = 9'h117 == _GEN_11183 ? phv_data_279 : _GEN_4838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4840 = 9'h118 == _GEN_11183 ? phv_data_280 : _GEN_4839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4841 = 9'h119 == _GEN_11183 ? phv_data_281 : _GEN_4840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4842 = 9'h11a == _GEN_11183 ? phv_data_282 : _GEN_4841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4843 = 9'h11b == _GEN_11183 ? phv_data_283 : _GEN_4842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4844 = 9'h11c == _GEN_11183 ? phv_data_284 : _GEN_4843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4845 = 9'h11d == _GEN_11183 ? phv_data_285 : _GEN_4844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4846 = 9'h11e == _GEN_11183 ? phv_data_286 : _GEN_4845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4847 = 9'h11f == _GEN_11183 ? phv_data_287 : _GEN_4846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4848 = 9'h120 == _GEN_11183 ? phv_data_288 : _GEN_4847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4849 = 9'h121 == _GEN_11183 ? phv_data_289 : _GEN_4848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4850 = 9'h122 == _GEN_11183 ? phv_data_290 : _GEN_4849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4851 = 9'h123 == _GEN_11183 ? phv_data_291 : _GEN_4850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4852 = 9'h124 == _GEN_11183 ? phv_data_292 : _GEN_4851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4853 = 9'h125 == _GEN_11183 ? phv_data_293 : _GEN_4852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4854 = 9'h126 == _GEN_11183 ? phv_data_294 : _GEN_4853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4855 = 9'h127 == _GEN_11183 ? phv_data_295 : _GEN_4854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4856 = 9'h128 == _GEN_11183 ? phv_data_296 : _GEN_4855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4857 = 9'h129 == _GEN_11183 ? phv_data_297 : _GEN_4856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4858 = 9'h12a == _GEN_11183 ? phv_data_298 : _GEN_4857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4859 = 9'h12b == _GEN_11183 ? phv_data_299 : _GEN_4858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4860 = 9'h12c == _GEN_11183 ? phv_data_300 : _GEN_4859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4861 = 9'h12d == _GEN_11183 ? phv_data_301 : _GEN_4860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4862 = 9'h12e == _GEN_11183 ? phv_data_302 : _GEN_4861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4863 = 9'h12f == _GEN_11183 ? phv_data_303 : _GEN_4862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4864 = 9'h130 == _GEN_11183 ? phv_data_304 : _GEN_4863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4865 = 9'h131 == _GEN_11183 ? phv_data_305 : _GEN_4864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4866 = 9'h132 == _GEN_11183 ? phv_data_306 : _GEN_4865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4867 = 9'h133 == _GEN_11183 ? phv_data_307 : _GEN_4866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4868 = 9'h134 == _GEN_11183 ? phv_data_308 : _GEN_4867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4869 = 9'h135 == _GEN_11183 ? phv_data_309 : _GEN_4868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4870 = 9'h136 == _GEN_11183 ? phv_data_310 : _GEN_4869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4871 = 9'h137 == _GEN_11183 ? phv_data_311 : _GEN_4870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4872 = 9'h138 == _GEN_11183 ? phv_data_312 : _GEN_4871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4873 = 9'h139 == _GEN_11183 ? phv_data_313 : _GEN_4872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4874 = 9'h13a == _GEN_11183 ? phv_data_314 : _GEN_4873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4875 = 9'h13b == _GEN_11183 ? phv_data_315 : _GEN_4874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4876 = 9'h13c == _GEN_11183 ? phv_data_316 : _GEN_4875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4877 = 9'h13d == _GEN_11183 ? phv_data_317 : _GEN_4876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4878 = 9'h13e == _GEN_11183 ? phv_data_318 : _GEN_4877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4879 = 9'h13f == _GEN_11183 ? phv_data_319 : _GEN_4878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4880 = 9'h140 == _GEN_11183 ? phv_data_320 : _GEN_4879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4881 = 9'h141 == _GEN_11183 ? phv_data_321 : _GEN_4880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4882 = 9'h142 == _GEN_11183 ? phv_data_322 : _GEN_4881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4883 = 9'h143 == _GEN_11183 ? phv_data_323 : _GEN_4882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4884 = 9'h144 == _GEN_11183 ? phv_data_324 : _GEN_4883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4885 = 9'h145 == _GEN_11183 ? phv_data_325 : _GEN_4884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4886 = 9'h146 == _GEN_11183 ? phv_data_326 : _GEN_4885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4887 = 9'h147 == _GEN_11183 ? phv_data_327 : _GEN_4886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4888 = 9'h148 == _GEN_11183 ? phv_data_328 : _GEN_4887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4889 = 9'h149 == _GEN_11183 ? phv_data_329 : _GEN_4888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4890 = 9'h14a == _GEN_11183 ? phv_data_330 : _GEN_4889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4891 = 9'h14b == _GEN_11183 ? phv_data_331 : _GEN_4890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4892 = 9'h14c == _GEN_11183 ? phv_data_332 : _GEN_4891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4893 = 9'h14d == _GEN_11183 ? phv_data_333 : _GEN_4892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4894 = 9'h14e == _GEN_11183 ? phv_data_334 : _GEN_4893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4895 = 9'h14f == _GEN_11183 ? phv_data_335 : _GEN_4894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4896 = 9'h150 == _GEN_11183 ? phv_data_336 : _GEN_4895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4897 = 9'h151 == _GEN_11183 ? phv_data_337 : _GEN_4896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4898 = 9'h152 == _GEN_11183 ? phv_data_338 : _GEN_4897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4899 = 9'h153 == _GEN_11183 ? phv_data_339 : _GEN_4898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4900 = 9'h154 == _GEN_11183 ? phv_data_340 : _GEN_4899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4901 = 9'h155 == _GEN_11183 ? phv_data_341 : _GEN_4900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4902 = 9'h156 == _GEN_11183 ? phv_data_342 : _GEN_4901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4903 = 9'h157 == _GEN_11183 ? phv_data_343 : _GEN_4902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4904 = 9'h158 == _GEN_11183 ? phv_data_344 : _GEN_4903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4905 = 9'h159 == _GEN_11183 ? phv_data_345 : _GEN_4904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4906 = 9'h15a == _GEN_11183 ? phv_data_346 : _GEN_4905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4907 = 9'h15b == _GEN_11183 ? phv_data_347 : _GEN_4906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4908 = 9'h15c == _GEN_11183 ? phv_data_348 : _GEN_4907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4909 = 9'h15d == _GEN_11183 ? phv_data_349 : _GEN_4908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4910 = 9'h15e == _GEN_11183 ? phv_data_350 : _GEN_4909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4911 = 9'h15f == _GEN_11183 ? phv_data_351 : _GEN_4910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4912 = 9'h160 == _GEN_11183 ? phv_data_352 : _GEN_4911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4913 = 9'h161 == _GEN_11183 ? phv_data_353 : _GEN_4912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4914 = 9'h162 == _GEN_11183 ? phv_data_354 : _GEN_4913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4915 = 9'h163 == _GEN_11183 ? phv_data_355 : _GEN_4914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4916 = 9'h164 == _GEN_11183 ? phv_data_356 : _GEN_4915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4917 = 9'h165 == _GEN_11183 ? phv_data_357 : _GEN_4916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4918 = 9'h166 == _GEN_11183 ? phv_data_358 : _GEN_4917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4919 = 9'h167 == _GEN_11183 ? phv_data_359 : _GEN_4918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4920 = 9'h168 == _GEN_11183 ? phv_data_360 : _GEN_4919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4921 = 9'h169 == _GEN_11183 ? phv_data_361 : _GEN_4920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4922 = 9'h16a == _GEN_11183 ? phv_data_362 : _GEN_4921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4923 = 9'h16b == _GEN_11183 ? phv_data_363 : _GEN_4922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4924 = 9'h16c == _GEN_11183 ? phv_data_364 : _GEN_4923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4925 = 9'h16d == _GEN_11183 ? phv_data_365 : _GEN_4924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4926 = 9'h16e == _GEN_11183 ? phv_data_366 : _GEN_4925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4927 = 9'h16f == _GEN_11183 ? phv_data_367 : _GEN_4926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4928 = 9'h170 == _GEN_11183 ? phv_data_368 : _GEN_4927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4929 = 9'h171 == _GEN_11183 ? phv_data_369 : _GEN_4928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4930 = 9'h172 == _GEN_11183 ? phv_data_370 : _GEN_4929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4931 = 9'h173 == _GEN_11183 ? phv_data_371 : _GEN_4930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4932 = 9'h174 == _GEN_11183 ? phv_data_372 : _GEN_4931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4933 = 9'h175 == _GEN_11183 ? phv_data_373 : _GEN_4932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4934 = 9'h176 == _GEN_11183 ? phv_data_374 : _GEN_4933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4935 = 9'h177 == _GEN_11183 ? phv_data_375 : _GEN_4934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4936 = 9'h178 == _GEN_11183 ? phv_data_376 : _GEN_4935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4937 = 9'h179 == _GEN_11183 ? phv_data_377 : _GEN_4936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4938 = 9'h17a == _GEN_11183 ? phv_data_378 : _GEN_4937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4939 = 9'h17b == _GEN_11183 ? phv_data_379 : _GEN_4938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4940 = 9'h17c == _GEN_11183 ? phv_data_380 : _GEN_4939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4941 = 9'h17d == _GEN_11183 ? phv_data_381 : _GEN_4940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4942 = 9'h17e == _GEN_11183 ? phv_data_382 : _GEN_4941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4943 = 9'h17f == _GEN_11183 ? phv_data_383 : _GEN_4942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4944 = 9'h180 == _GEN_11183 ? phv_data_384 : _GEN_4943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4945 = 9'h181 == _GEN_11183 ? phv_data_385 : _GEN_4944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4946 = 9'h182 == _GEN_11183 ? phv_data_386 : _GEN_4945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4947 = 9'h183 == _GEN_11183 ? phv_data_387 : _GEN_4946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4948 = 9'h184 == _GEN_11183 ? phv_data_388 : _GEN_4947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4949 = 9'h185 == _GEN_11183 ? phv_data_389 : _GEN_4948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4950 = 9'h186 == _GEN_11183 ? phv_data_390 : _GEN_4949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4951 = 9'h187 == _GEN_11183 ? phv_data_391 : _GEN_4950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4952 = 9'h188 == _GEN_11183 ? phv_data_392 : _GEN_4951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4953 = 9'h189 == _GEN_11183 ? phv_data_393 : _GEN_4952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4954 = 9'h18a == _GEN_11183 ? phv_data_394 : _GEN_4953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4955 = 9'h18b == _GEN_11183 ? phv_data_395 : _GEN_4954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4956 = 9'h18c == _GEN_11183 ? phv_data_396 : _GEN_4955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4957 = 9'h18d == _GEN_11183 ? phv_data_397 : _GEN_4956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4958 = 9'h18e == _GEN_11183 ? phv_data_398 : _GEN_4957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4959 = 9'h18f == _GEN_11183 ? phv_data_399 : _GEN_4958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4960 = 9'h190 == _GEN_11183 ? phv_data_400 : _GEN_4959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4961 = 9'h191 == _GEN_11183 ? phv_data_401 : _GEN_4960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4962 = 9'h192 == _GEN_11183 ? phv_data_402 : _GEN_4961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4963 = 9'h193 == _GEN_11183 ? phv_data_403 : _GEN_4962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4964 = 9'h194 == _GEN_11183 ? phv_data_404 : _GEN_4963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4965 = 9'h195 == _GEN_11183 ? phv_data_405 : _GEN_4964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4966 = 9'h196 == _GEN_11183 ? phv_data_406 : _GEN_4965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4967 = 9'h197 == _GEN_11183 ? phv_data_407 : _GEN_4966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4968 = 9'h198 == _GEN_11183 ? phv_data_408 : _GEN_4967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4969 = 9'h199 == _GEN_11183 ? phv_data_409 : _GEN_4968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4970 = 9'h19a == _GEN_11183 ? phv_data_410 : _GEN_4969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4971 = 9'h19b == _GEN_11183 ? phv_data_411 : _GEN_4970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4972 = 9'h19c == _GEN_11183 ? phv_data_412 : _GEN_4971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4973 = 9'h19d == _GEN_11183 ? phv_data_413 : _GEN_4972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4974 = 9'h19e == _GEN_11183 ? phv_data_414 : _GEN_4973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4975 = 9'h19f == _GEN_11183 ? phv_data_415 : _GEN_4974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4976 = 9'h1a0 == _GEN_11183 ? phv_data_416 : _GEN_4975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4977 = 9'h1a1 == _GEN_11183 ? phv_data_417 : _GEN_4976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4978 = 9'h1a2 == _GEN_11183 ? phv_data_418 : _GEN_4977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4979 = 9'h1a3 == _GEN_11183 ? phv_data_419 : _GEN_4978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4980 = 9'h1a4 == _GEN_11183 ? phv_data_420 : _GEN_4979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4981 = 9'h1a5 == _GEN_11183 ? phv_data_421 : _GEN_4980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4982 = 9'h1a6 == _GEN_11183 ? phv_data_422 : _GEN_4981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4983 = 9'h1a7 == _GEN_11183 ? phv_data_423 : _GEN_4982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4984 = 9'h1a8 == _GEN_11183 ? phv_data_424 : _GEN_4983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4985 = 9'h1a9 == _GEN_11183 ? phv_data_425 : _GEN_4984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4986 = 9'h1aa == _GEN_11183 ? phv_data_426 : _GEN_4985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4987 = 9'h1ab == _GEN_11183 ? phv_data_427 : _GEN_4986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4988 = 9'h1ac == _GEN_11183 ? phv_data_428 : _GEN_4987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4989 = 9'h1ad == _GEN_11183 ? phv_data_429 : _GEN_4988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4990 = 9'h1ae == _GEN_11183 ? phv_data_430 : _GEN_4989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4991 = 9'h1af == _GEN_11183 ? phv_data_431 : _GEN_4990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4992 = 9'h1b0 == _GEN_11183 ? phv_data_432 : _GEN_4991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4993 = 9'h1b1 == _GEN_11183 ? phv_data_433 : _GEN_4992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4994 = 9'h1b2 == _GEN_11183 ? phv_data_434 : _GEN_4993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4995 = 9'h1b3 == _GEN_11183 ? phv_data_435 : _GEN_4994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4996 = 9'h1b4 == _GEN_11183 ? phv_data_436 : _GEN_4995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4997 = 9'h1b5 == _GEN_11183 ? phv_data_437 : _GEN_4996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4998 = 9'h1b6 == _GEN_11183 ? phv_data_438 : _GEN_4997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_4999 = 9'h1b7 == _GEN_11183 ? phv_data_439 : _GEN_4998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5000 = 9'h1b8 == _GEN_11183 ? phv_data_440 : _GEN_4999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5001 = 9'h1b9 == _GEN_11183 ? phv_data_441 : _GEN_5000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5002 = 9'h1ba == _GEN_11183 ? phv_data_442 : _GEN_5001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5003 = 9'h1bb == _GEN_11183 ? phv_data_443 : _GEN_5002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5004 = 9'h1bc == _GEN_11183 ? phv_data_444 : _GEN_5003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5005 = 9'h1bd == _GEN_11183 ? phv_data_445 : _GEN_5004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5006 = 9'h1be == _GEN_11183 ? phv_data_446 : _GEN_5005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5007 = 9'h1bf == _GEN_11183 ? phv_data_447 : _GEN_5006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5008 = 9'h1c0 == _GEN_11183 ? phv_data_448 : _GEN_5007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5009 = 9'h1c1 == _GEN_11183 ? phv_data_449 : _GEN_5008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5010 = 9'h1c2 == _GEN_11183 ? phv_data_450 : _GEN_5009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5011 = 9'h1c3 == _GEN_11183 ? phv_data_451 : _GEN_5010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5012 = 9'h1c4 == _GEN_11183 ? phv_data_452 : _GEN_5011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5013 = 9'h1c5 == _GEN_11183 ? phv_data_453 : _GEN_5012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5014 = 9'h1c6 == _GEN_11183 ? phv_data_454 : _GEN_5013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5015 = 9'h1c7 == _GEN_11183 ? phv_data_455 : _GEN_5014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5016 = 9'h1c8 == _GEN_11183 ? phv_data_456 : _GEN_5015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5017 = 9'h1c9 == _GEN_11183 ? phv_data_457 : _GEN_5016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5018 = 9'h1ca == _GEN_11183 ? phv_data_458 : _GEN_5017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5019 = 9'h1cb == _GEN_11183 ? phv_data_459 : _GEN_5018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5020 = 9'h1cc == _GEN_11183 ? phv_data_460 : _GEN_5019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5021 = 9'h1cd == _GEN_11183 ? phv_data_461 : _GEN_5020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5022 = 9'h1ce == _GEN_11183 ? phv_data_462 : _GEN_5021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5023 = 9'h1cf == _GEN_11183 ? phv_data_463 : _GEN_5022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5024 = 9'h1d0 == _GEN_11183 ? phv_data_464 : _GEN_5023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5025 = 9'h1d1 == _GEN_11183 ? phv_data_465 : _GEN_5024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5026 = 9'h1d2 == _GEN_11183 ? phv_data_466 : _GEN_5025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5027 = 9'h1d3 == _GEN_11183 ? phv_data_467 : _GEN_5026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5028 = 9'h1d4 == _GEN_11183 ? phv_data_468 : _GEN_5027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5029 = 9'h1d5 == _GEN_11183 ? phv_data_469 : _GEN_5028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5030 = 9'h1d6 == _GEN_11183 ? phv_data_470 : _GEN_5029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5031 = 9'h1d7 == _GEN_11183 ? phv_data_471 : _GEN_5030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5032 = 9'h1d8 == _GEN_11183 ? phv_data_472 : _GEN_5031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5033 = 9'h1d9 == _GEN_11183 ? phv_data_473 : _GEN_5032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5034 = 9'h1da == _GEN_11183 ? phv_data_474 : _GEN_5033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5035 = 9'h1db == _GEN_11183 ? phv_data_475 : _GEN_5034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5036 = 9'h1dc == _GEN_11183 ? phv_data_476 : _GEN_5035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5037 = 9'h1dd == _GEN_11183 ? phv_data_477 : _GEN_5036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5038 = 9'h1de == _GEN_11183 ? phv_data_478 : _GEN_5037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5039 = 9'h1df == _GEN_11183 ? phv_data_479 : _GEN_5038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5040 = 9'h1e0 == _GEN_11183 ? phv_data_480 : _GEN_5039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5041 = 9'h1e1 == _GEN_11183 ? phv_data_481 : _GEN_5040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5042 = 9'h1e2 == _GEN_11183 ? phv_data_482 : _GEN_5041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5043 = 9'h1e3 == _GEN_11183 ? phv_data_483 : _GEN_5042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5044 = 9'h1e4 == _GEN_11183 ? phv_data_484 : _GEN_5043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5045 = 9'h1e5 == _GEN_11183 ? phv_data_485 : _GEN_5044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5046 = 9'h1e6 == _GEN_11183 ? phv_data_486 : _GEN_5045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5047 = 9'h1e7 == _GEN_11183 ? phv_data_487 : _GEN_5046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5048 = 9'h1e8 == _GEN_11183 ? phv_data_488 : _GEN_5047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5049 = 9'h1e9 == _GEN_11183 ? phv_data_489 : _GEN_5048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5050 = 9'h1ea == _GEN_11183 ? phv_data_490 : _GEN_5049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5051 = 9'h1eb == _GEN_11183 ? phv_data_491 : _GEN_5050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5052 = 9'h1ec == _GEN_11183 ? phv_data_492 : _GEN_5051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5053 = 9'h1ed == _GEN_11183 ? phv_data_493 : _GEN_5052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5054 = 9'h1ee == _GEN_11183 ? phv_data_494 : _GEN_5053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5055 = 9'h1ef == _GEN_11183 ? phv_data_495 : _GEN_5054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5056 = 9'h1f0 == _GEN_11183 ? phv_data_496 : _GEN_5055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5057 = 9'h1f1 == _GEN_11183 ? phv_data_497 : _GEN_5056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5058 = 9'h1f2 == _GEN_11183 ? phv_data_498 : _GEN_5057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5059 = 9'h1f3 == _GEN_11183 ? phv_data_499 : _GEN_5058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5060 = 9'h1f4 == _GEN_11183 ? phv_data_500 : _GEN_5059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5061 = 9'h1f5 == _GEN_11183 ? phv_data_501 : _GEN_5060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5062 = 9'h1f6 == _GEN_11183 ? phv_data_502 : _GEN_5061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5063 = 9'h1f7 == _GEN_11183 ? phv_data_503 : _GEN_5062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5064 = 9'h1f8 == _GEN_11183 ? phv_data_504 : _GEN_5063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5065 = 9'h1f9 == _GEN_11183 ? phv_data_505 : _GEN_5064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5066 = 9'h1fa == _GEN_11183 ? phv_data_506 : _GEN_5065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5067 = 9'h1fb == _GEN_11183 ? phv_data_507 : _GEN_5066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5068 = 9'h1fc == _GEN_11183 ? phv_data_508 : _GEN_5067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5069 = 9'h1fd == _GEN_11183 ? phv_data_509 : _GEN_5068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5070 = 9'h1fe == _GEN_11183 ? phv_data_510 : _GEN_5069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_3 = 9'h1ff == _GEN_11183 ? phv_data_511 : _GEN_5070; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_17 = ending_2 == 2'h0; // @[executor.scala 199:88]
  wire  mask_2_3 = 2'h0 >= offset_2[1:0] & (2'h0 < ending_2 | ending_2 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_9 = {total_offset_hi_2,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_5073 = 8'h1 == total_offset_9 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5074 = 8'h2 == total_offset_9 ? phv_data_2 : _GEN_5073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5075 = 8'h3 == total_offset_9 ? phv_data_3 : _GEN_5074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5076 = 8'h4 == total_offset_9 ? phv_data_4 : _GEN_5075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5077 = 8'h5 == total_offset_9 ? phv_data_5 : _GEN_5076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5078 = 8'h6 == total_offset_9 ? phv_data_6 : _GEN_5077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5079 = 8'h7 == total_offset_9 ? phv_data_7 : _GEN_5078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5080 = 8'h8 == total_offset_9 ? phv_data_8 : _GEN_5079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5081 = 8'h9 == total_offset_9 ? phv_data_9 : _GEN_5080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5082 = 8'ha == total_offset_9 ? phv_data_10 : _GEN_5081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5083 = 8'hb == total_offset_9 ? phv_data_11 : _GEN_5082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5084 = 8'hc == total_offset_9 ? phv_data_12 : _GEN_5083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5085 = 8'hd == total_offset_9 ? phv_data_13 : _GEN_5084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5086 = 8'he == total_offset_9 ? phv_data_14 : _GEN_5085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5087 = 8'hf == total_offset_9 ? phv_data_15 : _GEN_5086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5088 = 8'h10 == total_offset_9 ? phv_data_16 : _GEN_5087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5089 = 8'h11 == total_offset_9 ? phv_data_17 : _GEN_5088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5090 = 8'h12 == total_offset_9 ? phv_data_18 : _GEN_5089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5091 = 8'h13 == total_offset_9 ? phv_data_19 : _GEN_5090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5092 = 8'h14 == total_offset_9 ? phv_data_20 : _GEN_5091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5093 = 8'h15 == total_offset_9 ? phv_data_21 : _GEN_5092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5094 = 8'h16 == total_offset_9 ? phv_data_22 : _GEN_5093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5095 = 8'h17 == total_offset_9 ? phv_data_23 : _GEN_5094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5096 = 8'h18 == total_offset_9 ? phv_data_24 : _GEN_5095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5097 = 8'h19 == total_offset_9 ? phv_data_25 : _GEN_5096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5098 = 8'h1a == total_offset_9 ? phv_data_26 : _GEN_5097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5099 = 8'h1b == total_offset_9 ? phv_data_27 : _GEN_5098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5100 = 8'h1c == total_offset_9 ? phv_data_28 : _GEN_5099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5101 = 8'h1d == total_offset_9 ? phv_data_29 : _GEN_5100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5102 = 8'h1e == total_offset_9 ? phv_data_30 : _GEN_5101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5103 = 8'h1f == total_offset_9 ? phv_data_31 : _GEN_5102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5104 = 8'h20 == total_offset_9 ? phv_data_32 : _GEN_5103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5105 = 8'h21 == total_offset_9 ? phv_data_33 : _GEN_5104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5106 = 8'h22 == total_offset_9 ? phv_data_34 : _GEN_5105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5107 = 8'h23 == total_offset_9 ? phv_data_35 : _GEN_5106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5108 = 8'h24 == total_offset_9 ? phv_data_36 : _GEN_5107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5109 = 8'h25 == total_offset_9 ? phv_data_37 : _GEN_5108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5110 = 8'h26 == total_offset_9 ? phv_data_38 : _GEN_5109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5111 = 8'h27 == total_offset_9 ? phv_data_39 : _GEN_5110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5112 = 8'h28 == total_offset_9 ? phv_data_40 : _GEN_5111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5113 = 8'h29 == total_offset_9 ? phv_data_41 : _GEN_5112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5114 = 8'h2a == total_offset_9 ? phv_data_42 : _GEN_5113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5115 = 8'h2b == total_offset_9 ? phv_data_43 : _GEN_5114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5116 = 8'h2c == total_offset_9 ? phv_data_44 : _GEN_5115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5117 = 8'h2d == total_offset_9 ? phv_data_45 : _GEN_5116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5118 = 8'h2e == total_offset_9 ? phv_data_46 : _GEN_5117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5119 = 8'h2f == total_offset_9 ? phv_data_47 : _GEN_5118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5120 = 8'h30 == total_offset_9 ? phv_data_48 : _GEN_5119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5121 = 8'h31 == total_offset_9 ? phv_data_49 : _GEN_5120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5122 = 8'h32 == total_offset_9 ? phv_data_50 : _GEN_5121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5123 = 8'h33 == total_offset_9 ? phv_data_51 : _GEN_5122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5124 = 8'h34 == total_offset_9 ? phv_data_52 : _GEN_5123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5125 = 8'h35 == total_offset_9 ? phv_data_53 : _GEN_5124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5126 = 8'h36 == total_offset_9 ? phv_data_54 : _GEN_5125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5127 = 8'h37 == total_offset_9 ? phv_data_55 : _GEN_5126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5128 = 8'h38 == total_offset_9 ? phv_data_56 : _GEN_5127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5129 = 8'h39 == total_offset_9 ? phv_data_57 : _GEN_5128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5130 = 8'h3a == total_offset_9 ? phv_data_58 : _GEN_5129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5131 = 8'h3b == total_offset_9 ? phv_data_59 : _GEN_5130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5132 = 8'h3c == total_offset_9 ? phv_data_60 : _GEN_5131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5133 = 8'h3d == total_offset_9 ? phv_data_61 : _GEN_5132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5134 = 8'h3e == total_offset_9 ? phv_data_62 : _GEN_5133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5135 = 8'h3f == total_offset_9 ? phv_data_63 : _GEN_5134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5136 = 8'h40 == total_offset_9 ? phv_data_64 : _GEN_5135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5137 = 8'h41 == total_offset_9 ? phv_data_65 : _GEN_5136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5138 = 8'h42 == total_offset_9 ? phv_data_66 : _GEN_5137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5139 = 8'h43 == total_offset_9 ? phv_data_67 : _GEN_5138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5140 = 8'h44 == total_offset_9 ? phv_data_68 : _GEN_5139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5141 = 8'h45 == total_offset_9 ? phv_data_69 : _GEN_5140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5142 = 8'h46 == total_offset_9 ? phv_data_70 : _GEN_5141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5143 = 8'h47 == total_offset_9 ? phv_data_71 : _GEN_5142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5144 = 8'h48 == total_offset_9 ? phv_data_72 : _GEN_5143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5145 = 8'h49 == total_offset_9 ? phv_data_73 : _GEN_5144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5146 = 8'h4a == total_offset_9 ? phv_data_74 : _GEN_5145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5147 = 8'h4b == total_offset_9 ? phv_data_75 : _GEN_5146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5148 = 8'h4c == total_offset_9 ? phv_data_76 : _GEN_5147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5149 = 8'h4d == total_offset_9 ? phv_data_77 : _GEN_5148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5150 = 8'h4e == total_offset_9 ? phv_data_78 : _GEN_5149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5151 = 8'h4f == total_offset_9 ? phv_data_79 : _GEN_5150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5152 = 8'h50 == total_offset_9 ? phv_data_80 : _GEN_5151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5153 = 8'h51 == total_offset_9 ? phv_data_81 : _GEN_5152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5154 = 8'h52 == total_offset_9 ? phv_data_82 : _GEN_5153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5155 = 8'h53 == total_offset_9 ? phv_data_83 : _GEN_5154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5156 = 8'h54 == total_offset_9 ? phv_data_84 : _GEN_5155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5157 = 8'h55 == total_offset_9 ? phv_data_85 : _GEN_5156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5158 = 8'h56 == total_offset_9 ? phv_data_86 : _GEN_5157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5159 = 8'h57 == total_offset_9 ? phv_data_87 : _GEN_5158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5160 = 8'h58 == total_offset_9 ? phv_data_88 : _GEN_5159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5161 = 8'h59 == total_offset_9 ? phv_data_89 : _GEN_5160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5162 = 8'h5a == total_offset_9 ? phv_data_90 : _GEN_5161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5163 = 8'h5b == total_offset_9 ? phv_data_91 : _GEN_5162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5164 = 8'h5c == total_offset_9 ? phv_data_92 : _GEN_5163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5165 = 8'h5d == total_offset_9 ? phv_data_93 : _GEN_5164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5166 = 8'h5e == total_offset_9 ? phv_data_94 : _GEN_5165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5167 = 8'h5f == total_offset_9 ? phv_data_95 : _GEN_5166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5168 = 8'h60 == total_offset_9 ? phv_data_96 : _GEN_5167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5169 = 8'h61 == total_offset_9 ? phv_data_97 : _GEN_5168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5170 = 8'h62 == total_offset_9 ? phv_data_98 : _GEN_5169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5171 = 8'h63 == total_offset_9 ? phv_data_99 : _GEN_5170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5172 = 8'h64 == total_offset_9 ? phv_data_100 : _GEN_5171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5173 = 8'h65 == total_offset_9 ? phv_data_101 : _GEN_5172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5174 = 8'h66 == total_offset_9 ? phv_data_102 : _GEN_5173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5175 = 8'h67 == total_offset_9 ? phv_data_103 : _GEN_5174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5176 = 8'h68 == total_offset_9 ? phv_data_104 : _GEN_5175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5177 = 8'h69 == total_offset_9 ? phv_data_105 : _GEN_5176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5178 = 8'h6a == total_offset_9 ? phv_data_106 : _GEN_5177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5179 = 8'h6b == total_offset_9 ? phv_data_107 : _GEN_5178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5180 = 8'h6c == total_offset_9 ? phv_data_108 : _GEN_5179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5181 = 8'h6d == total_offset_9 ? phv_data_109 : _GEN_5180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5182 = 8'h6e == total_offset_9 ? phv_data_110 : _GEN_5181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5183 = 8'h6f == total_offset_9 ? phv_data_111 : _GEN_5182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5184 = 8'h70 == total_offset_9 ? phv_data_112 : _GEN_5183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5185 = 8'h71 == total_offset_9 ? phv_data_113 : _GEN_5184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5186 = 8'h72 == total_offset_9 ? phv_data_114 : _GEN_5185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5187 = 8'h73 == total_offset_9 ? phv_data_115 : _GEN_5186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5188 = 8'h74 == total_offset_9 ? phv_data_116 : _GEN_5187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5189 = 8'h75 == total_offset_9 ? phv_data_117 : _GEN_5188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5190 = 8'h76 == total_offset_9 ? phv_data_118 : _GEN_5189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5191 = 8'h77 == total_offset_9 ? phv_data_119 : _GEN_5190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5192 = 8'h78 == total_offset_9 ? phv_data_120 : _GEN_5191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5193 = 8'h79 == total_offset_9 ? phv_data_121 : _GEN_5192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5194 = 8'h7a == total_offset_9 ? phv_data_122 : _GEN_5193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5195 = 8'h7b == total_offset_9 ? phv_data_123 : _GEN_5194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5196 = 8'h7c == total_offset_9 ? phv_data_124 : _GEN_5195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5197 = 8'h7d == total_offset_9 ? phv_data_125 : _GEN_5196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5198 = 8'h7e == total_offset_9 ? phv_data_126 : _GEN_5197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5199 = 8'h7f == total_offset_9 ? phv_data_127 : _GEN_5198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5200 = 8'h80 == total_offset_9 ? phv_data_128 : _GEN_5199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5201 = 8'h81 == total_offset_9 ? phv_data_129 : _GEN_5200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5202 = 8'h82 == total_offset_9 ? phv_data_130 : _GEN_5201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5203 = 8'h83 == total_offset_9 ? phv_data_131 : _GEN_5202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5204 = 8'h84 == total_offset_9 ? phv_data_132 : _GEN_5203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5205 = 8'h85 == total_offset_9 ? phv_data_133 : _GEN_5204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5206 = 8'h86 == total_offset_9 ? phv_data_134 : _GEN_5205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5207 = 8'h87 == total_offset_9 ? phv_data_135 : _GEN_5206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5208 = 8'h88 == total_offset_9 ? phv_data_136 : _GEN_5207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5209 = 8'h89 == total_offset_9 ? phv_data_137 : _GEN_5208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5210 = 8'h8a == total_offset_9 ? phv_data_138 : _GEN_5209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5211 = 8'h8b == total_offset_9 ? phv_data_139 : _GEN_5210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5212 = 8'h8c == total_offset_9 ? phv_data_140 : _GEN_5211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5213 = 8'h8d == total_offset_9 ? phv_data_141 : _GEN_5212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5214 = 8'h8e == total_offset_9 ? phv_data_142 : _GEN_5213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5215 = 8'h8f == total_offset_9 ? phv_data_143 : _GEN_5214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5216 = 8'h90 == total_offset_9 ? phv_data_144 : _GEN_5215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5217 = 8'h91 == total_offset_9 ? phv_data_145 : _GEN_5216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5218 = 8'h92 == total_offset_9 ? phv_data_146 : _GEN_5217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5219 = 8'h93 == total_offset_9 ? phv_data_147 : _GEN_5218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5220 = 8'h94 == total_offset_9 ? phv_data_148 : _GEN_5219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5221 = 8'h95 == total_offset_9 ? phv_data_149 : _GEN_5220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5222 = 8'h96 == total_offset_9 ? phv_data_150 : _GEN_5221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5223 = 8'h97 == total_offset_9 ? phv_data_151 : _GEN_5222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5224 = 8'h98 == total_offset_9 ? phv_data_152 : _GEN_5223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5225 = 8'h99 == total_offset_9 ? phv_data_153 : _GEN_5224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5226 = 8'h9a == total_offset_9 ? phv_data_154 : _GEN_5225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5227 = 8'h9b == total_offset_9 ? phv_data_155 : _GEN_5226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5228 = 8'h9c == total_offset_9 ? phv_data_156 : _GEN_5227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5229 = 8'h9d == total_offset_9 ? phv_data_157 : _GEN_5228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5230 = 8'h9e == total_offset_9 ? phv_data_158 : _GEN_5229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5231 = 8'h9f == total_offset_9 ? phv_data_159 : _GEN_5230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5232 = 8'ha0 == total_offset_9 ? phv_data_160 : _GEN_5231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5233 = 8'ha1 == total_offset_9 ? phv_data_161 : _GEN_5232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5234 = 8'ha2 == total_offset_9 ? phv_data_162 : _GEN_5233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5235 = 8'ha3 == total_offset_9 ? phv_data_163 : _GEN_5234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5236 = 8'ha4 == total_offset_9 ? phv_data_164 : _GEN_5235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5237 = 8'ha5 == total_offset_9 ? phv_data_165 : _GEN_5236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5238 = 8'ha6 == total_offset_9 ? phv_data_166 : _GEN_5237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5239 = 8'ha7 == total_offset_9 ? phv_data_167 : _GEN_5238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5240 = 8'ha8 == total_offset_9 ? phv_data_168 : _GEN_5239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5241 = 8'ha9 == total_offset_9 ? phv_data_169 : _GEN_5240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5242 = 8'haa == total_offset_9 ? phv_data_170 : _GEN_5241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5243 = 8'hab == total_offset_9 ? phv_data_171 : _GEN_5242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5244 = 8'hac == total_offset_9 ? phv_data_172 : _GEN_5243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5245 = 8'had == total_offset_9 ? phv_data_173 : _GEN_5244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5246 = 8'hae == total_offset_9 ? phv_data_174 : _GEN_5245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5247 = 8'haf == total_offset_9 ? phv_data_175 : _GEN_5246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5248 = 8'hb0 == total_offset_9 ? phv_data_176 : _GEN_5247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5249 = 8'hb1 == total_offset_9 ? phv_data_177 : _GEN_5248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5250 = 8'hb2 == total_offset_9 ? phv_data_178 : _GEN_5249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5251 = 8'hb3 == total_offset_9 ? phv_data_179 : _GEN_5250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5252 = 8'hb4 == total_offset_9 ? phv_data_180 : _GEN_5251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5253 = 8'hb5 == total_offset_9 ? phv_data_181 : _GEN_5252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5254 = 8'hb6 == total_offset_9 ? phv_data_182 : _GEN_5253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5255 = 8'hb7 == total_offset_9 ? phv_data_183 : _GEN_5254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5256 = 8'hb8 == total_offset_9 ? phv_data_184 : _GEN_5255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5257 = 8'hb9 == total_offset_9 ? phv_data_185 : _GEN_5256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5258 = 8'hba == total_offset_9 ? phv_data_186 : _GEN_5257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5259 = 8'hbb == total_offset_9 ? phv_data_187 : _GEN_5258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5260 = 8'hbc == total_offset_9 ? phv_data_188 : _GEN_5259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5261 = 8'hbd == total_offset_9 ? phv_data_189 : _GEN_5260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5262 = 8'hbe == total_offset_9 ? phv_data_190 : _GEN_5261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5263 = 8'hbf == total_offset_9 ? phv_data_191 : _GEN_5262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5264 = 8'hc0 == total_offset_9 ? phv_data_192 : _GEN_5263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5265 = 8'hc1 == total_offset_9 ? phv_data_193 : _GEN_5264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5266 = 8'hc2 == total_offset_9 ? phv_data_194 : _GEN_5265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5267 = 8'hc3 == total_offset_9 ? phv_data_195 : _GEN_5266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5268 = 8'hc4 == total_offset_9 ? phv_data_196 : _GEN_5267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5269 = 8'hc5 == total_offset_9 ? phv_data_197 : _GEN_5268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5270 = 8'hc6 == total_offset_9 ? phv_data_198 : _GEN_5269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5271 = 8'hc7 == total_offset_9 ? phv_data_199 : _GEN_5270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5272 = 8'hc8 == total_offset_9 ? phv_data_200 : _GEN_5271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5273 = 8'hc9 == total_offset_9 ? phv_data_201 : _GEN_5272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5274 = 8'hca == total_offset_9 ? phv_data_202 : _GEN_5273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5275 = 8'hcb == total_offset_9 ? phv_data_203 : _GEN_5274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5276 = 8'hcc == total_offset_9 ? phv_data_204 : _GEN_5275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5277 = 8'hcd == total_offset_9 ? phv_data_205 : _GEN_5276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5278 = 8'hce == total_offset_9 ? phv_data_206 : _GEN_5277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5279 = 8'hcf == total_offset_9 ? phv_data_207 : _GEN_5278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5280 = 8'hd0 == total_offset_9 ? phv_data_208 : _GEN_5279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5281 = 8'hd1 == total_offset_9 ? phv_data_209 : _GEN_5280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5282 = 8'hd2 == total_offset_9 ? phv_data_210 : _GEN_5281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5283 = 8'hd3 == total_offset_9 ? phv_data_211 : _GEN_5282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5284 = 8'hd4 == total_offset_9 ? phv_data_212 : _GEN_5283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5285 = 8'hd5 == total_offset_9 ? phv_data_213 : _GEN_5284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5286 = 8'hd6 == total_offset_9 ? phv_data_214 : _GEN_5285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5287 = 8'hd7 == total_offset_9 ? phv_data_215 : _GEN_5286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5288 = 8'hd8 == total_offset_9 ? phv_data_216 : _GEN_5287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5289 = 8'hd9 == total_offset_9 ? phv_data_217 : _GEN_5288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5290 = 8'hda == total_offset_9 ? phv_data_218 : _GEN_5289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5291 = 8'hdb == total_offset_9 ? phv_data_219 : _GEN_5290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5292 = 8'hdc == total_offset_9 ? phv_data_220 : _GEN_5291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5293 = 8'hdd == total_offset_9 ? phv_data_221 : _GEN_5292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5294 = 8'hde == total_offset_9 ? phv_data_222 : _GEN_5293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5295 = 8'hdf == total_offset_9 ? phv_data_223 : _GEN_5294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5296 = 8'he0 == total_offset_9 ? phv_data_224 : _GEN_5295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5297 = 8'he1 == total_offset_9 ? phv_data_225 : _GEN_5296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5298 = 8'he2 == total_offset_9 ? phv_data_226 : _GEN_5297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5299 = 8'he3 == total_offset_9 ? phv_data_227 : _GEN_5298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5300 = 8'he4 == total_offset_9 ? phv_data_228 : _GEN_5299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5301 = 8'he5 == total_offset_9 ? phv_data_229 : _GEN_5300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5302 = 8'he6 == total_offset_9 ? phv_data_230 : _GEN_5301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5303 = 8'he7 == total_offset_9 ? phv_data_231 : _GEN_5302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5304 = 8'he8 == total_offset_9 ? phv_data_232 : _GEN_5303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5305 = 8'he9 == total_offset_9 ? phv_data_233 : _GEN_5304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5306 = 8'hea == total_offset_9 ? phv_data_234 : _GEN_5305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5307 = 8'heb == total_offset_9 ? phv_data_235 : _GEN_5306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5308 = 8'hec == total_offset_9 ? phv_data_236 : _GEN_5307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5309 = 8'hed == total_offset_9 ? phv_data_237 : _GEN_5308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5310 = 8'hee == total_offset_9 ? phv_data_238 : _GEN_5309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5311 = 8'hef == total_offset_9 ? phv_data_239 : _GEN_5310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5312 = 8'hf0 == total_offset_9 ? phv_data_240 : _GEN_5311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5313 = 8'hf1 == total_offset_9 ? phv_data_241 : _GEN_5312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5314 = 8'hf2 == total_offset_9 ? phv_data_242 : _GEN_5313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5315 = 8'hf3 == total_offset_9 ? phv_data_243 : _GEN_5314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5316 = 8'hf4 == total_offset_9 ? phv_data_244 : _GEN_5315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5317 = 8'hf5 == total_offset_9 ? phv_data_245 : _GEN_5316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5318 = 8'hf6 == total_offset_9 ? phv_data_246 : _GEN_5317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5319 = 8'hf7 == total_offset_9 ? phv_data_247 : _GEN_5318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5320 = 8'hf8 == total_offset_9 ? phv_data_248 : _GEN_5319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5321 = 8'hf9 == total_offset_9 ? phv_data_249 : _GEN_5320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5322 = 8'hfa == total_offset_9 ? phv_data_250 : _GEN_5321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5323 = 8'hfb == total_offset_9 ? phv_data_251 : _GEN_5322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5324 = 8'hfc == total_offset_9 ? phv_data_252 : _GEN_5323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5325 = 8'hfd == total_offset_9 ? phv_data_253 : _GEN_5324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5326 = 8'hfe == total_offset_9 ? phv_data_254 : _GEN_5325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5327 = 8'hff == total_offset_9 ? phv_data_255 : _GEN_5326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_11439 = {{1'd0}, total_offset_9}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5328 = 9'h100 == _GEN_11439 ? phv_data_256 : _GEN_5327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5329 = 9'h101 == _GEN_11439 ? phv_data_257 : _GEN_5328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5330 = 9'h102 == _GEN_11439 ? phv_data_258 : _GEN_5329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5331 = 9'h103 == _GEN_11439 ? phv_data_259 : _GEN_5330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5332 = 9'h104 == _GEN_11439 ? phv_data_260 : _GEN_5331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5333 = 9'h105 == _GEN_11439 ? phv_data_261 : _GEN_5332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5334 = 9'h106 == _GEN_11439 ? phv_data_262 : _GEN_5333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5335 = 9'h107 == _GEN_11439 ? phv_data_263 : _GEN_5334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5336 = 9'h108 == _GEN_11439 ? phv_data_264 : _GEN_5335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5337 = 9'h109 == _GEN_11439 ? phv_data_265 : _GEN_5336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5338 = 9'h10a == _GEN_11439 ? phv_data_266 : _GEN_5337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5339 = 9'h10b == _GEN_11439 ? phv_data_267 : _GEN_5338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5340 = 9'h10c == _GEN_11439 ? phv_data_268 : _GEN_5339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5341 = 9'h10d == _GEN_11439 ? phv_data_269 : _GEN_5340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5342 = 9'h10e == _GEN_11439 ? phv_data_270 : _GEN_5341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5343 = 9'h10f == _GEN_11439 ? phv_data_271 : _GEN_5342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5344 = 9'h110 == _GEN_11439 ? phv_data_272 : _GEN_5343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5345 = 9'h111 == _GEN_11439 ? phv_data_273 : _GEN_5344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5346 = 9'h112 == _GEN_11439 ? phv_data_274 : _GEN_5345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5347 = 9'h113 == _GEN_11439 ? phv_data_275 : _GEN_5346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5348 = 9'h114 == _GEN_11439 ? phv_data_276 : _GEN_5347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5349 = 9'h115 == _GEN_11439 ? phv_data_277 : _GEN_5348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5350 = 9'h116 == _GEN_11439 ? phv_data_278 : _GEN_5349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5351 = 9'h117 == _GEN_11439 ? phv_data_279 : _GEN_5350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5352 = 9'h118 == _GEN_11439 ? phv_data_280 : _GEN_5351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5353 = 9'h119 == _GEN_11439 ? phv_data_281 : _GEN_5352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5354 = 9'h11a == _GEN_11439 ? phv_data_282 : _GEN_5353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5355 = 9'h11b == _GEN_11439 ? phv_data_283 : _GEN_5354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5356 = 9'h11c == _GEN_11439 ? phv_data_284 : _GEN_5355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5357 = 9'h11d == _GEN_11439 ? phv_data_285 : _GEN_5356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5358 = 9'h11e == _GEN_11439 ? phv_data_286 : _GEN_5357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5359 = 9'h11f == _GEN_11439 ? phv_data_287 : _GEN_5358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5360 = 9'h120 == _GEN_11439 ? phv_data_288 : _GEN_5359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5361 = 9'h121 == _GEN_11439 ? phv_data_289 : _GEN_5360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5362 = 9'h122 == _GEN_11439 ? phv_data_290 : _GEN_5361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5363 = 9'h123 == _GEN_11439 ? phv_data_291 : _GEN_5362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5364 = 9'h124 == _GEN_11439 ? phv_data_292 : _GEN_5363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5365 = 9'h125 == _GEN_11439 ? phv_data_293 : _GEN_5364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5366 = 9'h126 == _GEN_11439 ? phv_data_294 : _GEN_5365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5367 = 9'h127 == _GEN_11439 ? phv_data_295 : _GEN_5366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5368 = 9'h128 == _GEN_11439 ? phv_data_296 : _GEN_5367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5369 = 9'h129 == _GEN_11439 ? phv_data_297 : _GEN_5368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5370 = 9'h12a == _GEN_11439 ? phv_data_298 : _GEN_5369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5371 = 9'h12b == _GEN_11439 ? phv_data_299 : _GEN_5370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5372 = 9'h12c == _GEN_11439 ? phv_data_300 : _GEN_5371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5373 = 9'h12d == _GEN_11439 ? phv_data_301 : _GEN_5372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5374 = 9'h12e == _GEN_11439 ? phv_data_302 : _GEN_5373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5375 = 9'h12f == _GEN_11439 ? phv_data_303 : _GEN_5374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5376 = 9'h130 == _GEN_11439 ? phv_data_304 : _GEN_5375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5377 = 9'h131 == _GEN_11439 ? phv_data_305 : _GEN_5376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5378 = 9'h132 == _GEN_11439 ? phv_data_306 : _GEN_5377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5379 = 9'h133 == _GEN_11439 ? phv_data_307 : _GEN_5378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5380 = 9'h134 == _GEN_11439 ? phv_data_308 : _GEN_5379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5381 = 9'h135 == _GEN_11439 ? phv_data_309 : _GEN_5380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5382 = 9'h136 == _GEN_11439 ? phv_data_310 : _GEN_5381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5383 = 9'h137 == _GEN_11439 ? phv_data_311 : _GEN_5382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5384 = 9'h138 == _GEN_11439 ? phv_data_312 : _GEN_5383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5385 = 9'h139 == _GEN_11439 ? phv_data_313 : _GEN_5384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5386 = 9'h13a == _GEN_11439 ? phv_data_314 : _GEN_5385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5387 = 9'h13b == _GEN_11439 ? phv_data_315 : _GEN_5386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5388 = 9'h13c == _GEN_11439 ? phv_data_316 : _GEN_5387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5389 = 9'h13d == _GEN_11439 ? phv_data_317 : _GEN_5388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5390 = 9'h13e == _GEN_11439 ? phv_data_318 : _GEN_5389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5391 = 9'h13f == _GEN_11439 ? phv_data_319 : _GEN_5390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5392 = 9'h140 == _GEN_11439 ? phv_data_320 : _GEN_5391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5393 = 9'h141 == _GEN_11439 ? phv_data_321 : _GEN_5392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5394 = 9'h142 == _GEN_11439 ? phv_data_322 : _GEN_5393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5395 = 9'h143 == _GEN_11439 ? phv_data_323 : _GEN_5394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5396 = 9'h144 == _GEN_11439 ? phv_data_324 : _GEN_5395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5397 = 9'h145 == _GEN_11439 ? phv_data_325 : _GEN_5396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5398 = 9'h146 == _GEN_11439 ? phv_data_326 : _GEN_5397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5399 = 9'h147 == _GEN_11439 ? phv_data_327 : _GEN_5398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5400 = 9'h148 == _GEN_11439 ? phv_data_328 : _GEN_5399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5401 = 9'h149 == _GEN_11439 ? phv_data_329 : _GEN_5400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5402 = 9'h14a == _GEN_11439 ? phv_data_330 : _GEN_5401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5403 = 9'h14b == _GEN_11439 ? phv_data_331 : _GEN_5402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5404 = 9'h14c == _GEN_11439 ? phv_data_332 : _GEN_5403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5405 = 9'h14d == _GEN_11439 ? phv_data_333 : _GEN_5404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5406 = 9'h14e == _GEN_11439 ? phv_data_334 : _GEN_5405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5407 = 9'h14f == _GEN_11439 ? phv_data_335 : _GEN_5406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5408 = 9'h150 == _GEN_11439 ? phv_data_336 : _GEN_5407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5409 = 9'h151 == _GEN_11439 ? phv_data_337 : _GEN_5408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5410 = 9'h152 == _GEN_11439 ? phv_data_338 : _GEN_5409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5411 = 9'h153 == _GEN_11439 ? phv_data_339 : _GEN_5410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5412 = 9'h154 == _GEN_11439 ? phv_data_340 : _GEN_5411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5413 = 9'h155 == _GEN_11439 ? phv_data_341 : _GEN_5412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5414 = 9'h156 == _GEN_11439 ? phv_data_342 : _GEN_5413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5415 = 9'h157 == _GEN_11439 ? phv_data_343 : _GEN_5414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5416 = 9'h158 == _GEN_11439 ? phv_data_344 : _GEN_5415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5417 = 9'h159 == _GEN_11439 ? phv_data_345 : _GEN_5416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5418 = 9'h15a == _GEN_11439 ? phv_data_346 : _GEN_5417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5419 = 9'h15b == _GEN_11439 ? phv_data_347 : _GEN_5418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5420 = 9'h15c == _GEN_11439 ? phv_data_348 : _GEN_5419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5421 = 9'h15d == _GEN_11439 ? phv_data_349 : _GEN_5420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5422 = 9'h15e == _GEN_11439 ? phv_data_350 : _GEN_5421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5423 = 9'h15f == _GEN_11439 ? phv_data_351 : _GEN_5422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5424 = 9'h160 == _GEN_11439 ? phv_data_352 : _GEN_5423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5425 = 9'h161 == _GEN_11439 ? phv_data_353 : _GEN_5424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5426 = 9'h162 == _GEN_11439 ? phv_data_354 : _GEN_5425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5427 = 9'h163 == _GEN_11439 ? phv_data_355 : _GEN_5426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5428 = 9'h164 == _GEN_11439 ? phv_data_356 : _GEN_5427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5429 = 9'h165 == _GEN_11439 ? phv_data_357 : _GEN_5428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5430 = 9'h166 == _GEN_11439 ? phv_data_358 : _GEN_5429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5431 = 9'h167 == _GEN_11439 ? phv_data_359 : _GEN_5430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5432 = 9'h168 == _GEN_11439 ? phv_data_360 : _GEN_5431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5433 = 9'h169 == _GEN_11439 ? phv_data_361 : _GEN_5432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5434 = 9'h16a == _GEN_11439 ? phv_data_362 : _GEN_5433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5435 = 9'h16b == _GEN_11439 ? phv_data_363 : _GEN_5434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5436 = 9'h16c == _GEN_11439 ? phv_data_364 : _GEN_5435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5437 = 9'h16d == _GEN_11439 ? phv_data_365 : _GEN_5436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5438 = 9'h16e == _GEN_11439 ? phv_data_366 : _GEN_5437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5439 = 9'h16f == _GEN_11439 ? phv_data_367 : _GEN_5438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5440 = 9'h170 == _GEN_11439 ? phv_data_368 : _GEN_5439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5441 = 9'h171 == _GEN_11439 ? phv_data_369 : _GEN_5440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5442 = 9'h172 == _GEN_11439 ? phv_data_370 : _GEN_5441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5443 = 9'h173 == _GEN_11439 ? phv_data_371 : _GEN_5442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5444 = 9'h174 == _GEN_11439 ? phv_data_372 : _GEN_5443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5445 = 9'h175 == _GEN_11439 ? phv_data_373 : _GEN_5444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5446 = 9'h176 == _GEN_11439 ? phv_data_374 : _GEN_5445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5447 = 9'h177 == _GEN_11439 ? phv_data_375 : _GEN_5446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5448 = 9'h178 == _GEN_11439 ? phv_data_376 : _GEN_5447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5449 = 9'h179 == _GEN_11439 ? phv_data_377 : _GEN_5448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5450 = 9'h17a == _GEN_11439 ? phv_data_378 : _GEN_5449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5451 = 9'h17b == _GEN_11439 ? phv_data_379 : _GEN_5450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5452 = 9'h17c == _GEN_11439 ? phv_data_380 : _GEN_5451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5453 = 9'h17d == _GEN_11439 ? phv_data_381 : _GEN_5452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5454 = 9'h17e == _GEN_11439 ? phv_data_382 : _GEN_5453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5455 = 9'h17f == _GEN_11439 ? phv_data_383 : _GEN_5454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5456 = 9'h180 == _GEN_11439 ? phv_data_384 : _GEN_5455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5457 = 9'h181 == _GEN_11439 ? phv_data_385 : _GEN_5456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5458 = 9'h182 == _GEN_11439 ? phv_data_386 : _GEN_5457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5459 = 9'h183 == _GEN_11439 ? phv_data_387 : _GEN_5458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5460 = 9'h184 == _GEN_11439 ? phv_data_388 : _GEN_5459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5461 = 9'h185 == _GEN_11439 ? phv_data_389 : _GEN_5460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5462 = 9'h186 == _GEN_11439 ? phv_data_390 : _GEN_5461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5463 = 9'h187 == _GEN_11439 ? phv_data_391 : _GEN_5462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5464 = 9'h188 == _GEN_11439 ? phv_data_392 : _GEN_5463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5465 = 9'h189 == _GEN_11439 ? phv_data_393 : _GEN_5464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5466 = 9'h18a == _GEN_11439 ? phv_data_394 : _GEN_5465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5467 = 9'h18b == _GEN_11439 ? phv_data_395 : _GEN_5466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5468 = 9'h18c == _GEN_11439 ? phv_data_396 : _GEN_5467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5469 = 9'h18d == _GEN_11439 ? phv_data_397 : _GEN_5468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5470 = 9'h18e == _GEN_11439 ? phv_data_398 : _GEN_5469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5471 = 9'h18f == _GEN_11439 ? phv_data_399 : _GEN_5470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5472 = 9'h190 == _GEN_11439 ? phv_data_400 : _GEN_5471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5473 = 9'h191 == _GEN_11439 ? phv_data_401 : _GEN_5472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5474 = 9'h192 == _GEN_11439 ? phv_data_402 : _GEN_5473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5475 = 9'h193 == _GEN_11439 ? phv_data_403 : _GEN_5474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5476 = 9'h194 == _GEN_11439 ? phv_data_404 : _GEN_5475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5477 = 9'h195 == _GEN_11439 ? phv_data_405 : _GEN_5476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5478 = 9'h196 == _GEN_11439 ? phv_data_406 : _GEN_5477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5479 = 9'h197 == _GEN_11439 ? phv_data_407 : _GEN_5478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5480 = 9'h198 == _GEN_11439 ? phv_data_408 : _GEN_5479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5481 = 9'h199 == _GEN_11439 ? phv_data_409 : _GEN_5480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5482 = 9'h19a == _GEN_11439 ? phv_data_410 : _GEN_5481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5483 = 9'h19b == _GEN_11439 ? phv_data_411 : _GEN_5482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5484 = 9'h19c == _GEN_11439 ? phv_data_412 : _GEN_5483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5485 = 9'h19d == _GEN_11439 ? phv_data_413 : _GEN_5484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5486 = 9'h19e == _GEN_11439 ? phv_data_414 : _GEN_5485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5487 = 9'h19f == _GEN_11439 ? phv_data_415 : _GEN_5486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5488 = 9'h1a0 == _GEN_11439 ? phv_data_416 : _GEN_5487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5489 = 9'h1a1 == _GEN_11439 ? phv_data_417 : _GEN_5488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5490 = 9'h1a2 == _GEN_11439 ? phv_data_418 : _GEN_5489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5491 = 9'h1a3 == _GEN_11439 ? phv_data_419 : _GEN_5490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5492 = 9'h1a4 == _GEN_11439 ? phv_data_420 : _GEN_5491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5493 = 9'h1a5 == _GEN_11439 ? phv_data_421 : _GEN_5492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5494 = 9'h1a6 == _GEN_11439 ? phv_data_422 : _GEN_5493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5495 = 9'h1a7 == _GEN_11439 ? phv_data_423 : _GEN_5494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5496 = 9'h1a8 == _GEN_11439 ? phv_data_424 : _GEN_5495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5497 = 9'h1a9 == _GEN_11439 ? phv_data_425 : _GEN_5496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5498 = 9'h1aa == _GEN_11439 ? phv_data_426 : _GEN_5497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5499 = 9'h1ab == _GEN_11439 ? phv_data_427 : _GEN_5498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5500 = 9'h1ac == _GEN_11439 ? phv_data_428 : _GEN_5499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5501 = 9'h1ad == _GEN_11439 ? phv_data_429 : _GEN_5500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5502 = 9'h1ae == _GEN_11439 ? phv_data_430 : _GEN_5501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5503 = 9'h1af == _GEN_11439 ? phv_data_431 : _GEN_5502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5504 = 9'h1b0 == _GEN_11439 ? phv_data_432 : _GEN_5503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5505 = 9'h1b1 == _GEN_11439 ? phv_data_433 : _GEN_5504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5506 = 9'h1b2 == _GEN_11439 ? phv_data_434 : _GEN_5505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5507 = 9'h1b3 == _GEN_11439 ? phv_data_435 : _GEN_5506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5508 = 9'h1b4 == _GEN_11439 ? phv_data_436 : _GEN_5507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5509 = 9'h1b5 == _GEN_11439 ? phv_data_437 : _GEN_5508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5510 = 9'h1b6 == _GEN_11439 ? phv_data_438 : _GEN_5509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5511 = 9'h1b7 == _GEN_11439 ? phv_data_439 : _GEN_5510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5512 = 9'h1b8 == _GEN_11439 ? phv_data_440 : _GEN_5511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5513 = 9'h1b9 == _GEN_11439 ? phv_data_441 : _GEN_5512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5514 = 9'h1ba == _GEN_11439 ? phv_data_442 : _GEN_5513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5515 = 9'h1bb == _GEN_11439 ? phv_data_443 : _GEN_5514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5516 = 9'h1bc == _GEN_11439 ? phv_data_444 : _GEN_5515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5517 = 9'h1bd == _GEN_11439 ? phv_data_445 : _GEN_5516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5518 = 9'h1be == _GEN_11439 ? phv_data_446 : _GEN_5517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5519 = 9'h1bf == _GEN_11439 ? phv_data_447 : _GEN_5518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5520 = 9'h1c0 == _GEN_11439 ? phv_data_448 : _GEN_5519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5521 = 9'h1c1 == _GEN_11439 ? phv_data_449 : _GEN_5520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5522 = 9'h1c2 == _GEN_11439 ? phv_data_450 : _GEN_5521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5523 = 9'h1c3 == _GEN_11439 ? phv_data_451 : _GEN_5522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5524 = 9'h1c4 == _GEN_11439 ? phv_data_452 : _GEN_5523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5525 = 9'h1c5 == _GEN_11439 ? phv_data_453 : _GEN_5524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5526 = 9'h1c6 == _GEN_11439 ? phv_data_454 : _GEN_5525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5527 = 9'h1c7 == _GEN_11439 ? phv_data_455 : _GEN_5526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5528 = 9'h1c8 == _GEN_11439 ? phv_data_456 : _GEN_5527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5529 = 9'h1c9 == _GEN_11439 ? phv_data_457 : _GEN_5528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5530 = 9'h1ca == _GEN_11439 ? phv_data_458 : _GEN_5529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5531 = 9'h1cb == _GEN_11439 ? phv_data_459 : _GEN_5530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5532 = 9'h1cc == _GEN_11439 ? phv_data_460 : _GEN_5531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5533 = 9'h1cd == _GEN_11439 ? phv_data_461 : _GEN_5532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5534 = 9'h1ce == _GEN_11439 ? phv_data_462 : _GEN_5533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5535 = 9'h1cf == _GEN_11439 ? phv_data_463 : _GEN_5534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5536 = 9'h1d0 == _GEN_11439 ? phv_data_464 : _GEN_5535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5537 = 9'h1d1 == _GEN_11439 ? phv_data_465 : _GEN_5536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5538 = 9'h1d2 == _GEN_11439 ? phv_data_466 : _GEN_5537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5539 = 9'h1d3 == _GEN_11439 ? phv_data_467 : _GEN_5538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5540 = 9'h1d4 == _GEN_11439 ? phv_data_468 : _GEN_5539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5541 = 9'h1d5 == _GEN_11439 ? phv_data_469 : _GEN_5540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5542 = 9'h1d6 == _GEN_11439 ? phv_data_470 : _GEN_5541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5543 = 9'h1d7 == _GEN_11439 ? phv_data_471 : _GEN_5542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5544 = 9'h1d8 == _GEN_11439 ? phv_data_472 : _GEN_5543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5545 = 9'h1d9 == _GEN_11439 ? phv_data_473 : _GEN_5544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5546 = 9'h1da == _GEN_11439 ? phv_data_474 : _GEN_5545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5547 = 9'h1db == _GEN_11439 ? phv_data_475 : _GEN_5546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5548 = 9'h1dc == _GEN_11439 ? phv_data_476 : _GEN_5547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5549 = 9'h1dd == _GEN_11439 ? phv_data_477 : _GEN_5548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5550 = 9'h1de == _GEN_11439 ? phv_data_478 : _GEN_5549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5551 = 9'h1df == _GEN_11439 ? phv_data_479 : _GEN_5550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5552 = 9'h1e0 == _GEN_11439 ? phv_data_480 : _GEN_5551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5553 = 9'h1e1 == _GEN_11439 ? phv_data_481 : _GEN_5552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5554 = 9'h1e2 == _GEN_11439 ? phv_data_482 : _GEN_5553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5555 = 9'h1e3 == _GEN_11439 ? phv_data_483 : _GEN_5554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5556 = 9'h1e4 == _GEN_11439 ? phv_data_484 : _GEN_5555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5557 = 9'h1e5 == _GEN_11439 ? phv_data_485 : _GEN_5556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5558 = 9'h1e6 == _GEN_11439 ? phv_data_486 : _GEN_5557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5559 = 9'h1e7 == _GEN_11439 ? phv_data_487 : _GEN_5558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5560 = 9'h1e8 == _GEN_11439 ? phv_data_488 : _GEN_5559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5561 = 9'h1e9 == _GEN_11439 ? phv_data_489 : _GEN_5560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5562 = 9'h1ea == _GEN_11439 ? phv_data_490 : _GEN_5561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5563 = 9'h1eb == _GEN_11439 ? phv_data_491 : _GEN_5562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5564 = 9'h1ec == _GEN_11439 ? phv_data_492 : _GEN_5563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5565 = 9'h1ed == _GEN_11439 ? phv_data_493 : _GEN_5564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5566 = 9'h1ee == _GEN_11439 ? phv_data_494 : _GEN_5565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5567 = 9'h1ef == _GEN_11439 ? phv_data_495 : _GEN_5566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5568 = 9'h1f0 == _GEN_11439 ? phv_data_496 : _GEN_5567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5569 = 9'h1f1 == _GEN_11439 ? phv_data_497 : _GEN_5568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5570 = 9'h1f2 == _GEN_11439 ? phv_data_498 : _GEN_5569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5571 = 9'h1f3 == _GEN_11439 ? phv_data_499 : _GEN_5570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5572 = 9'h1f4 == _GEN_11439 ? phv_data_500 : _GEN_5571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5573 = 9'h1f5 == _GEN_11439 ? phv_data_501 : _GEN_5572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5574 = 9'h1f6 == _GEN_11439 ? phv_data_502 : _GEN_5573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5575 = 9'h1f7 == _GEN_11439 ? phv_data_503 : _GEN_5574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5576 = 9'h1f8 == _GEN_11439 ? phv_data_504 : _GEN_5575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5577 = 9'h1f9 == _GEN_11439 ? phv_data_505 : _GEN_5576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5578 = 9'h1fa == _GEN_11439 ? phv_data_506 : _GEN_5577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5579 = 9'h1fb == _GEN_11439 ? phv_data_507 : _GEN_5578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5580 = 9'h1fc == _GEN_11439 ? phv_data_508 : _GEN_5579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5581 = 9'h1fd == _GEN_11439 ? phv_data_509 : _GEN_5580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5582 = 9'h1fe == _GEN_11439 ? phv_data_510 : _GEN_5581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_2 = 9'h1ff == _GEN_11439 ? phv_data_511 : _GEN_5582; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_2_2 = 2'h1 >= offset_2[1:0] & (2'h1 < ending_2 | ending_2 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_10 = {total_offset_hi_2,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_5585 = 8'h1 == total_offset_10 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5586 = 8'h2 == total_offset_10 ? phv_data_2 : _GEN_5585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5587 = 8'h3 == total_offset_10 ? phv_data_3 : _GEN_5586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5588 = 8'h4 == total_offset_10 ? phv_data_4 : _GEN_5587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5589 = 8'h5 == total_offset_10 ? phv_data_5 : _GEN_5588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5590 = 8'h6 == total_offset_10 ? phv_data_6 : _GEN_5589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5591 = 8'h7 == total_offset_10 ? phv_data_7 : _GEN_5590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5592 = 8'h8 == total_offset_10 ? phv_data_8 : _GEN_5591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5593 = 8'h9 == total_offset_10 ? phv_data_9 : _GEN_5592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5594 = 8'ha == total_offset_10 ? phv_data_10 : _GEN_5593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5595 = 8'hb == total_offset_10 ? phv_data_11 : _GEN_5594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5596 = 8'hc == total_offset_10 ? phv_data_12 : _GEN_5595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5597 = 8'hd == total_offset_10 ? phv_data_13 : _GEN_5596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5598 = 8'he == total_offset_10 ? phv_data_14 : _GEN_5597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5599 = 8'hf == total_offset_10 ? phv_data_15 : _GEN_5598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5600 = 8'h10 == total_offset_10 ? phv_data_16 : _GEN_5599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5601 = 8'h11 == total_offset_10 ? phv_data_17 : _GEN_5600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5602 = 8'h12 == total_offset_10 ? phv_data_18 : _GEN_5601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5603 = 8'h13 == total_offset_10 ? phv_data_19 : _GEN_5602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5604 = 8'h14 == total_offset_10 ? phv_data_20 : _GEN_5603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5605 = 8'h15 == total_offset_10 ? phv_data_21 : _GEN_5604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5606 = 8'h16 == total_offset_10 ? phv_data_22 : _GEN_5605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5607 = 8'h17 == total_offset_10 ? phv_data_23 : _GEN_5606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5608 = 8'h18 == total_offset_10 ? phv_data_24 : _GEN_5607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5609 = 8'h19 == total_offset_10 ? phv_data_25 : _GEN_5608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5610 = 8'h1a == total_offset_10 ? phv_data_26 : _GEN_5609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5611 = 8'h1b == total_offset_10 ? phv_data_27 : _GEN_5610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5612 = 8'h1c == total_offset_10 ? phv_data_28 : _GEN_5611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5613 = 8'h1d == total_offset_10 ? phv_data_29 : _GEN_5612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5614 = 8'h1e == total_offset_10 ? phv_data_30 : _GEN_5613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5615 = 8'h1f == total_offset_10 ? phv_data_31 : _GEN_5614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5616 = 8'h20 == total_offset_10 ? phv_data_32 : _GEN_5615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5617 = 8'h21 == total_offset_10 ? phv_data_33 : _GEN_5616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5618 = 8'h22 == total_offset_10 ? phv_data_34 : _GEN_5617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5619 = 8'h23 == total_offset_10 ? phv_data_35 : _GEN_5618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5620 = 8'h24 == total_offset_10 ? phv_data_36 : _GEN_5619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5621 = 8'h25 == total_offset_10 ? phv_data_37 : _GEN_5620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5622 = 8'h26 == total_offset_10 ? phv_data_38 : _GEN_5621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5623 = 8'h27 == total_offset_10 ? phv_data_39 : _GEN_5622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5624 = 8'h28 == total_offset_10 ? phv_data_40 : _GEN_5623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5625 = 8'h29 == total_offset_10 ? phv_data_41 : _GEN_5624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5626 = 8'h2a == total_offset_10 ? phv_data_42 : _GEN_5625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5627 = 8'h2b == total_offset_10 ? phv_data_43 : _GEN_5626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5628 = 8'h2c == total_offset_10 ? phv_data_44 : _GEN_5627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5629 = 8'h2d == total_offset_10 ? phv_data_45 : _GEN_5628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5630 = 8'h2e == total_offset_10 ? phv_data_46 : _GEN_5629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5631 = 8'h2f == total_offset_10 ? phv_data_47 : _GEN_5630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5632 = 8'h30 == total_offset_10 ? phv_data_48 : _GEN_5631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5633 = 8'h31 == total_offset_10 ? phv_data_49 : _GEN_5632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5634 = 8'h32 == total_offset_10 ? phv_data_50 : _GEN_5633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5635 = 8'h33 == total_offset_10 ? phv_data_51 : _GEN_5634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5636 = 8'h34 == total_offset_10 ? phv_data_52 : _GEN_5635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5637 = 8'h35 == total_offset_10 ? phv_data_53 : _GEN_5636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5638 = 8'h36 == total_offset_10 ? phv_data_54 : _GEN_5637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5639 = 8'h37 == total_offset_10 ? phv_data_55 : _GEN_5638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5640 = 8'h38 == total_offset_10 ? phv_data_56 : _GEN_5639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5641 = 8'h39 == total_offset_10 ? phv_data_57 : _GEN_5640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5642 = 8'h3a == total_offset_10 ? phv_data_58 : _GEN_5641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5643 = 8'h3b == total_offset_10 ? phv_data_59 : _GEN_5642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5644 = 8'h3c == total_offset_10 ? phv_data_60 : _GEN_5643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5645 = 8'h3d == total_offset_10 ? phv_data_61 : _GEN_5644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5646 = 8'h3e == total_offset_10 ? phv_data_62 : _GEN_5645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5647 = 8'h3f == total_offset_10 ? phv_data_63 : _GEN_5646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5648 = 8'h40 == total_offset_10 ? phv_data_64 : _GEN_5647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5649 = 8'h41 == total_offset_10 ? phv_data_65 : _GEN_5648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5650 = 8'h42 == total_offset_10 ? phv_data_66 : _GEN_5649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5651 = 8'h43 == total_offset_10 ? phv_data_67 : _GEN_5650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5652 = 8'h44 == total_offset_10 ? phv_data_68 : _GEN_5651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5653 = 8'h45 == total_offset_10 ? phv_data_69 : _GEN_5652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5654 = 8'h46 == total_offset_10 ? phv_data_70 : _GEN_5653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5655 = 8'h47 == total_offset_10 ? phv_data_71 : _GEN_5654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5656 = 8'h48 == total_offset_10 ? phv_data_72 : _GEN_5655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5657 = 8'h49 == total_offset_10 ? phv_data_73 : _GEN_5656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5658 = 8'h4a == total_offset_10 ? phv_data_74 : _GEN_5657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5659 = 8'h4b == total_offset_10 ? phv_data_75 : _GEN_5658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5660 = 8'h4c == total_offset_10 ? phv_data_76 : _GEN_5659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5661 = 8'h4d == total_offset_10 ? phv_data_77 : _GEN_5660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5662 = 8'h4e == total_offset_10 ? phv_data_78 : _GEN_5661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5663 = 8'h4f == total_offset_10 ? phv_data_79 : _GEN_5662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5664 = 8'h50 == total_offset_10 ? phv_data_80 : _GEN_5663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5665 = 8'h51 == total_offset_10 ? phv_data_81 : _GEN_5664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5666 = 8'h52 == total_offset_10 ? phv_data_82 : _GEN_5665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5667 = 8'h53 == total_offset_10 ? phv_data_83 : _GEN_5666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5668 = 8'h54 == total_offset_10 ? phv_data_84 : _GEN_5667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5669 = 8'h55 == total_offset_10 ? phv_data_85 : _GEN_5668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5670 = 8'h56 == total_offset_10 ? phv_data_86 : _GEN_5669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5671 = 8'h57 == total_offset_10 ? phv_data_87 : _GEN_5670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5672 = 8'h58 == total_offset_10 ? phv_data_88 : _GEN_5671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5673 = 8'h59 == total_offset_10 ? phv_data_89 : _GEN_5672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5674 = 8'h5a == total_offset_10 ? phv_data_90 : _GEN_5673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5675 = 8'h5b == total_offset_10 ? phv_data_91 : _GEN_5674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5676 = 8'h5c == total_offset_10 ? phv_data_92 : _GEN_5675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5677 = 8'h5d == total_offset_10 ? phv_data_93 : _GEN_5676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5678 = 8'h5e == total_offset_10 ? phv_data_94 : _GEN_5677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5679 = 8'h5f == total_offset_10 ? phv_data_95 : _GEN_5678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5680 = 8'h60 == total_offset_10 ? phv_data_96 : _GEN_5679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5681 = 8'h61 == total_offset_10 ? phv_data_97 : _GEN_5680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5682 = 8'h62 == total_offset_10 ? phv_data_98 : _GEN_5681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5683 = 8'h63 == total_offset_10 ? phv_data_99 : _GEN_5682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5684 = 8'h64 == total_offset_10 ? phv_data_100 : _GEN_5683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5685 = 8'h65 == total_offset_10 ? phv_data_101 : _GEN_5684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5686 = 8'h66 == total_offset_10 ? phv_data_102 : _GEN_5685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5687 = 8'h67 == total_offset_10 ? phv_data_103 : _GEN_5686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5688 = 8'h68 == total_offset_10 ? phv_data_104 : _GEN_5687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5689 = 8'h69 == total_offset_10 ? phv_data_105 : _GEN_5688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5690 = 8'h6a == total_offset_10 ? phv_data_106 : _GEN_5689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5691 = 8'h6b == total_offset_10 ? phv_data_107 : _GEN_5690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5692 = 8'h6c == total_offset_10 ? phv_data_108 : _GEN_5691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5693 = 8'h6d == total_offset_10 ? phv_data_109 : _GEN_5692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5694 = 8'h6e == total_offset_10 ? phv_data_110 : _GEN_5693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5695 = 8'h6f == total_offset_10 ? phv_data_111 : _GEN_5694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5696 = 8'h70 == total_offset_10 ? phv_data_112 : _GEN_5695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5697 = 8'h71 == total_offset_10 ? phv_data_113 : _GEN_5696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5698 = 8'h72 == total_offset_10 ? phv_data_114 : _GEN_5697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5699 = 8'h73 == total_offset_10 ? phv_data_115 : _GEN_5698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5700 = 8'h74 == total_offset_10 ? phv_data_116 : _GEN_5699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5701 = 8'h75 == total_offset_10 ? phv_data_117 : _GEN_5700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5702 = 8'h76 == total_offset_10 ? phv_data_118 : _GEN_5701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5703 = 8'h77 == total_offset_10 ? phv_data_119 : _GEN_5702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5704 = 8'h78 == total_offset_10 ? phv_data_120 : _GEN_5703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5705 = 8'h79 == total_offset_10 ? phv_data_121 : _GEN_5704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5706 = 8'h7a == total_offset_10 ? phv_data_122 : _GEN_5705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5707 = 8'h7b == total_offset_10 ? phv_data_123 : _GEN_5706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5708 = 8'h7c == total_offset_10 ? phv_data_124 : _GEN_5707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5709 = 8'h7d == total_offset_10 ? phv_data_125 : _GEN_5708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5710 = 8'h7e == total_offset_10 ? phv_data_126 : _GEN_5709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5711 = 8'h7f == total_offset_10 ? phv_data_127 : _GEN_5710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5712 = 8'h80 == total_offset_10 ? phv_data_128 : _GEN_5711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5713 = 8'h81 == total_offset_10 ? phv_data_129 : _GEN_5712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5714 = 8'h82 == total_offset_10 ? phv_data_130 : _GEN_5713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5715 = 8'h83 == total_offset_10 ? phv_data_131 : _GEN_5714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5716 = 8'h84 == total_offset_10 ? phv_data_132 : _GEN_5715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5717 = 8'h85 == total_offset_10 ? phv_data_133 : _GEN_5716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5718 = 8'h86 == total_offset_10 ? phv_data_134 : _GEN_5717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5719 = 8'h87 == total_offset_10 ? phv_data_135 : _GEN_5718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5720 = 8'h88 == total_offset_10 ? phv_data_136 : _GEN_5719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5721 = 8'h89 == total_offset_10 ? phv_data_137 : _GEN_5720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5722 = 8'h8a == total_offset_10 ? phv_data_138 : _GEN_5721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5723 = 8'h8b == total_offset_10 ? phv_data_139 : _GEN_5722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5724 = 8'h8c == total_offset_10 ? phv_data_140 : _GEN_5723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5725 = 8'h8d == total_offset_10 ? phv_data_141 : _GEN_5724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5726 = 8'h8e == total_offset_10 ? phv_data_142 : _GEN_5725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5727 = 8'h8f == total_offset_10 ? phv_data_143 : _GEN_5726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5728 = 8'h90 == total_offset_10 ? phv_data_144 : _GEN_5727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5729 = 8'h91 == total_offset_10 ? phv_data_145 : _GEN_5728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5730 = 8'h92 == total_offset_10 ? phv_data_146 : _GEN_5729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5731 = 8'h93 == total_offset_10 ? phv_data_147 : _GEN_5730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5732 = 8'h94 == total_offset_10 ? phv_data_148 : _GEN_5731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5733 = 8'h95 == total_offset_10 ? phv_data_149 : _GEN_5732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5734 = 8'h96 == total_offset_10 ? phv_data_150 : _GEN_5733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5735 = 8'h97 == total_offset_10 ? phv_data_151 : _GEN_5734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5736 = 8'h98 == total_offset_10 ? phv_data_152 : _GEN_5735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5737 = 8'h99 == total_offset_10 ? phv_data_153 : _GEN_5736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5738 = 8'h9a == total_offset_10 ? phv_data_154 : _GEN_5737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5739 = 8'h9b == total_offset_10 ? phv_data_155 : _GEN_5738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5740 = 8'h9c == total_offset_10 ? phv_data_156 : _GEN_5739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5741 = 8'h9d == total_offset_10 ? phv_data_157 : _GEN_5740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5742 = 8'h9e == total_offset_10 ? phv_data_158 : _GEN_5741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5743 = 8'h9f == total_offset_10 ? phv_data_159 : _GEN_5742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5744 = 8'ha0 == total_offset_10 ? phv_data_160 : _GEN_5743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5745 = 8'ha1 == total_offset_10 ? phv_data_161 : _GEN_5744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5746 = 8'ha2 == total_offset_10 ? phv_data_162 : _GEN_5745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5747 = 8'ha3 == total_offset_10 ? phv_data_163 : _GEN_5746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5748 = 8'ha4 == total_offset_10 ? phv_data_164 : _GEN_5747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5749 = 8'ha5 == total_offset_10 ? phv_data_165 : _GEN_5748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5750 = 8'ha6 == total_offset_10 ? phv_data_166 : _GEN_5749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5751 = 8'ha7 == total_offset_10 ? phv_data_167 : _GEN_5750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5752 = 8'ha8 == total_offset_10 ? phv_data_168 : _GEN_5751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5753 = 8'ha9 == total_offset_10 ? phv_data_169 : _GEN_5752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5754 = 8'haa == total_offset_10 ? phv_data_170 : _GEN_5753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5755 = 8'hab == total_offset_10 ? phv_data_171 : _GEN_5754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5756 = 8'hac == total_offset_10 ? phv_data_172 : _GEN_5755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5757 = 8'had == total_offset_10 ? phv_data_173 : _GEN_5756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5758 = 8'hae == total_offset_10 ? phv_data_174 : _GEN_5757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5759 = 8'haf == total_offset_10 ? phv_data_175 : _GEN_5758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5760 = 8'hb0 == total_offset_10 ? phv_data_176 : _GEN_5759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5761 = 8'hb1 == total_offset_10 ? phv_data_177 : _GEN_5760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5762 = 8'hb2 == total_offset_10 ? phv_data_178 : _GEN_5761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5763 = 8'hb3 == total_offset_10 ? phv_data_179 : _GEN_5762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5764 = 8'hb4 == total_offset_10 ? phv_data_180 : _GEN_5763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5765 = 8'hb5 == total_offset_10 ? phv_data_181 : _GEN_5764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5766 = 8'hb6 == total_offset_10 ? phv_data_182 : _GEN_5765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5767 = 8'hb7 == total_offset_10 ? phv_data_183 : _GEN_5766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5768 = 8'hb8 == total_offset_10 ? phv_data_184 : _GEN_5767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5769 = 8'hb9 == total_offset_10 ? phv_data_185 : _GEN_5768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5770 = 8'hba == total_offset_10 ? phv_data_186 : _GEN_5769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5771 = 8'hbb == total_offset_10 ? phv_data_187 : _GEN_5770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5772 = 8'hbc == total_offset_10 ? phv_data_188 : _GEN_5771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5773 = 8'hbd == total_offset_10 ? phv_data_189 : _GEN_5772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5774 = 8'hbe == total_offset_10 ? phv_data_190 : _GEN_5773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5775 = 8'hbf == total_offset_10 ? phv_data_191 : _GEN_5774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5776 = 8'hc0 == total_offset_10 ? phv_data_192 : _GEN_5775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5777 = 8'hc1 == total_offset_10 ? phv_data_193 : _GEN_5776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5778 = 8'hc2 == total_offset_10 ? phv_data_194 : _GEN_5777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5779 = 8'hc3 == total_offset_10 ? phv_data_195 : _GEN_5778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5780 = 8'hc4 == total_offset_10 ? phv_data_196 : _GEN_5779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5781 = 8'hc5 == total_offset_10 ? phv_data_197 : _GEN_5780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5782 = 8'hc6 == total_offset_10 ? phv_data_198 : _GEN_5781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5783 = 8'hc7 == total_offset_10 ? phv_data_199 : _GEN_5782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5784 = 8'hc8 == total_offset_10 ? phv_data_200 : _GEN_5783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5785 = 8'hc9 == total_offset_10 ? phv_data_201 : _GEN_5784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5786 = 8'hca == total_offset_10 ? phv_data_202 : _GEN_5785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5787 = 8'hcb == total_offset_10 ? phv_data_203 : _GEN_5786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5788 = 8'hcc == total_offset_10 ? phv_data_204 : _GEN_5787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5789 = 8'hcd == total_offset_10 ? phv_data_205 : _GEN_5788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5790 = 8'hce == total_offset_10 ? phv_data_206 : _GEN_5789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5791 = 8'hcf == total_offset_10 ? phv_data_207 : _GEN_5790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5792 = 8'hd0 == total_offset_10 ? phv_data_208 : _GEN_5791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5793 = 8'hd1 == total_offset_10 ? phv_data_209 : _GEN_5792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5794 = 8'hd2 == total_offset_10 ? phv_data_210 : _GEN_5793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5795 = 8'hd3 == total_offset_10 ? phv_data_211 : _GEN_5794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5796 = 8'hd4 == total_offset_10 ? phv_data_212 : _GEN_5795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5797 = 8'hd5 == total_offset_10 ? phv_data_213 : _GEN_5796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5798 = 8'hd6 == total_offset_10 ? phv_data_214 : _GEN_5797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5799 = 8'hd7 == total_offset_10 ? phv_data_215 : _GEN_5798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5800 = 8'hd8 == total_offset_10 ? phv_data_216 : _GEN_5799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5801 = 8'hd9 == total_offset_10 ? phv_data_217 : _GEN_5800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5802 = 8'hda == total_offset_10 ? phv_data_218 : _GEN_5801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5803 = 8'hdb == total_offset_10 ? phv_data_219 : _GEN_5802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5804 = 8'hdc == total_offset_10 ? phv_data_220 : _GEN_5803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5805 = 8'hdd == total_offset_10 ? phv_data_221 : _GEN_5804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5806 = 8'hde == total_offset_10 ? phv_data_222 : _GEN_5805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5807 = 8'hdf == total_offset_10 ? phv_data_223 : _GEN_5806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5808 = 8'he0 == total_offset_10 ? phv_data_224 : _GEN_5807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5809 = 8'he1 == total_offset_10 ? phv_data_225 : _GEN_5808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5810 = 8'he2 == total_offset_10 ? phv_data_226 : _GEN_5809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5811 = 8'he3 == total_offset_10 ? phv_data_227 : _GEN_5810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5812 = 8'he4 == total_offset_10 ? phv_data_228 : _GEN_5811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5813 = 8'he5 == total_offset_10 ? phv_data_229 : _GEN_5812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5814 = 8'he6 == total_offset_10 ? phv_data_230 : _GEN_5813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5815 = 8'he7 == total_offset_10 ? phv_data_231 : _GEN_5814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5816 = 8'he8 == total_offset_10 ? phv_data_232 : _GEN_5815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5817 = 8'he9 == total_offset_10 ? phv_data_233 : _GEN_5816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5818 = 8'hea == total_offset_10 ? phv_data_234 : _GEN_5817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5819 = 8'heb == total_offset_10 ? phv_data_235 : _GEN_5818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5820 = 8'hec == total_offset_10 ? phv_data_236 : _GEN_5819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5821 = 8'hed == total_offset_10 ? phv_data_237 : _GEN_5820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5822 = 8'hee == total_offset_10 ? phv_data_238 : _GEN_5821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5823 = 8'hef == total_offset_10 ? phv_data_239 : _GEN_5822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5824 = 8'hf0 == total_offset_10 ? phv_data_240 : _GEN_5823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5825 = 8'hf1 == total_offset_10 ? phv_data_241 : _GEN_5824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5826 = 8'hf2 == total_offset_10 ? phv_data_242 : _GEN_5825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5827 = 8'hf3 == total_offset_10 ? phv_data_243 : _GEN_5826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5828 = 8'hf4 == total_offset_10 ? phv_data_244 : _GEN_5827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5829 = 8'hf5 == total_offset_10 ? phv_data_245 : _GEN_5828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5830 = 8'hf6 == total_offset_10 ? phv_data_246 : _GEN_5829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5831 = 8'hf7 == total_offset_10 ? phv_data_247 : _GEN_5830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5832 = 8'hf8 == total_offset_10 ? phv_data_248 : _GEN_5831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5833 = 8'hf9 == total_offset_10 ? phv_data_249 : _GEN_5832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5834 = 8'hfa == total_offset_10 ? phv_data_250 : _GEN_5833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5835 = 8'hfb == total_offset_10 ? phv_data_251 : _GEN_5834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5836 = 8'hfc == total_offset_10 ? phv_data_252 : _GEN_5835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5837 = 8'hfd == total_offset_10 ? phv_data_253 : _GEN_5836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5838 = 8'hfe == total_offset_10 ? phv_data_254 : _GEN_5837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5839 = 8'hff == total_offset_10 ? phv_data_255 : _GEN_5838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_11695 = {{1'd0}, total_offset_10}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5840 = 9'h100 == _GEN_11695 ? phv_data_256 : _GEN_5839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5841 = 9'h101 == _GEN_11695 ? phv_data_257 : _GEN_5840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5842 = 9'h102 == _GEN_11695 ? phv_data_258 : _GEN_5841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5843 = 9'h103 == _GEN_11695 ? phv_data_259 : _GEN_5842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5844 = 9'h104 == _GEN_11695 ? phv_data_260 : _GEN_5843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5845 = 9'h105 == _GEN_11695 ? phv_data_261 : _GEN_5844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5846 = 9'h106 == _GEN_11695 ? phv_data_262 : _GEN_5845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5847 = 9'h107 == _GEN_11695 ? phv_data_263 : _GEN_5846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5848 = 9'h108 == _GEN_11695 ? phv_data_264 : _GEN_5847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5849 = 9'h109 == _GEN_11695 ? phv_data_265 : _GEN_5848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5850 = 9'h10a == _GEN_11695 ? phv_data_266 : _GEN_5849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5851 = 9'h10b == _GEN_11695 ? phv_data_267 : _GEN_5850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5852 = 9'h10c == _GEN_11695 ? phv_data_268 : _GEN_5851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5853 = 9'h10d == _GEN_11695 ? phv_data_269 : _GEN_5852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5854 = 9'h10e == _GEN_11695 ? phv_data_270 : _GEN_5853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5855 = 9'h10f == _GEN_11695 ? phv_data_271 : _GEN_5854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5856 = 9'h110 == _GEN_11695 ? phv_data_272 : _GEN_5855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5857 = 9'h111 == _GEN_11695 ? phv_data_273 : _GEN_5856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5858 = 9'h112 == _GEN_11695 ? phv_data_274 : _GEN_5857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5859 = 9'h113 == _GEN_11695 ? phv_data_275 : _GEN_5858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5860 = 9'h114 == _GEN_11695 ? phv_data_276 : _GEN_5859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5861 = 9'h115 == _GEN_11695 ? phv_data_277 : _GEN_5860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5862 = 9'h116 == _GEN_11695 ? phv_data_278 : _GEN_5861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5863 = 9'h117 == _GEN_11695 ? phv_data_279 : _GEN_5862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5864 = 9'h118 == _GEN_11695 ? phv_data_280 : _GEN_5863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5865 = 9'h119 == _GEN_11695 ? phv_data_281 : _GEN_5864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5866 = 9'h11a == _GEN_11695 ? phv_data_282 : _GEN_5865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5867 = 9'h11b == _GEN_11695 ? phv_data_283 : _GEN_5866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5868 = 9'h11c == _GEN_11695 ? phv_data_284 : _GEN_5867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5869 = 9'h11d == _GEN_11695 ? phv_data_285 : _GEN_5868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5870 = 9'h11e == _GEN_11695 ? phv_data_286 : _GEN_5869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5871 = 9'h11f == _GEN_11695 ? phv_data_287 : _GEN_5870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5872 = 9'h120 == _GEN_11695 ? phv_data_288 : _GEN_5871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5873 = 9'h121 == _GEN_11695 ? phv_data_289 : _GEN_5872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5874 = 9'h122 == _GEN_11695 ? phv_data_290 : _GEN_5873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5875 = 9'h123 == _GEN_11695 ? phv_data_291 : _GEN_5874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5876 = 9'h124 == _GEN_11695 ? phv_data_292 : _GEN_5875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5877 = 9'h125 == _GEN_11695 ? phv_data_293 : _GEN_5876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5878 = 9'h126 == _GEN_11695 ? phv_data_294 : _GEN_5877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5879 = 9'h127 == _GEN_11695 ? phv_data_295 : _GEN_5878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5880 = 9'h128 == _GEN_11695 ? phv_data_296 : _GEN_5879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5881 = 9'h129 == _GEN_11695 ? phv_data_297 : _GEN_5880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5882 = 9'h12a == _GEN_11695 ? phv_data_298 : _GEN_5881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5883 = 9'h12b == _GEN_11695 ? phv_data_299 : _GEN_5882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5884 = 9'h12c == _GEN_11695 ? phv_data_300 : _GEN_5883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5885 = 9'h12d == _GEN_11695 ? phv_data_301 : _GEN_5884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5886 = 9'h12e == _GEN_11695 ? phv_data_302 : _GEN_5885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5887 = 9'h12f == _GEN_11695 ? phv_data_303 : _GEN_5886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5888 = 9'h130 == _GEN_11695 ? phv_data_304 : _GEN_5887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5889 = 9'h131 == _GEN_11695 ? phv_data_305 : _GEN_5888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5890 = 9'h132 == _GEN_11695 ? phv_data_306 : _GEN_5889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5891 = 9'h133 == _GEN_11695 ? phv_data_307 : _GEN_5890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5892 = 9'h134 == _GEN_11695 ? phv_data_308 : _GEN_5891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5893 = 9'h135 == _GEN_11695 ? phv_data_309 : _GEN_5892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5894 = 9'h136 == _GEN_11695 ? phv_data_310 : _GEN_5893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5895 = 9'h137 == _GEN_11695 ? phv_data_311 : _GEN_5894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5896 = 9'h138 == _GEN_11695 ? phv_data_312 : _GEN_5895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5897 = 9'h139 == _GEN_11695 ? phv_data_313 : _GEN_5896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5898 = 9'h13a == _GEN_11695 ? phv_data_314 : _GEN_5897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5899 = 9'h13b == _GEN_11695 ? phv_data_315 : _GEN_5898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5900 = 9'h13c == _GEN_11695 ? phv_data_316 : _GEN_5899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5901 = 9'h13d == _GEN_11695 ? phv_data_317 : _GEN_5900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5902 = 9'h13e == _GEN_11695 ? phv_data_318 : _GEN_5901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5903 = 9'h13f == _GEN_11695 ? phv_data_319 : _GEN_5902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5904 = 9'h140 == _GEN_11695 ? phv_data_320 : _GEN_5903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5905 = 9'h141 == _GEN_11695 ? phv_data_321 : _GEN_5904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5906 = 9'h142 == _GEN_11695 ? phv_data_322 : _GEN_5905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5907 = 9'h143 == _GEN_11695 ? phv_data_323 : _GEN_5906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5908 = 9'h144 == _GEN_11695 ? phv_data_324 : _GEN_5907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5909 = 9'h145 == _GEN_11695 ? phv_data_325 : _GEN_5908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5910 = 9'h146 == _GEN_11695 ? phv_data_326 : _GEN_5909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5911 = 9'h147 == _GEN_11695 ? phv_data_327 : _GEN_5910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5912 = 9'h148 == _GEN_11695 ? phv_data_328 : _GEN_5911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5913 = 9'h149 == _GEN_11695 ? phv_data_329 : _GEN_5912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5914 = 9'h14a == _GEN_11695 ? phv_data_330 : _GEN_5913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5915 = 9'h14b == _GEN_11695 ? phv_data_331 : _GEN_5914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5916 = 9'h14c == _GEN_11695 ? phv_data_332 : _GEN_5915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5917 = 9'h14d == _GEN_11695 ? phv_data_333 : _GEN_5916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5918 = 9'h14e == _GEN_11695 ? phv_data_334 : _GEN_5917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5919 = 9'h14f == _GEN_11695 ? phv_data_335 : _GEN_5918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5920 = 9'h150 == _GEN_11695 ? phv_data_336 : _GEN_5919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5921 = 9'h151 == _GEN_11695 ? phv_data_337 : _GEN_5920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5922 = 9'h152 == _GEN_11695 ? phv_data_338 : _GEN_5921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5923 = 9'h153 == _GEN_11695 ? phv_data_339 : _GEN_5922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5924 = 9'h154 == _GEN_11695 ? phv_data_340 : _GEN_5923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5925 = 9'h155 == _GEN_11695 ? phv_data_341 : _GEN_5924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5926 = 9'h156 == _GEN_11695 ? phv_data_342 : _GEN_5925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5927 = 9'h157 == _GEN_11695 ? phv_data_343 : _GEN_5926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5928 = 9'h158 == _GEN_11695 ? phv_data_344 : _GEN_5927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5929 = 9'h159 == _GEN_11695 ? phv_data_345 : _GEN_5928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5930 = 9'h15a == _GEN_11695 ? phv_data_346 : _GEN_5929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5931 = 9'h15b == _GEN_11695 ? phv_data_347 : _GEN_5930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5932 = 9'h15c == _GEN_11695 ? phv_data_348 : _GEN_5931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5933 = 9'h15d == _GEN_11695 ? phv_data_349 : _GEN_5932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5934 = 9'h15e == _GEN_11695 ? phv_data_350 : _GEN_5933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5935 = 9'h15f == _GEN_11695 ? phv_data_351 : _GEN_5934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5936 = 9'h160 == _GEN_11695 ? phv_data_352 : _GEN_5935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5937 = 9'h161 == _GEN_11695 ? phv_data_353 : _GEN_5936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5938 = 9'h162 == _GEN_11695 ? phv_data_354 : _GEN_5937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5939 = 9'h163 == _GEN_11695 ? phv_data_355 : _GEN_5938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5940 = 9'h164 == _GEN_11695 ? phv_data_356 : _GEN_5939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5941 = 9'h165 == _GEN_11695 ? phv_data_357 : _GEN_5940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5942 = 9'h166 == _GEN_11695 ? phv_data_358 : _GEN_5941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5943 = 9'h167 == _GEN_11695 ? phv_data_359 : _GEN_5942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5944 = 9'h168 == _GEN_11695 ? phv_data_360 : _GEN_5943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5945 = 9'h169 == _GEN_11695 ? phv_data_361 : _GEN_5944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5946 = 9'h16a == _GEN_11695 ? phv_data_362 : _GEN_5945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5947 = 9'h16b == _GEN_11695 ? phv_data_363 : _GEN_5946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5948 = 9'h16c == _GEN_11695 ? phv_data_364 : _GEN_5947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5949 = 9'h16d == _GEN_11695 ? phv_data_365 : _GEN_5948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5950 = 9'h16e == _GEN_11695 ? phv_data_366 : _GEN_5949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5951 = 9'h16f == _GEN_11695 ? phv_data_367 : _GEN_5950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5952 = 9'h170 == _GEN_11695 ? phv_data_368 : _GEN_5951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5953 = 9'h171 == _GEN_11695 ? phv_data_369 : _GEN_5952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5954 = 9'h172 == _GEN_11695 ? phv_data_370 : _GEN_5953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5955 = 9'h173 == _GEN_11695 ? phv_data_371 : _GEN_5954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5956 = 9'h174 == _GEN_11695 ? phv_data_372 : _GEN_5955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5957 = 9'h175 == _GEN_11695 ? phv_data_373 : _GEN_5956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5958 = 9'h176 == _GEN_11695 ? phv_data_374 : _GEN_5957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5959 = 9'h177 == _GEN_11695 ? phv_data_375 : _GEN_5958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5960 = 9'h178 == _GEN_11695 ? phv_data_376 : _GEN_5959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5961 = 9'h179 == _GEN_11695 ? phv_data_377 : _GEN_5960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5962 = 9'h17a == _GEN_11695 ? phv_data_378 : _GEN_5961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5963 = 9'h17b == _GEN_11695 ? phv_data_379 : _GEN_5962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5964 = 9'h17c == _GEN_11695 ? phv_data_380 : _GEN_5963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5965 = 9'h17d == _GEN_11695 ? phv_data_381 : _GEN_5964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5966 = 9'h17e == _GEN_11695 ? phv_data_382 : _GEN_5965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5967 = 9'h17f == _GEN_11695 ? phv_data_383 : _GEN_5966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5968 = 9'h180 == _GEN_11695 ? phv_data_384 : _GEN_5967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5969 = 9'h181 == _GEN_11695 ? phv_data_385 : _GEN_5968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5970 = 9'h182 == _GEN_11695 ? phv_data_386 : _GEN_5969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5971 = 9'h183 == _GEN_11695 ? phv_data_387 : _GEN_5970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5972 = 9'h184 == _GEN_11695 ? phv_data_388 : _GEN_5971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5973 = 9'h185 == _GEN_11695 ? phv_data_389 : _GEN_5972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5974 = 9'h186 == _GEN_11695 ? phv_data_390 : _GEN_5973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5975 = 9'h187 == _GEN_11695 ? phv_data_391 : _GEN_5974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5976 = 9'h188 == _GEN_11695 ? phv_data_392 : _GEN_5975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5977 = 9'h189 == _GEN_11695 ? phv_data_393 : _GEN_5976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5978 = 9'h18a == _GEN_11695 ? phv_data_394 : _GEN_5977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5979 = 9'h18b == _GEN_11695 ? phv_data_395 : _GEN_5978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5980 = 9'h18c == _GEN_11695 ? phv_data_396 : _GEN_5979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5981 = 9'h18d == _GEN_11695 ? phv_data_397 : _GEN_5980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5982 = 9'h18e == _GEN_11695 ? phv_data_398 : _GEN_5981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5983 = 9'h18f == _GEN_11695 ? phv_data_399 : _GEN_5982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5984 = 9'h190 == _GEN_11695 ? phv_data_400 : _GEN_5983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5985 = 9'h191 == _GEN_11695 ? phv_data_401 : _GEN_5984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5986 = 9'h192 == _GEN_11695 ? phv_data_402 : _GEN_5985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5987 = 9'h193 == _GEN_11695 ? phv_data_403 : _GEN_5986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5988 = 9'h194 == _GEN_11695 ? phv_data_404 : _GEN_5987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5989 = 9'h195 == _GEN_11695 ? phv_data_405 : _GEN_5988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5990 = 9'h196 == _GEN_11695 ? phv_data_406 : _GEN_5989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5991 = 9'h197 == _GEN_11695 ? phv_data_407 : _GEN_5990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5992 = 9'h198 == _GEN_11695 ? phv_data_408 : _GEN_5991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5993 = 9'h199 == _GEN_11695 ? phv_data_409 : _GEN_5992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5994 = 9'h19a == _GEN_11695 ? phv_data_410 : _GEN_5993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5995 = 9'h19b == _GEN_11695 ? phv_data_411 : _GEN_5994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5996 = 9'h19c == _GEN_11695 ? phv_data_412 : _GEN_5995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5997 = 9'h19d == _GEN_11695 ? phv_data_413 : _GEN_5996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5998 = 9'h19e == _GEN_11695 ? phv_data_414 : _GEN_5997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_5999 = 9'h19f == _GEN_11695 ? phv_data_415 : _GEN_5998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6000 = 9'h1a0 == _GEN_11695 ? phv_data_416 : _GEN_5999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6001 = 9'h1a1 == _GEN_11695 ? phv_data_417 : _GEN_6000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6002 = 9'h1a2 == _GEN_11695 ? phv_data_418 : _GEN_6001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6003 = 9'h1a3 == _GEN_11695 ? phv_data_419 : _GEN_6002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6004 = 9'h1a4 == _GEN_11695 ? phv_data_420 : _GEN_6003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6005 = 9'h1a5 == _GEN_11695 ? phv_data_421 : _GEN_6004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6006 = 9'h1a6 == _GEN_11695 ? phv_data_422 : _GEN_6005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6007 = 9'h1a7 == _GEN_11695 ? phv_data_423 : _GEN_6006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6008 = 9'h1a8 == _GEN_11695 ? phv_data_424 : _GEN_6007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6009 = 9'h1a9 == _GEN_11695 ? phv_data_425 : _GEN_6008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6010 = 9'h1aa == _GEN_11695 ? phv_data_426 : _GEN_6009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6011 = 9'h1ab == _GEN_11695 ? phv_data_427 : _GEN_6010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6012 = 9'h1ac == _GEN_11695 ? phv_data_428 : _GEN_6011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6013 = 9'h1ad == _GEN_11695 ? phv_data_429 : _GEN_6012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6014 = 9'h1ae == _GEN_11695 ? phv_data_430 : _GEN_6013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6015 = 9'h1af == _GEN_11695 ? phv_data_431 : _GEN_6014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6016 = 9'h1b0 == _GEN_11695 ? phv_data_432 : _GEN_6015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6017 = 9'h1b1 == _GEN_11695 ? phv_data_433 : _GEN_6016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6018 = 9'h1b2 == _GEN_11695 ? phv_data_434 : _GEN_6017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6019 = 9'h1b3 == _GEN_11695 ? phv_data_435 : _GEN_6018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6020 = 9'h1b4 == _GEN_11695 ? phv_data_436 : _GEN_6019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6021 = 9'h1b5 == _GEN_11695 ? phv_data_437 : _GEN_6020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6022 = 9'h1b6 == _GEN_11695 ? phv_data_438 : _GEN_6021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6023 = 9'h1b7 == _GEN_11695 ? phv_data_439 : _GEN_6022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6024 = 9'h1b8 == _GEN_11695 ? phv_data_440 : _GEN_6023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6025 = 9'h1b9 == _GEN_11695 ? phv_data_441 : _GEN_6024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6026 = 9'h1ba == _GEN_11695 ? phv_data_442 : _GEN_6025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6027 = 9'h1bb == _GEN_11695 ? phv_data_443 : _GEN_6026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6028 = 9'h1bc == _GEN_11695 ? phv_data_444 : _GEN_6027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6029 = 9'h1bd == _GEN_11695 ? phv_data_445 : _GEN_6028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6030 = 9'h1be == _GEN_11695 ? phv_data_446 : _GEN_6029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6031 = 9'h1bf == _GEN_11695 ? phv_data_447 : _GEN_6030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6032 = 9'h1c0 == _GEN_11695 ? phv_data_448 : _GEN_6031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6033 = 9'h1c1 == _GEN_11695 ? phv_data_449 : _GEN_6032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6034 = 9'h1c2 == _GEN_11695 ? phv_data_450 : _GEN_6033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6035 = 9'h1c3 == _GEN_11695 ? phv_data_451 : _GEN_6034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6036 = 9'h1c4 == _GEN_11695 ? phv_data_452 : _GEN_6035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6037 = 9'h1c5 == _GEN_11695 ? phv_data_453 : _GEN_6036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6038 = 9'h1c6 == _GEN_11695 ? phv_data_454 : _GEN_6037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6039 = 9'h1c7 == _GEN_11695 ? phv_data_455 : _GEN_6038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6040 = 9'h1c8 == _GEN_11695 ? phv_data_456 : _GEN_6039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6041 = 9'h1c9 == _GEN_11695 ? phv_data_457 : _GEN_6040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6042 = 9'h1ca == _GEN_11695 ? phv_data_458 : _GEN_6041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6043 = 9'h1cb == _GEN_11695 ? phv_data_459 : _GEN_6042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6044 = 9'h1cc == _GEN_11695 ? phv_data_460 : _GEN_6043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6045 = 9'h1cd == _GEN_11695 ? phv_data_461 : _GEN_6044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6046 = 9'h1ce == _GEN_11695 ? phv_data_462 : _GEN_6045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6047 = 9'h1cf == _GEN_11695 ? phv_data_463 : _GEN_6046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6048 = 9'h1d0 == _GEN_11695 ? phv_data_464 : _GEN_6047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6049 = 9'h1d1 == _GEN_11695 ? phv_data_465 : _GEN_6048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6050 = 9'h1d2 == _GEN_11695 ? phv_data_466 : _GEN_6049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6051 = 9'h1d3 == _GEN_11695 ? phv_data_467 : _GEN_6050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6052 = 9'h1d4 == _GEN_11695 ? phv_data_468 : _GEN_6051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6053 = 9'h1d5 == _GEN_11695 ? phv_data_469 : _GEN_6052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6054 = 9'h1d6 == _GEN_11695 ? phv_data_470 : _GEN_6053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6055 = 9'h1d7 == _GEN_11695 ? phv_data_471 : _GEN_6054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6056 = 9'h1d8 == _GEN_11695 ? phv_data_472 : _GEN_6055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6057 = 9'h1d9 == _GEN_11695 ? phv_data_473 : _GEN_6056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6058 = 9'h1da == _GEN_11695 ? phv_data_474 : _GEN_6057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6059 = 9'h1db == _GEN_11695 ? phv_data_475 : _GEN_6058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6060 = 9'h1dc == _GEN_11695 ? phv_data_476 : _GEN_6059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6061 = 9'h1dd == _GEN_11695 ? phv_data_477 : _GEN_6060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6062 = 9'h1de == _GEN_11695 ? phv_data_478 : _GEN_6061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6063 = 9'h1df == _GEN_11695 ? phv_data_479 : _GEN_6062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6064 = 9'h1e0 == _GEN_11695 ? phv_data_480 : _GEN_6063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6065 = 9'h1e1 == _GEN_11695 ? phv_data_481 : _GEN_6064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6066 = 9'h1e2 == _GEN_11695 ? phv_data_482 : _GEN_6065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6067 = 9'h1e3 == _GEN_11695 ? phv_data_483 : _GEN_6066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6068 = 9'h1e4 == _GEN_11695 ? phv_data_484 : _GEN_6067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6069 = 9'h1e5 == _GEN_11695 ? phv_data_485 : _GEN_6068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6070 = 9'h1e6 == _GEN_11695 ? phv_data_486 : _GEN_6069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6071 = 9'h1e7 == _GEN_11695 ? phv_data_487 : _GEN_6070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6072 = 9'h1e8 == _GEN_11695 ? phv_data_488 : _GEN_6071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6073 = 9'h1e9 == _GEN_11695 ? phv_data_489 : _GEN_6072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6074 = 9'h1ea == _GEN_11695 ? phv_data_490 : _GEN_6073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6075 = 9'h1eb == _GEN_11695 ? phv_data_491 : _GEN_6074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6076 = 9'h1ec == _GEN_11695 ? phv_data_492 : _GEN_6075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6077 = 9'h1ed == _GEN_11695 ? phv_data_493 : _GEN_6076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6078 = 9'h1ee == _GEN_11695 ? phv_data_494 : _GEN_6077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6079 = 9'h1ef == _GEN_11695 ? phv_data_495 : _GEN_6078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6080 = 9'h1f0 == _GEN_11695 ? phv_data_496 : _GEN_6079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6081 = 9'h1f1 == _GEN_11695 ? phv_data_497 : _GEN_6080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6082 = 9'h1f2 == _GEN_11695 ? phv_data_498 : _GEN_6081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6083 = 9'h1f3 == _GEN_11695 ? phv_data_499 : _GEN_6082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6084 = 9'h1f4 == _GEN_11695 ? phv_data_500 : _GEN_6083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6085 = 9'h1f5 == _GEN_11695 ? phv_data_501 : _GEN_6084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6086 = 9'h1f6 == _GEN_11695 ? phv_data_502 : _GEN_6085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6087 = 9'h1f7 == _GEN_11695 ? phv_data_503 : _GEN_6086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6088 = 9'h1f8 == _GEN_11695 ? phv_data_504 : _GEN_6087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6089 = 9'h1f9 == _GEN_11695 ? phv_data_505 : _GEN_6088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6090 = 9'h1fa == _GEN_11695 ? phv_data_506 : _GEN_6089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6091 = 9'h1fb == _GEN_11695 ? phv_data_507 : _GEN_6090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6092 = 9'h1fc == _GEN_11695 ? phv_data_508 : _GEN_6091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6093 = 9'h1fd == _GEN_11695 ? phv_data_509 : _GEN_6092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6094 = 9'h1fe == _GEN_11695 ? phv_data_510 : _GEN_6093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_1 = 9'h1ff == _GEN_11695 ? phv_data_511 : _GEN_6094; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_2_1 = 2'h2 >= offset_2[1:0] & (2'h2 < ending_2 | ending_2 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_11 = {total_offset_hi_2,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_6097 = 8'h1 == total_offset_11 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6098 = 8'h2 == total_offset_11 ? phv_data_2 : _GEN_6097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6099 = 8'h3 == total_offset_11 ? phv_data_3 : _GEN_6098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6100 = 8'h4 == total_offset_11 ? phv_data_4 : _GEN_6099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6101 = 8'h5 == total_offset_11 ? phv_data_5 : _GEN_6100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6102 = 8'h6 == total_offset_11 ? phv_data_6 : _GEN_6101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6103 = 8'h7 == total_offset_11 ? phv_data_7 : _GEN_6102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6104 = 8'h8 == total_offset_11 ? phv_data_8 : _GEN_6103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6105 = 8'h9 == total_offset_11 ? phv_data_9 : _GEN_6104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6106 = 8'ha == total_offset_11 ? phv_data_10 : _GEN_6105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6107 = 8'hb == total_offset_11 ? phv_data_11 : _GEN_6106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6108 = 8'hc == total_offset_11 ? phv_data_12 : _GEN_6107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6109 = 8'hd == total_offset_11 ? phv_data_13 : _GEN_6108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6110 = 8'he == total_offset_11 ? phv_data_14 : _GEN_6109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6111 = 8'hf == total_offset_11 ? phv_data_15 : _GEN_6110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6112 = 8'h10 == total_offset_11 ? phv_data_16 : _GEN_6111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6113 = 8'h11 == total_offset_11 ? phv_data_17 : _GEN_6112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6114 = 8'h12 == total_offset_11 ? phv_data_18 : _GEN_6113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6115 = 8'h13 == total_offset_11 ? phv_data_19 : _GEN_6114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6116 = 8'h14 == total_offset_11 ? phv_data_20 : _GEN_6115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6117 = 8'h15 == total_offset_11 ? phv_data_21 : _GEN_6116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6118 = 8'h16 == total_offset_11 ? phv_data_22 : _GEN_6117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6119 = 8'h17 == total_offset_11 ? phv_data_23 : _GEN_6118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6120 = 8'h18 == total_offset_11 ? phv_data_24 : _GEN_6119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6121 = 8'h19 == total_offset_11 ? phv_data_25 : _GEN_6120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6122 = 8'h1a == total_offset_11 ? phv_data_26 : _GEN_6121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6123 = 8'h1b == total_offset_11 ? phv_data_27 : _GEN_6122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6124 = 8'h1c == total_offset_11 ? phv_data_28 : _GEN_6123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6125 = 8'h1d == total_offset_11 ? phv_data_29 : _GEN_6124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6126 = 8'h1e == total_offset_11 ? phv_data_30 : _GEN_6125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6127 = 8'h1f == total_offset_11 ? phv_data_31 : _GEN_6126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6128 = 8'h20 == total_offset_11 ? phv_data_32 : _GEN_6127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6129 = 8'h21 == total_offset_11 ? phv_data_33 : _GEN_6128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6130 = 8'h22 == total_offset_11 ? phv_data_34 : _GEN_6129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6131 = 8'h23 == total_offset_11 ? phv_data_35 : _GEN_6130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6132 = 8'h24 == total_offset_11 ? phv_data_36 : _GEN_6131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6133 = 8'h25 == total_offset_11 ? phv_data_37 : _GEN_6132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6134 = 8'h26 == total_offset_11 ? phv_data_38 : _GEN_6133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6135 = 8'h27 == total_offset_11 ? phv_data_39 : _GEN_6134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6136 = 8'h28 == total_offset_11 ? phv_data_40 : _GEN_6135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6137 = 8'h29 == total_offset_11 ? phv_data_41 : _GEN_6136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6138 = 8'h2a == total_offset_11 ? phv_data_42 : _GEN_6137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6139 = 8'h2b == total_offset_11 ? phv_data_43 : _GEN_6138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6140 = 8'h2c == total_offset_11 ? phv_data_44 : _GEN_6139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6141 = 8'h2d == total_offset_11 ? phv_data_45 : _GEN_6140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6142 = 8'h2e == total_offset_11 ? phv_data_46 : _GEN_6141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6143 = 8'h2f == total_offset_11 ? phv_data_47 : _GEN_6142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6144 = 8'h30 == total_offset_11 ? phv_data_48 : _GEN_6143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6145 = 8'h31 == total_offset_11 ? phv_data_49 : _GEN_6144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6146 = 8'h32 == total_offset_11 ? phv_data_50 : _GEN_6145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6147 = 8'h33 == total_offset_11 ? phv_data_51 : _GEN_6146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6148 = 8'h34 == total_offset_11 ? phv_data_52 : _GEN_6147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6149 = 8'h35 == total_offset_11 ? phv_data_53 : _GEN_6148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6150 = 8'h36 == total_offset_11 ? phv_data_54 : _GEN_6149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6151 = 8'h37 == total_offset_11 ? phv_data_55 : _GEN_6150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6152 = 8'h38 == total_offset_11 ? phv_data_56 : _GEN_6151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6153 = 8'h39 == total_offset_11 ? phv_data_57 : _GEN_6152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6154 = 8'h3a == total_offset_11 ? phv_data_58 : _GEN_6153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6155 = 8'h3b == total_offset_11 ? phv_data_59 : _GEN_6154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6156 = 8'h3c == total_offset_11 ? phv_data_60 : _GEN_6155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6157 = 8'h3d == total_offset_11 ? phv_data_61 : _GEN_6156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6158 = 8'h3e == total_offset_11 ? phv_data_62 : _GEN_6157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6159 = 8'h3f == total_offset_11 ? phv_data_63 : _GEN_6158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6160 = 8'h40 == total_offset_11 ? phv_data_64 : _GEN_6159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6161 = 8'h41 == total_offset_11 ? phv_data_65 : _GEN_6160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6162 = 8'h42 == total_offset_11 ? phv_data_66 : _GEN_6161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6163 = 8'h43 == total_offset_11 ? phv_data_67 : _GEN_6162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6164 = 8'h44 == total_offset_11 ? phv_data_68 : _GEN_6163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6165 = 8'h45 == total_offset_11 ? phv_data_69 : _GEN_6164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6166 = 8'h46 == total_offset_11 ? phv_data_70 : _GEN_6165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6167 = 8'h47 == total_offset_11 ? phv_data_71 : _GEN_6166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6168 = 8'h48 == total_offset_11 ? phv_data_72 : _GEN_6167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6169 = 8'h49 == total_offset_11 ? phv_data_73 : _GEN_6168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6170 = 8'h4a == total_offset_11 ? phv_data_74 : _GEN_6169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6171 = 8'h4b == total_offset_11 ? phv_data_75 : _GEN_6170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6172 = 8'h4c == total_offset_11 ? phv_data_76 : _GEN_6171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6173 = 8'h4d == total_offset_11 ? phv_data_77 : _GEN_6172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6174 = 8'h4e == total_offset_11 ? phv_data_78 : _GEN_6173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6175 = 8'h4f == total_offset_11 ? phv_data_79 : _GEN_6174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6176 = 8'h50 == total_offset_11 ? phv_data_80 : _GEN_6175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6177 = 8'h51 == total_offset_11 ? phv_data_81 : _GEN_6176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6178 = 8'h52 == total_offset_11 ? phv_data_82 : _GEN_6177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6179 = 8'h53 == total_offset_11 ? phv_data_83 : _GEN_6178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6180 = 8'h54 == total_offset_11 ? phv_data_84 : _GEN_6179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6181 = 8'h55 == total_offset_11 ? phv_data_85 : _GEN_6180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6182 = 8'h56 == total_offset_11 ? phv_data_86 : _GEN_6181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6183 = 8'h57 == total_offset_11 ? phv_data_87 : _GEN_6182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6184 = 8'h58 == total_offset_11 ? phv_data_88 : _GEN_6183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6185 = 8'h59 == total_offset_11 ? phv_data_89 : _GEN_6184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6186 = 8'h5a == total_offset_11 ? phv_data_90 : _GEN_6185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6187 = 8'h5b == total_offset_11 ? phv_data_91 : _GEN_6186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6188 = 8'h5c == total_offset_11 ? phv_data_92 : _GEN_6187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6189 = 8'h5d == total_offset_11 ? phv_data_93 : _GEN_6188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6190 = 8'h5e == total_offset_11 ? phv_data_94 : _GEN_6189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6191 = 8'h5f == total_offset_11 ? phv_data_95 : _GEN_6190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6192 = 8'h60 == total_offset_11 ? phv_data_96 : _GEN_6191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6193 = 8'h61 == total_offset_11 ? phv_data_97 : _GEN_6192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6194 = 8'h62 == total_offset_11 ? phv_data_98 : _GEN_6193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6195 = 8'h63 == total_offset_11 ? phv_data_99 : _GEN_6194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6196 = 8'h64 == total_offset_11 ? phv_data_100 : _GEN_6195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6197 = 8'h65 == total_offset_11 ? phv_data_101 : _GEN_6196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6198 = 8'h66 == total_offset_11 ? phv_data_102 : _GEN_6197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6199 = 8'h67 == total_offset_11 ? phv_data_103 : _GEN_6198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6200 = 8'h68 == total_offset_11 ? phv_data_104 : _GEN_6199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6201 = 8'h69 == total_offset_11 ? phv_data_105 : _GEN_6200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6202 = 8'h6a == total_offset_11 ? phv_data_106 : _GEN_6201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6203 = 8'h6b == total_offset_11 ? phv_data_107 : _GEN_6202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6204 = 8'h6c == total_offset_11 ? phv_data_108 : _GEN_6203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6205 = 8'h6d == total_offset_11 ? phv_data_109 : _GEN_6204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6206 = 8'h6e == total_offset_11 ? phv_data_110 : _GEN_6205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6207 = 8'h6f == total_offset_11 ? phv_data_111 : _GEN_6206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6208 = 8'h70 == total_offset_11 ? phv_data_112 : _GEN_6207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6209 = 8'h71 == total_offset_11 ? phv_data_113 : _GEN_6208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6210 = 8'h72 == total_offset_11 ? phv_data_114 : _GEN_6209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6211 = 8'h73 == total_offset_11 ? phv_data_115 : _GEN_6210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6212 = 8'h74 == total_offset_11 ? phv_data_116 : _GEN_6211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6213 = 8'h75 == total_offset_11 ? phv_data_117 : _GEN_6212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6214 = 8'h76 == total_offset_11 ? phv_data_118 : _GEN_6213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6215 = 8'h77 == total_offset_11 ? phv_data_119 : _GEN_6214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6216 = 8'h78 == total_offset_11 ? phv_data_120 : _GEN_6215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6217 = 8'h79 == total_offset_11 ? phv_data_121 : _GEN_6216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6218 = 8'h7a == total_offset_11 ? phv_data_122 : _GEN_6217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6219 = 8'h7b == total_offset_11 ? phv_data_123 : _GEN_6218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6220 = 8'h7c == total_offset_11 ? phv_data_124 : _GEN_6219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6221 = 8'h7d == total_offset_11 ? phv_data_125 : _GEN_6220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6222 = 8'h7e == total_offset_11 ? phv_data_126 : _GEN_6221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6223 = 8'h7f == total_offset_11 ? phv_data_127 : _GEN_6222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6224 = 8'h80 == total_offset_11 ? phv_data_128 : _GEN_6223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6225 = 8'h81 == total_offset_11 ? phv_data_129 : _GEN_6224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6226 = 8'h82 == total_offset_11 ? phv_data_130 : _GEN_6225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6227 = 8'h83 == total_offset_11 ? phv_data_131 : _GEN_6226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6228 = 8'h84 == total_offset_11 ? phv_data_132 : _GEN_6227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6229 = 8'h85 == total_offset_11 ? phv_data_133 : _GEN_6228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6230 = 8'h86 == total_offset_11 ? phv_data_134 : _GEN_6229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6231 = 8'h87 == total_offset_11 ? phv_data_135 : _GEN_6230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6232 = 8'h88 == total_offset_11 ? phv_data_136 : _GEN_6231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6233 = 8'h89 == total_offset_11 ? phv_data_137 : _GEN_6232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6234 = 8'h8a == total_offset_11 ? phv_data_138 : _GEN_6233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6235 = 8'h8b == total_offset_11 ? phv_data_139 : _GEN_6234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6236 = 8'h8c == total_offset_11 ? phv_data_140 : _GEN_6235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6237 = 8'h8d == total_offset_11 ? phv_data_141 : _GEN_6236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6238 = 8'h8e == total_offset_11 ? phv_data_142 : _GEN_6237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6239 = 8'h8f == total_offset_11 ? phv_data_143 : _GEN_6238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6240 = 8'h90 == total_offset_11 ? phv_data_144 : _GEN_6239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6241 = 8'h91 == total_offset_11 ? phv_data_145 : _GEN_6240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6242 = 8'h92 == total_offset_11 ? phv_data_146 : _GEN_6241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6243 = 8'h93 == total_offset_11 ? phv_data_147 : _GEN_6242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6244 = 8'h94 == total_offset_11 ? phv_data_148 : _GEN_6243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6245 = 8'h95 == total_offset_11 ? phv_data_149 : _GEN_6244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6246 = 8'h96 == total_offset_11 ? phv_data_150 : _GEN_6245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6247 = 8'h97 == total_offset_11 ? phv_data_151 : _GEN_6246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6248 = 8'h98 == total_offset_11 ? phv_data_152 : _GEN_6247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6249 = 8'h99 == total_offset_11 ? phv_data_153 : _GEN_6248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6250 = 8'h9a == total_offset_11 ? phv_data_154 : _GEN_6249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6251 = 8'h9b == total_offset_11 ? phv_data_155 : _GEN_6250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6252 = 8'h9c == total_offset_11 ? phv_data_156 : _GEN_6251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6253 = 8'h9d == total_offset_11 ? phv_data_157 : _GEN_6252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6254 = 8'h9e == total_offset_11 ? phv_data_158 : _GEN_6253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6255 = 8'h9f == total_offset_11 ? phv_data_159 : _GEN_6254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6256 = 8'ha0 == total_offset_11 ? phv_data_160 : _GEN_6255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6257 = 8'ha1 == total_offset_11 ? phv_data_161 : _GEN_6256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6258 = 8'ha2 == total_offset_11 ? phv_data_162 : _GEN_6257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6259 = 8'ha3 == total_offset_11 ? phv_data_163 : _GEN_6258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6260 = 8'ha4 == total_offset_11 ? phv_data_164 : _GEN_6259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6261 = 8'ha5 == total_offset_11 ? phv_data_165 : _GEN_6260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6262 = 8'ha6 == total_offset_11 ? phv_data_166 : _GEN_6261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6263 = 8'ha7 == total_offset_11 ? phv_data_167 : _GEN_6262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6264 = 8'ha8 == total_offset_11 ? phv_data_168 : _GEN_6263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6265 = 8'ha9 == total_offset_11 ? phv_data_169 : _GEN_6264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6266 = 8'haa == total_offset_11 ? phv_data_170 : _GEN_6265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6267 = 8'hab == total_offset_11 ? phv_data_171 : _GEN_6266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6268 = 8'hac == total_offset_11 ? phv_data_172 : _GEN_6267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6269 = 8'had == total_offset_11 ? phv_data_173 : _GEN_6268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6270 = 8'hae == total_offset_11 ? phv_data_174 : _GEN_6269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6271 = 8'haf == total_offset_11 ? phv_data_175 : _GEN_6270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6272 = 8'hb0 == total_offset_11 ? phv_data_176 : _GEN_6271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6273 = 8'hb1 == total_offset_11 ? phv_data_177 : _GEN_6272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6274 = 8'hb2 == total_offset_11 ? phv_data_178 : _GEN_6273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6275 = 8'hb3 == total_offset_11 ? phv_data_179 : _GEN_6274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6276 = 8'hb4 == total_offset_11 ? phv_data_180 : _GEN_6275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6277 = 8'hb5 == total_offset_11 ? phv_data_181 : _GEN_6276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6278 = 8'hb6 == total_offset_11 ? phv_data_182 : _GEN_6277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6279 = 8'hb7 == total_offset_11 ? phv_data_183 : _GEN_6278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6280 = 8'hb8 == total_offset_11 ? phv_data_184 : _GEN_6279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6281 = 8'hb9 == total_offset_11 ? phv_data_185 : _GEN_6280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6282 = 8'hba == total_offset_11 ? phv_data_186 : _GEN_6281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6283 = 8'hbb == total_offset_11 ? phv_data_187 : _GEN_6282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6284 = 8'hbc == total_offset_11 ? phv_data_188 : _GEN_6283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6285 = 8'hbd == total_offset_11 ? phv_data_189 : _GEN_6284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6286 = 8'hbe == total_offset_11 ? phv_data_190 : _GEN_6285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6287 = 8'hbf == total_offset_11 ? phv_data_191 : _GEN_6286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6288 = 8'hc0 == total_offset_11 ? phv_data_192 : _GEN_6287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6289 = 8'hc1 == total_offset_11 ? phv_data_193 : _GEN_6288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6290 = 8'hc2 == total_offset_11 ? phv_data_194 : _GEN_6289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6291 = 8'hc3 == total_offset_11 ? phv_data_195 : _GEN_6290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6292 = 8'hc4 == total_offset_11 ? phv_data_196 : _GEN_6291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6293 = 8'hc5 == total_offset_11 ? phv_data_197 : _GEN_6292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6294 = 8'hc6 == total_offset_11 ? phv_data_198 : _GEN_6293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6295 = 8'hc7 == total_offset_11 ? phv_data_199 : _GEN_6294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6296 = 8'hc8 == total_offset_11 ? phv_data_200 : _GEN_6295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6297 = 8'hc9 == total_offset_11 ? phv_data_201 : _GEN_6296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6298 = 8'hca == total_offset_11 ? phv_data_202 : _GEN_6297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6299 = 8'hcb == total_offset_11 ? phv_data_203 : _GEN_6298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6300 = 8'hcc == total_offset_11 ? phv_data_204 : _GEN_6299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6301 = 8'hcd == total_offset_11 ? phv_data_205 : _GEN_6300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6302 = 8'hce == total_offset_11 ? phv_data_206 : _GEN_6301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6303 = 8'hcf == total_offset_11 ? phv_data_207 : _GEN_6302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6304 = 8'hd0 == total_offset_11 ? phv_data_208 : _GEN_6303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6305 = 8'hd1 == total_offset_11 ? phv_data_209 : _GEN_6304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6306 = 8'hd2 == total_offset_11 ? phv_data_210 : _GEN_6305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6307 = 8'hd3 == total_offset_11 ? phv_data_211 : _GEN_6306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6308 = 8'hd4 == total_offset_11 ? phv_data_212 : _GEN_6307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6309 = 8'hd5 == total_offset_11 ? phv_data_213 : _GEN_6308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6310 = 8'hd6 == total_offset_11 ? phv_data_214 : _GEN_6309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6311 = 8'hd7 == total_offset_11 ? phv_data_215 : _GEN_6310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6312 = 8'hd8 == total_offset_11 ? phv_data_216 : _GEN_6311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6313 = 8'hd9 == total_offset_11 ? phv_data_217 : _GEN_6312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6314 = 8'hda == total_offset_11 ? phv_data_218 : _GEN_6313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6315 = 8'hdb == total_offset_11 ? phv_data_219 : _GEN_6314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6316 = 8'hdc == total_offset_11 ? phv_data_220 : _GEN_6315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6317 = 8'hdd == total_offset_11 ? phv_data_221 : _GEN_6316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6318 = 8'hde == total_offset_11 ? phv_data_222 : _GEN_6317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6319 = 8'hdf == total_offset_11 ? phv_data_223 : _GEN_6318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6320 = 8'he0 == total_offset_11 ? phv_data_224 : _GEN_6319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6321 = 8'he1 == total_offset_11 ? phv_data_225 : _GEN_6320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6322 = 8'he2 == total_offset_11 ? phv_data_226 : _GEN_6321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6323 = 8'he3 == total_offset_11 ? phv_data_227 : _GEN_6322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6324 = 8'he4 == total_offset_11 ? phv_data_228 : _GEN_6323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6325 = 8'he5 == total_offset_11 ? phv_data_229 : _GEN_6324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6326 = 8'he6 == total_offset_11 ? phv_data_230 : _GEN_6325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6327 = 8'he7 == total_offset_11 ? phv_data_231 : _GEN_6326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6328 = 8'he8 == total_offset_11 ? phv_data_232 : _GEN_6327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6329 = 8'he9 == total_offset_11 ? phv_data_233 : _GEN_6328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6330 = 8'hea == total_offset_11 ? phv_data_234 : _GEN_6329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6331 = 8'heb == total_offset_11 ? phv_data_235 : _GEN_6330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6332 = 8'hec == total_offset_11 ? phv_data_236 : _GEN_6331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6333 = 8'hed == total_offset_11 ? phv_data_237 : _GEN_6332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6334 = 8'hee == total_offset_11 ? phv_data_238 : _GEN_6333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6335 = 8'hef == total_offset_11 ? phv_data_239 : _GEN_6334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6336 = 8'hf0 == total_offset_11 ? phv_data_240 : _GEN_6335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6337 = 8'hf1 == total_offset_11 ? phv_data_241 : _GEN_6336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6338 = 8'hf2 == total_offset_11 ? phv_data_242 : _GEN_6337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6339 = 8'hf3 == total_offset_11 ? phv_data_243 : _GEN_6338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6340 = 8'hf4 == total_offset_11 ? phv_data_244 : _GEN_6339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6341 = 8'hf5 == total_offset_11 ? phv_data_245 : _GEN_6340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6342 = 8'hf6 == total_offset_11 ? phv_data_246 : _GEN_6341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6343 = 8'hf7 == total_offset_11 ? phv_data_247 : _GEN_6342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6344 = 8'hf8 == total_offset_11 ? phv_data_248 : _GEN_6343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6345 = 8'hf9 == total_offset_11 ? phv_data_249 : _GEN_6344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6346 = 8'hfa == total_offset_11 ? phv_data_250 : _GEN_6345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6347 = 8'hfb == total_offset_11 ? phv_data_251 : _GEN_6346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6348 = 8'hfc == total_offset_11 ? phv_data_252 : _GEN_6347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6349 = 8'hfd == total_offset_11 ? phv_data_253 : _GEN_6348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6350 = 8'hfe == total_offset_11 ? phv_data_254 : _GEN_6349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6351 = 8'hff == total_offset_11 ? phv_data_255 : _GEN_6350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_11951 = {{1'd0}, total_offset_11}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6352 = 9'h100 == _GEN_11951 ? phv_data_256 : _GEN_6351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6353 = 9'h101 == _GEN_11951 ? phv_data_257 : _GEN_6352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6354 = 9'h102 == _GEN_11951 ? phv_data_258 : _GEN_6353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6355 = 9'h103 == _GEN_11951 ? phv_data_259 : _GEN_6354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6356 = 9'h104 == _GEN_11951 ? phv_data_260 : _GEN_6355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6357 = 9'h105 == _GEN_11951 ? phv_data_261 : _GEN_6356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6358 = 9'h106 == _GEN_11951 ? phv_data_262 : _GEN_6357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6359 = 9'h107 == _GEN_11951 ? phv_data_263 : _GEN_6358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6360 = 9'h108 == _GEN_11951 ? phv_data_264 : _GEN_6359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6361 = 9'h109 == _GEN_11951 ? phv_data_265 : _GEN_6360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6362 = 9'h10a == _GEN_11951 ? phv_data_266 : _GEN_6361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6363 = 9'h10b == _GEN_11951 ? phv_data_267 : _GEN_6362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6364 = 9'h10c == _GEN_11951 ? phv_data_268 : _GEN_6363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6365 = 9'h10d == _GEN_11951 ? phv_data_269 : _GEN_6364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6366 = 9'h10e == _GEN_11951 ? phv_data_270 : _GEN_6365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6367 = 9'h10f == _GEN_11951 ? phv_data_271 : _GEN_6366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6368 = 9'h110 == _GEN_11951 ? phv_data_272 : _GEN_6367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6369 = 9'h111 == _GEN_11951 ? phv_data_273 : _GEN_6368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6370 = 9'h112 == _GEN_11951 ? phv_data_274 : _GEN_6369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6371 = 9'h113 == _GEN_11951 ? phv_data_275 : _GEN_6370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6372 = 9'h114 == _GEN_11951 ? phv_data_276 : _GEN_6371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6373 = 9'h115 == _GEN_11951 ? phv_data_277 : _GEN_6372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6374 = 9'h116 == _GEN_11951 ? phv_data_278 : _GEN_6373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6375 = 9'h117 == _GEN_11951 ? phv_data_279 : _GEN_6374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6376 = 9'h118 == _GEN_11951 ? phv_data_280 : _GEN_6375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6377 = 9'h119 == _GEN_11951 ? phv_data_281 : _GEN_6376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6378 = 9'h11a == _GEN_11951 ? phv_data_282 : _GEN_6377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6379 = 9'h11b == _GEN_11951 ? phv_data_283 : _GEN_6378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6380 = 9'h11c == _GEN_11951 ? phv_data_284 : _GEN_6379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6381 = 9'h11d == _GEN_11951 ? phv_data_285 : _GEN_6380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6382 = 9'h11e == _GEN_11951 ? phv_data_286 : _GEN_6381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6383 = 9'h11f == _GEN_11951 ? phv_data_287 : _GEN_6382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6384 = 9'h120 == _GEN_11951 ? phv_data_288 : _GEN_6383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6385 = 9'h121 == _GEN_11951 ? phv_data_289 : _GEN_6384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6386 = 9'h122 == _GEN_11951 ? phv_data_290 : _GEN_6385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6387 = 9'h123 == _GEN_11951 ? phv_data_291 : _GEN_6386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6388 = 9'h124 == _GEN_11951 ? phv_data_292 : _GEN_6387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6389 = 9'h125 == _GEN_11951 ? phv_data_293 : _GEN_6388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6390 = 9'h126 == _GEN_11951 ? phv_data_294 : _GEN_6389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6391 = 9'h127 == _GEN_11951 ? phv_data_295 : _GEN_6390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6392 = 9'h128 == _GEN_11951 ? phv_data_296 : _GEN_6391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6393 = 9'h129 == _GEN_11951 ? phv_data_297 : _GEN_6392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6394 = 9'h12a == _GEN_11951 ? phv_data_298 : _GEN_6393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6395 = 9'h12b == _GEN_11951 ? phv_data_299 : _GEN_6394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6396 = 9'h12c == _GEN_11951 ? phv_data_300 : _GEN_6395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6397 = 9'h12d == _GEN_11951 ? phv_data_301 : _GEN_6396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6398 = 9'h12e == _GEN_11951 ? phv_data_302 : _GEN_6397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6399 = 9'h12f == _GEN_11951 ? phv_data_303 : _GEN_6398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6400 = 9'h130 == _GEN_11951 ? phv_data_304 : _GEN_6399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6401 = 9'h131 == _GEN_11951 ? phv_data_305 : _GEN_6400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6402 = 9'h132 == _GEN_11951 ? phv_data_306 : _GEN_6401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6403 = 9'h133 == _GEN_11951 ? phv_data_307 : _GEN_6402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6404 = 9'h134 == _GEN_11951 ? phv_data_308 : _GEN_6403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6405 = 9'h135 == _GEN_11951 ? phv_data_309 : _GEN_6404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6406 = 9'h136 == _GEN_11951 ? phv_data_310 : _GEN_6405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6407 = 9'h137 == _GEN_11951 ? phv_data_311 : _GEN_6406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6408 = 9'h138 == _GEN_11951 ? phv_data_312 : _GEN_6407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6409 = 9'h139 == _GEN_11951 ? phv_data_313 : _GEN_6408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6410 = 9'h13a == _GEN_11951 ? phv_data_314 : _GEN_6409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6411 = 9'h13b == _GEN_11951 ? phv_data_315 : _GEN_6410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6412 = 9'h13c == _GEN_11951 ? phv_data_316 : _GEN_6411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6413 = 9'h13d == _GEN_11951 ? phv_data_317 : _GEN_6412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6414 = 9'h13e == _GEN_11951 ? phv_data_318 : _GEN_6413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6415 = 9'h13f == _GEN_11951 ? phv_data_319 : _GEN_6414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6416 = 9'h140 == _GEN_11951 ? phv_data_320 : _GEN_6415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6417 = 9'h141 == _GEN_11951 ? phv_data_321 : _GEN_6416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6418 = 9'h142 == _GEN_11951 ? phv_data_322 : _GEN_6417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6419 = 9'h143 == _GEN_11951 ? phv_data_323 : _GEN_6418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6420 = 9'h144 == _GEN_11951 ? phv_data_324 : _GEN_6419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6421 = 9'h145 == _GEN_11951 ? phv_data_325 : _GEN_6420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6422 = 9'h146 == _GEN_11951 ? phv_data_326 : _GEN_6421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6423 = 9'h147 == _GEN_11951 ? phv_data_327 : _GEN_6422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6424 = 9'h148 == _GEN_11951 ? phv_data_328 : _GEN_6423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6425 = 9'h149 == _GEN_11951 ? phv_data_329 : _GEN_6424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6426 = 9'h14a == _GEN_11951 ? phv_data_330 : _GEN_6425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6427 = 9'h14b == _GEN_11951 ? phv_data_331 : _GEN_6426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6428 = 9'h14c == _GEN_11951 ? phv_data_332 : _GEN_6427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6429 = 9'h14d == _GEN_11951 ? phv_data_333 : _GEN_6428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6430 = 9'h14e == _GEN_11951 ? phv_data_334 : _GEN_6429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6431 = 9'h14f == _GEN_11951 ? phv_data_335 : _GEN_6430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6432 = 9'h150 == _GEN_11951 ? phv_data_336 : _GEN_6431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6433 = 9'h151 == _GEN_11951 ? phv_data_337 : _GEN_6432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6434 = 9'h152 == _GEN_11951 ? phv_data_338 : _GEN_6433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6435 = 9'h153 == _GEN_11951 ? phv_data_339 : _GEN_6434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6436 = 9'h154 == _GEN_11951 ? phv_data_340 : _GEN_6435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6437 = 9'h155 == _GEN_11951 ? phv_data_341 : _GEN_6436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6438 = 9'h156 == _GEN_11951 ? phv_data_342 : _GEN_6437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6439 = 9'h157 == _GEN_11951 ? phv_data_343 : _GEN_6438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6440 = 9'h158 == _GEN_11951 ? phv_data_344 : _GEN_6439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6441 = 9'h159 == _GEN_11951 ? phv_data_345 : _GEN_6440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6442 = 9'h15a == _GEN_11951 ? phv_data_346 : _GEN_6441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6443 = 9'h15b == _GEN_11951 ? phv_data_347 : _GEN_6442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6444 = 9'h15c == _GEN_11951 ? phv_data_348 : _GEN_6443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6445 = 9'h15d == _GEN_11951 ? phv_data_349 : _GEN_6444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6446 = 9'h15e == _GEN_11951 ? phv_data_350 : _GEN_6445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6447 = 9'h15f == _GEN_11951 ? phv_data_351 : _GEN_6446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6448 = 9'h160 == _GEN_11951 ? phv_data_352 : _GEN_6447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6449 = 9'h161 == _GEN_11951 ? phv_data_353 : _GEN_6448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6450 = 9'h162 == _GEN_11951 ? phv_data_354 : _GEN_6449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6451 = 9'h163 == _GEN_11951 ? phv_data_355 : _GEN_6450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6452 = 9'h164 == _GEN_11951 ? phv_data_356 : _GEN_6451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6453 = 9'h165 == _GEN_11951 ? phv_data_357 : _GEN_6452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6454 = 9'h166 == _GEN_11951 ? phv_data_358 : _GEN_6453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6455 = 9'h167 == _GEN_11951 ? phv_data_359 : _GEN_6454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6456 = 9'h168 == _GEN_11951 ? phv_data_360 : _GEN_6455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6457 = 9'h169 == _GEN_11951 ? phv_data_361 : _GEN_6456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6458 = 9'h16a == _GEN_11951 ? phv_data_362 : _GEN_6457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6459 = 9'h16b == _GEN_11951 ? phv_data_363 : _GEN_6458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6460 = 9'h16c == _GEN_11951 ? phv_data_364 : _GEN_6459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6461 = 9'h16d == _GEN_11951 ? phv_data_365 : _GEN_6460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6462 = 9'h16e == _GEN_11951 ? phv_data_366 : _GEN_6461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6463 = 9'h16f == _GEN_11951 ? phv_data_367 : _GEN_6462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6464 = 9'h170 == _GEN_11951 ? phv_data_368 : _GEN_6463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6465 = 9'h171 == _GEN_11951 ? phv_data_369 : _GEN_6464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6466 = 9'h172 == _GEN_11951 ? phv_data_370 : _GEN_6465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6467 = 9'h173 == _GEN_11951 ? phv_data_371 : _GEN_6466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6468 = 9'h174 == _GEN_11951 ? phv_data_372 : _GEN_6467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6469 = 9'h175 == _GEN_11951 ? phv_data_373 : _GEN_6468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6470 = 9'h176 == _GEN_11951 ? phv_data_374 : _GEN_6469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6471 = 9'h177 == _GEN_11951 ? phv_data_375 : _GEN_6470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6472 = 9'h178 == _GEN_11951 ? phv_data_376 : _GEN_6471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6473 = 9'h179 == _GEN_11951 ? phv_data_377 : _GEN_6472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6474 = 9'h17a == _GEN_11951 ? phv_data_378 : _GEN_6473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6475 = 9'h17b == _GEN_11951 ? phv_data_379 : _GEN_6474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6476 = 9'h17c == _GEN_11951 ? phv_data_380 : _GEN_6475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6477 = 9'h17d == _GEN_11951 ? phv_data_381 : _GEN_6476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6478 = 9'h17e == _GEN_11951 ? phv_data_382 : _GEN_6477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6479 = 9'h17f == _GEN_11951 ? phv_data_383 : _GEN_6478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6480 = 9'h180 == _GEN_11951 ? phv_data_384 : _GEN_6479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6481 = 9'h181 == _GEN_11951 ? phv_data_385 : _GEN_6480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6482 = 9'h182 == _GEN_11951 ? phv_data_386 : _GEN_6481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6483 = 9'h183 == _GEN_11951 ? phv_data_387 : _GEN_6482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6484 = 9'h184 == _GEN_11951 ? phv_data_388 : _GEN_6483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6485 = 9'h185 == _GEN_11951 ? phv_data_389 : _GEN_6484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6486 = 9'h186 == _GEN_11951 ? phv_data_390 : _GEN_6485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6487 = 9'h187 == _GEN_11951 ? phv_data_391 : _GEN_6486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6488 = 9'h188 == _GEN_11951 ? phv_data_392 : _GEN_6487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6489 = 9'h189 == _GEN_11951 ? phv_data_393 : _GEN_6488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6490 = 9'h18a == _GEN_11951 ? phv_data_394 : _GEN_6489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6491 = 9'h18b == _GEN_11951 ? phv_data_395 : _GEN_6490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6492 = 9'h18c == _GEN_11951 ? phv_data_396 : _GEN_6491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6493 = 9'h18d == _GEN_11951 ? phv_data_397 : _GEN_6492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6494 = 9'h18e == _GEN_11951 ? phv_data_398 : _GEN_6493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6495 = 9'h18f == _GEN_11951 ? phv_data_399 : _GEN_6494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6496 = 9'h190 == _GEN_11951 ? phv_data_400 : _GEN_6495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6497 = 9'h191 == _GEN_11951 ? phv_data_401 : _GEN_6496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6498 = 9'h192 == _GEN_11951 ? phv_data_402 : _GEN_6497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6499 = 9'h193 == _GEN_11951 ? phv_data_403 : _GEN_6498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6500 = 9'h194 == _GEN_11951 ? phv_data_404 : _GEN_6499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6501 = 9'h195 == _GEN_11951 ? phv_data_405 : _GEN_6500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6502 = 9'h196 == _GEN_11951 ? phv_data_406 : _GEN_6501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6503 = 9'h197 == _GEN_11951 ? phv_data_407 : _GEN_6502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6504 = 9'h198 == _GEN_11951 ? phv_data_408 : _GEN_6503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6505 = 9'h199 == _GEN_11951 ? phv_data_409 : _GEN_6504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6506 = 9'h19a == _GEN_11951 ? phv_data_410 : _GEN_6505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6507 = 9'h19b == _GEN_11951 ? phv_data_411 : _GEN_6506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6508 = 9'h19c == _GEN_11951 ? phv_data_412 : _GEN_6507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6509 = 9'h19d == _GEN_11951 ? phv_data_413 : _GEN_6508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6510 = 9'h19e == _GEN_11951 ? phv_data_414 : _GEN_6509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6511 = 9'h19f == _GEN_11951 ? phv_data_415 : _GEN_6510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6512 = 9'h1a0 == _GEN_11951 ? phv_data_416 : _GEN_6511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6513 = 9'h1a1 == _GEN_11951 ? phv_data_417 : _GEN_6512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6514 = 9'h1a2 == _GEN_11951 ? phv_data_418 : _GEN_6513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6515 = 9'h1a3 == _GEN_11951 ? phv_data_419 : _GEN_6514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6516 = 9'h1a4 == _GEN_11951 ? phv_data_420 : _GEN_6515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6517 = 9'h1a5 == _GEN_11951 ? phv_data_421 : _GEN_6516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6518 = 9'h1a6 == _GEN_11951 ? phv_data_422 : _GEN_6517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6519 = 9'h1a7 == _GEN_11951 ? phv_data_423 : _GEN_6518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6520 = 9'h1a8 == _GEN_11951 ? phv_data_424 : _GEN_6519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6521 = 9'h1a9 == _GEN_11951 ? phv_data_425 : _GEN_6520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6522 = 9'h1aa == _GEN_11951 ? phv_data_426 : _GEN_6521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6523 = 9'h1ab == _GEN_11951 ? phv_data_427 : _GEN_6522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6524 = 9'h1ac == _GEN_11951 ? phv_data_428 : _GEN_6523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6525 = 9'h1ad == _GEN_11951 ? phv_data_429 : _GEN_6524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6526 = 9'h1ae == _GEN_11951 ? phv_data_430 : _GEN_6525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6527 = 9'h1af == _GEN_11951 ? phv_data_431 : _GEN_6526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6528 = 9'h1b0 == _GEN_11951 ? phv_data_432 : _GEN_6527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6529 = 9'h1b1 == _GEN_11951 ? phv_data_433 : _GEN_6528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6530 = 9'h1b2 == _GEN_11951 ? phv_data_434 : _GEN_6529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6531 = 9'h1b3 == _GEN_11951 ? phv_data_435 : _GEN_6530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6532 = 9'h1b4 == _GEN_11951 ? phv_data_436 : _GEN_6531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6533 = 9'h1b5 == _GEN_11951 ? phv_data_437 : _GEN_6532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6534 = 9'h1b6 == _GEN_11951 ? phv_data_438 : _GEN_6533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6535 = 9'h1b7 == _GEN_11951 ? phv_data_439 : _GEN_6534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6536 = 9'h1b8 == _GEN_11951 ? phv_data_440 : _GEN_6535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6537 = 9'h1b9 == _GEN_11951 ? phv_data_441 : _GEN_6536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6538 = 9'h1ba == _GEN_11951 ? phv_data_442 : _GEN_6537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6539 = 9'h1bb == _GEN_11951 ? phv_data_443 : _GEN_6538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6540 = 9'h1bc == _GEN_11951 ? phv_data_444 : _GEN_6539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6541 = 9'h1bd == _GEN_11951 ? phv_data_445 : _GEN_6540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6542 = 9'h1be == _GEN_11951 ? phv_data_446 : _GEN_6541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6543 = 9'h1bf == _GEN_11951 ? phv_data_447 : _GEN_6542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6544 = 9'h1c0 == _GEN_11951 ? phv_data_448 : _GEN_6543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6545 = 9'h1c1 == _GEN_11951 ? phv_data_449 : _GEN_6544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6546 = 9'h1c2 == _GEN_11951 ? phv_data_450 : _GEN_6545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6547 = 9'h1c3 == _GEN_11951 ? phv_data_451 : _GEN_6546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6548 = 9'h1c4 == _GEN_11951 ? phv_data_452 : _GEN_6547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6549 = 9'h1c5 == _GEN_11951 ? phv_data_453 : _GEN_6548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6550 = 9'h1c6 == _GEN_11951 ? phv_data_454 : _GEN_6549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6551 = 9'h1c7 == _GEN_11951 ? phv_data_455 : _GEN_6550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6552 = 9'h1c8 == _GEN_11951 ? phv_data_456 : _GEN_6551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6553 = 9'h1c9 == _GEN_11951 ? phv_data_457 : _GEN_6552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6554 = 9'h1ca == _GEN_11951 ? phv_data_458 : _GEN_6553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6555 = 9'h1cb == _GEN_11951 ? phv_data_459 : _GEN_6554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6556 = 9'h1cc == _GEN_11951 ? phv_data_460 : _GEN_6555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6557 = 9'h1cd == _GEN_11951 ? phv_data_461 : _GEN_6556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6558 = 9'h1ce == _GEN_11951 ? phv_data_462 : _GEN_6557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6559 = 9'h1cf == _GEN_11951 ? phv_data_463 : _GEN_6558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6560 = 9'h1d0 == _GEN_11951 ? phv_data_464 : _GEN_6559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6561 = 9'h1d1 == _GEN_11951 ? phv_data_465 : _GEN_6560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6562 = 9'h1d2 == _GEN_11951 ? phv_data_466 : _GEN_6561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6563 = 9'h1d3 == _GEN_11951 ? phv_data_467 : _GEN_6562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6564 = 9'h1d4 == _GEN_11951 ? phv_data_468 : _GEN_6563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6565 = 9'h1d5 == _GEN_11951 ? phv_data_469 : _GEN_6564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6566 = 9'h1d6 == _GEN_11951 ? phv_data_470 : _GEN_6565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6567 = 9'h1d7 == _GEN_11951 ? phv_data_471 : _GEN_6566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6568 = 9'h1d8 == _GEN_11951 ? phv_data_472 : _GEN_6567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6569 = 9'h1d9 == _GEN_11951 ? phv_data_473 : _GEN_6568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6570 = 9'h1da == _GEN_11951 ? phv_data_474 : _GEN_6569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6571 = 9'h1db == _GEN_11951 ? phv_data_475 : _GEN_6570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6572 = 9'h1dc == _GEN_11951 ? phv_data_476 : _GEN_6571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6573 = 9'h1dd == _GEN_11951 ? phv_data_477 : _GEN_6572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6574 = 9'h1de == _GEN_11951 ? phv_data_478 : _GEN_6573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6575 = 9'h1df == _GEN_11951 ? phv_data_479 : _GEN_6574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6576 = 9'h1e0 == _GEN_11951 ? phv_data_480 : _GEN_6575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6577 = 9'h1e1 == _GEN_11951 ? phv_data_481 : _GEN_6576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6578 = 9'h1e2 == _GEN_11951 ? phv_data_482 : _GEN_6577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6579 = 9'h1e3 == _GEN_11951 ? phv_data_483 : _GEN_6578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6580 = 9'h1e4 == _GEN_11951 ? phv_data_484 : _GEN_6579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6581 = 9'h1e5 == _GEN_11951 ? phv_data_485 : _GEN_6580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6582 = 9'h1e6 == _GEN_11951 ? phv_data_486 : _GEN_6581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6583 = 9'h1e7 == _GEN_11951 ? phv_data_487 : _GEN_6582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6584 = 9'h1e8 == _GEN_11951 ? phv_data_488 : _GEN_6583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6585 = 9'h1e9 == _GEN_11951 ? phv_data_489 : _GEN_6584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6586 = 9'h1ea == _GEN_11951 ? phv_data_490 : _GEN_6585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6587 = 9'h1eb == _GEN_11951 ? phv_data_491 : _GEN_6586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6588 = 9'h1ec == _GEN_11951 ? phv_data_492 : _GEN_6587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6589 = 9'h1ed == _GEN_11951 ? phv_data_493 : _GEN_6588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6590 = 9'h1ee == _GEN_11951 ? phv_data_494 : _GEN_6589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6591 = 9'h1ef == _GEN_11951 ? phv_data_495 : _GEN_6590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6592 = 9'h1f0 == _GEN_11951 ? phv_data_496 : _GEN_6591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6593 = 9'h1f1 == _GEN_11951 ? phv_data_497 : _GEN_6592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6594 = 9'h1f2 == _GEN_11951 ? phv_data_498 : _GEN_6593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6595 = 9'h1f3 == _GEN_11951 ? phv_data_499 : _GEN_6594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6596 = 9'h1f4 == _GEN_11951 ? phv_data_500 : _GEN_6595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6597 = 9'h1f5 == _GEN_11951 ? phv_data_501 : _GEN_6596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6598 = 9'h1f6 == _GEN_11951 ? phv_data_502 : _GEN_6597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6599 = 9'h1f7 == _GEN_11951 ? phv_data_503 : _GEN_6598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6600 = 9'h1f8 == _GEN_11951 ? phv_data_504 : _GEN_6599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6601 = 9'h1f9 == _GEN_11951 ? phv_data_505 : _GEN_6600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6602 = 9'h1fa == _GEN_11951 ? phv_data_506 : _GEN_6601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6603 = 9'h1fb == _GEN_11951 ? phv_data_507 : _GEN_6602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6604 = 9'h1fc == _GEN_11951 ? phv_data_508 : _GEN_6603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6605 = 9'h1fd == _GEN_11951 ? phv_data_509 : _GEN_6604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6606 = 9'h1fe == _GEN_11951 ? phv_data_510 : _GEN_6605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_2_0 = 9'h1ff == _GEN_11951 ? phv_data_511 : _GEN_6606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_2_T = {bytes_2_0,bytes_2_1,bytes_2_2,bytes_2_3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_2_T = {_mask_3_T_17,mask_2_1,mask_2_2,mask_2_3}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_2 = io_field_out_2_lo[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_2 = io_field_out_2_lo[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _local_offset_T_113 = {{1'd0}, args_offset_2}; // @[executor.scala 222:61]
  wire [2:0] local_offset_56 = _local_offset_T_113[2:0]; // @[executor.scala 222:61]
  wire [7:0] _GEN_6609 = 3'h1 == local_offset_56 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6610 = 3'h2 == local_offset_56 ? args_2 : _GEN_6609; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6611 = 3'h3 == local_offset_56 ? args_3 : _GEN_6610; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6612 = 3'h4 == local_offset_56 ? args_4 : _GEN_6611; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6613 = 3'h5 == local_offset_56 ? args_5 : _GEN_6612; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6614 = 3'h6 == local_offset_56 ? args_6 : _GEN_6613; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6615 = 3'h1 == args_length_2 ? _GEN_6614 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [2:0] local_offset_57 = 3'h1 + args_offset_2; // @[executor.scala 222:61]
  wire [7:0] _GEN_6617 = 3'h1 == local_offset_57 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6618 = 3'h2 == local_offset_57 ? args_2 : _GEN_6617; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6619 = 3'h3 == local_offset_57 ? args_3 : _GEN_6618; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6620 = 3'h4 == local_offset_57 ? args_4 : _GEN_6619; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6621 = 3'h5 == local_offset_57 ? args_5 : _GEN_6620; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6622 = 3'h6 == local_offset_57 ? args_6 : _GEN_6621; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6623 = 3'h2 == args_length_2 ? _GEN_6622 : _GEN_6615; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_58 = 3'h2 + args_offset_2; // @[executor.scala 222:61]
  wire [7:0] _GEN_6625 = 3'h1 == local_offset_58 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6626 = 3'h2 == local_offset_58 ? args_2 : _GEN_6625; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6627 = 3'h3 == local_offset_58 ? args_3 : _GEN_6626; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6628 = 3'h4 == local_offset_58 ? args_4 : _GEN_6627; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6629 = 3'h5 == local_offset_58 ? args_5 : _GEN_6628; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6630 = 3'h6 == local_offset_58 ? args_6 : _GEN_6629; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6631 = 3'h3 == args_length_2 ? _GEN_6630 : _GEN_6623; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_59 = 3'h3 + args_offset_2; // @[executor.scala 222:61]
  wire [7:0] _GEN_6633 = 3'h1 == local_offset_59 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6634 = 3'h2 == local_offset_59 ? args_2 : _GEN_6633; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6635 = 3'h3 == local_offset_59 ? args_3 : _GEN_6634; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6636 = 3'h4 == local_offset_59 ? args_4 : _GEN_6635; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6637 = 3'h5 == local_offset_59 ? args_5 : _GEN_6636; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6638 = 3'h6 == local_offset_59 ? args_6 : _GEN_6637; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6639 = 3'h4 == args_length_2 ? _GEN_6638 : _GEN_6631; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_60 = 3'h4 + args_offset_2; // @[executor.scala 222:61]
  wire [7:0] _GEN_6641 = 3'h1 == local_offset_60 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6642 = 3'h2 == local_offset_60 ? args_2 : _GEN_6641; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6643 = 3'h3 == local_offset_60 ? args_3 : _GEN_6642; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6644 = 3'h4 == local_offset_60 ? args_4 : _GEN_6643; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6645 = 3'h5 == local_offset_60 ? args_5 : _GEN_6644; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6646 = 3'h6 == local_offset_60 ? args_6 : _GEN_6645; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6647 = 3'h5 == args_length_2 ? _GEN_6646 : _GEN_6639; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_61 = 3'h5 + args_offset_2; // @[executor.scala 222:61]
  wire [7:0] _GEN_6649 = 3'h1 == local_offset_61 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6650 = 3'h2 == local_offset_61 ? args_2 : _GEN_6649; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6651 = 3'h3 == local_offset_61 ? args_3 : _GEN_6650; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6652 = 3'h4 == local_offset_61 ? args_4 : _GEN_6651; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6653 = 3'h5 == local_offset_61 ? args_5 : _GEN_6652; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6654 = 3'h6 == local_offset_61 ? args_6 : _GEN_6653; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6655 = 3'h6 == args_length_2 ? _GEN_6654 : _GEN_6647; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_62 = 3'h6 + args_offset_2; // @[executor.scala 222:61]
  wire [7:0] _GEN_6657 = 3'h1 == local_offset_62 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6658 = 3'h2 == local_offset_62 ? args_2 : _GEN_6657; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6659 = 3'h3 == local_offset_62 ? args_3 : _GEN_6658; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6660 = 3'h4 == local_offset_62 ? args_4 : _GEN_6659; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6661 = 3'h5 == local_offset_62 ? args_5 : _GEN_6660; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_6662 = 3'h6 == local_offset_62 ? args_6 : _GEN_6661; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] field_bytes_5_0 = 3'h7 == args_length_2 ? _GEN_6662 : _GEN_6655; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6671 = 3'h2 == args_length_2 ? _GEN_6614 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_6679 = 3'h3 == args_length_2 ? _GEN_6622 : _GEN_6671; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6687 = 3'h4 == args_length_2 ? _GEN_6630 : _GEN_6679; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6695 = 3'h5 == args_length_2 ? _GEN_6638 : _GEN_6687; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6703 = 3'h6 == args_length_2 ? _GEN_6646 : _GEN_6695; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6711 = 3'h7 == args_length_2 ? _GEN_6654 : _GEN_6703; // @[executor.scala 223:66 executor.scala 224:52]
  wire [3:0] _GEN_12207 = {{1'd0}, args_length_2}; // @[executor.scala 223:49]
  wire [7:0] field_bytes_5_1 = 4'h8 == _GEN_12207 ? _GEN_6662 : _GEN_6711; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6727 = 3'h3 == args_length_2 ? _GEN_6614 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_6735 = 3'h4 == args_length_2 ? _GEN_6622 : _GEN_6727; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6743 = 3'h5 == args_length_2 ? _GEN_6630 : _GEN_6735; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6751 = 3'h6 == args_length_2 ? _GEN_6638 : _GEN_6743; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6759 = 3'h7 == args_length_2 ? _GEN_6646 : _GEN_6751; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6767 = 4'h8 == _GEN_12207 ? _GEN_6654 : _GEN_6759; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_5_2 = 4'h9 == _GEN_12207 ? _GEN_6662 : _GEN_6767; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6783 = 3'h4 == args_length_2 ? _GEN_6614 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_6791 = 3'h5 == args_length_2 ? _GEN_6622 : _GEN_6783; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6799 = 3'h6 == args_length_2 ? _GEN_6630 : _GEN_6791; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6807 = 3'h7 == args_length_2 ? _GEN_6638 : _GEN_6799; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6815 = 4'h8 == _GEN_12207 ? _GEN_6646 : _GEN_6807; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_6823 = 4'h9 == _GEN_12207 ? _GEN_6654 : _GEN_6815; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_5_3 = 4'ha == _GEN_12207 ? _GEN_6662 : _GEN_6823; // @[executor.scala 223:66 executor.scala 224:52]
  wire [31:0] _io_field_out_2_T_1 = {field_bytes_5_0,field_bytes_5_1,field_bytes_5_2,field_bytes_5_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_6832 = 4'ha == opcode_2 ? _io_field_out_2_T_1 : 32'h0; // @[executor.scala 207:55 executor.scala 228:41 executor.scala 172:29]
  wire [17:0] io_field_out_2_hi_4 = io_field_out_2_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_2_T_4 = {io_field_out_2_hi_4,io_field_out_2_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_6833 = 4'hb == opcode_2 ? _io_field_out_2_T_4 : _GEN_6832; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_6834 = from_header_2 ? bias_2 : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_6835 = from_header_2 ? _io_field_out_2_T : _GEN_6833; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_6836 = from_header_2 ? _io_mask_out_2_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  wire [3:0] opcode_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] io_field_out_3_lo = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire  from_header_3 = length_3 != 8'h0; // @[executor.scala 177:45]
  wire [5:0] total_offset_hi_3 = offset_3[7:2]; // @[executor.scala 191:57]
  wire [7:0] _ending_T_7 = offset_3 + length_3; // @[executor.scala 193:46]
  wire [1:0] ending_3 = _ending_T_7[1:0]; // @[executor.scala 193:58]
  wire [3:0] _GEN_12213 = {{2'd0}, ending_3}; // @[executor.scala 194:45]
  wire [3:0] _bias_T_7 = 4'h4 - _GEN_12213; // @[executor.scala 194:45]
  wire [1:0] bias_3 = _bias_T_7[1:0]; // @[executor.scala 194:54]
  wire [7:0] total_offset_12 = {total_offset_hi_3,2'h0}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_6841 = 8'h1 == total_offset_12 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6842 = 8'h2 == total_offset_12 ? phv_data_2 : _GEN_6841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6843 = 8'h3 == total_offset_12 ? phv_data_3 : _GEN_6842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6844 = 8'h4 == total_offset_12 ? phv_data_4 : _GEN_6843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6845 = 8'h5 == total_offset_12 ? phv_data_5 : _GEN_6844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6846 = 8'h6 == total_offset_12 ? phv_data_6 : _GEN_6845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6847 = 8'h7 == total_offset_12 ? phv_data_7 : _GEN_6846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6848 = 8'h8 == total_offset_12 ? phv_data_8 : _GEN_6847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6849 = 8'h9 == total_offset_12 ? phv_data_9 : _GEN_6848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6850 = 8'ha == total_offset_12 ? phv_data_10 : _GEN_6849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6851 = 8'hb == total_offset_12 ? phv_data_11 : _GEN_6850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6852 = 8'hc == total_offset_12 ? phv_data_12 : _GEN_6851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6853 = 8'hd == total_offset_12 ? phv_data_13 : _GEN_6852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6854 = 8'he == total_offset_12 ? phv_data_14 : _GEN_6853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6855 = 8'hf == total_offset_12 ? phv_data_15 : _GEN_6854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6856 = 8'h10 == total_offset_12 ? phv_data_16 : _GEN_6855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6857 = 8'h11 == total_offset_12 ? phv_data_17 : _GEN_6856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6858 = 8'h12 == total_offset_12 ? phv_data_18 : _GEN_6857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6859 = 8'h13 == total_offset_12 ? phv_data_19 : _GEN_6858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6860 = 8'h14 == total_offset_12 ? phv_data_20 : _GEN_6859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6861 = 8'h15 == total_offset_12 ? phv_data_21 : _GEN_6860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6862 = 8'h16 == total_offset_12 ? phv_data_22 : _GEN_6861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6863 = 8'h17 == total_offset_12 ? phv_data_23 : _GEN_6862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6864 = 8'h18 == total_offset_12 ? phv_data_24 : _GEN_6863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6865 = 8'h19 == total_offset_12 ? phv_data_25 : _GEN_6864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6866 = 8'h1a == total_offset_12 ? phv_data_26 : _GEN_6865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6867 = 8'h1b == total_offset_12 ? phv_data_27 : _GEN_6866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6868 = 8'h1c == total_offset_12 ? phv_data_28 : _GEN_6867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6869 = 8'h1d == total_offset_12 ? phv_data_29 : _GEN_6868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6870 = 8'h1e == total_offset_12 ? phv_data_30 : _GEN_6869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6871 = 8'h1f == total_offset_12 ? phv_data_31 : _GEN_6870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6872 = 8'h20 == total_offset_12 ? phv_data_32 : _GEN_6871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6873 = 8'h21 == total_offset_12 ? phv_data_33 : _GEN_6872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6874 = 8'h22 == total_offset_12 ? phv_data_34 : _GEN_6873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6875 = 8'h23 == total_offset_12 ? phv_data_35 : _GEN_6874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6876 = 8'h24 == total_offset_12 ? phv_data_36 : _GEN_6875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6877 = 8'h25 == total_offset_12 ? phv_data_37 : _GEN_6876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6878 = 8'h26 == total_offset_12 ? phv_data_38 : _GEN_6877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6879 = 8'h27 == total_offset_12 ? phv_data_39 : _GEN_6878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6880 = 8'h28 == total_offset_12 ? phv_data_40 : _GEN_6879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6881 = 8'h29 == total_offset_12 ? phv_data_41 : _GEN_6880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6882 = 8'h2a == total_offset_12 ? phv_data_42 : _GEN_6881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6883 = 8'h2b == total_offset_12 ? phv_data_43 : _GEN_6882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6884 = 8'h2c == total_offset_12 ? phv_data_44 : _GEN_6883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6885 = 8'h2d == total_offset_12 ? phv_data_45 : _GEN_6884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6886 = 8'h2e == total_offset_12 ? phv_data_46 : _GEN_6885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6887 = 8'h2f == total_offset_12 ? phv_data_47 : _GEN_6886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6888 = 8'h30 == total_offset_12 ? phv_data_48 : _GEN_6887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6889 = 8'h31 == total_offset_12 ? phv_data_49 : _GEN_6888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6890 = 8'h32 == total_offset_12 ? phv_data_50 : _GEN_6889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6891 = 8'h33 == total_offset_12 ? phv_data_51 : _GEN_6890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6892 = 8'h34 == total_offset_12 ? phv_data_52 : _GEN_6891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6893 = 8'h35 == total_offset_12 ? phv_data_53 : _GEN_6892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6894 = 8'h36 == total_offset_12 ? phv_data_54 : _GEN_6893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6895 = 8'h37 == total_offset_12 ? phv_data_55 : _GEN_6894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6896 = 8'h38 == total_offset_12 ? phv_data_56 : _GEN_6895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6897 = 8'h39 == total_offset_12 ? phv_data_57 : _GEN_6896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6898 = 8'h3a == total_offset_12 ? phv_data_58 : _GEN_6897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6899 = 8'h3b == total_offset_12 ? phv_data_59 : _GEN_6898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6900 = 8'h3c == total_offset_12 ? phv_data_60 : _GEN_6899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6901 = 8'h3d == total_offset_12 ? phv_data_61 : _GEN_6900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6902 = 8'h3e == total_offset_12 ? phv_data_62 : _GEN_6901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6903 = 8'h3f == total_offset_12 ? phv_data_63 : _GEN_6902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6904 = 8'h40 == total_offset_12 ? phv_data_64 : _GEN_6903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6905 = 8'h41 == total_offset_12 ? phv_data_65 : _GEN_6904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6906 = 8'h42 == total_offset_12 ? phv_data_66 : _GEN_6905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6907 = 8'h43 == total_offset_12 ? phv_data_67 : _GEN_6906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6908 = 8'h44 == total_offset_12 ? phv_data_68 : _GEN_6907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6909 = 8'h45 == total_offset_12 ? phv_data_69 : _GEN_6908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6910 = 8'h46 == total_offset_12 ? phv_data_70 : _GEN_6909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6911 = 8'h47 == total_offset_12 ? phv_data_71 : _GEN_6910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6912 = 8'h48 == total_offset_12 ? phv_data_72 : _GEN_6911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6913 = 8'h49 == total_offset_12 ? phv_data_73 : _GEN_6912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6914 = 8'h4a == total_offset_12 ? phv_data_74 : _GEN_6913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6915 = 8'h4b == total_offset_12 ? phv_data_75 : _GEN_6914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6916 = 8'h4c == total_offset_12 ? phv_data_76 : _GEN_6915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6917 = 8'h4d == total_offset_12 ? phv_data_77 : _GEN_6916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6918 = 8'h4e == total_offset_12 ? phv_data_78 : _GEN_6917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6919 = 8'h4f == total_offset_12 ? phv_data_79 : _GEN_6918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6920 = 8'h50 == total_offset_12 ? phv_data_80 : _GEN_6919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6921 = 8'h51 == total_offset_12 ? phv_data_81 : _GEN_6920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6922 = 8'h52 == total_offset_12 ? phv_data_82 : _GEN_6921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6923 = 8'h53 == total_offset_12 ? phv_data_83 : _GEN_6922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6924 = 8'h54 == total_offset_12 ? phv_data_84 : _GEN_6923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6925 = 8'h55 == total_offset_12 ? phv_data_85 : _GEN_6924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6926 = 8'h56 == total_offset_12 ? phv_data_86 : _GEN_6925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6927 = 8'h57 == total_offset_12 ? phv_data_87 : _GEN_6926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6928 = 8'h58 == total_offset_12 ? phv_data_88 : _GEN_6927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6929 = 8'h59 == total_offset_12 ? phv_data_89 : _GEN_6928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6930 = 8'h5a == total_offset_12 ? phv_data_90 : _GEN_6929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6931 = 8'h5b == total_offset_12 ? phv_data_91 : _GEN_6930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6932 = 8'h5c == total_offset_12 ? phv_data_92 : _GEN_6931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6933 = 8'h5d == total_offset_12 ? phv_data_93 : _GEN_6932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6934 = 8'h5e == total_offset_12 ? phv_data_94 : _GEN_6933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6935 = 8'h5f == total_offset_12 ? phv_data_95 : _GEN_6934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6936 = 8'h60 == total_offset_12 ? phv_data_96 : _GEN_6935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6937 = 8'h61 == total_offset_12 ? phv_data_97 : _GEN_6936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6938 = 8'h62 == total_offset_12 ? phv_data_98 : _GEN_6937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6939 = 8'h63 == total_offset_12 ? phv_data_99 : _GEN_6938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6940 = 8'h64 == total_offset_12 ? phv_data_100 : _GEN_6939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6941 = 8'h65 == total_offset_12 ? phv_data_101 : _GEN_6940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6942 = 8'h66 == total_offset_12 ? phv_data_102 : _GEN_6941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6943 = 8'h67 == total_offset_12 ? phv_data_103 : _GEN_6942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6944 = 8'h68 == total_offset_12 ? phv_data_104 : _GEN_6943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6945 = 8'h69 == total_offset_12 ? phv_data_105 : _GEN_6944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6946 = 8'h6a == total_offset_12 ? phv_data_106 : _GEN_6945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6947 = 8'h6b == total_offset_12 ? phv_data_107 : _GEN_6946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6948 = 8'h6c == total_offset_12 ? phv_data_108 : _GEN_6947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6949 = 8'h6d == total_offset_12 ? phv_data_109 : _GEN_6948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6950 = 8'h6e == total_offset_12 ? phv_data_110 : _GEN_6949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6951 = 8'h6f == total_offset_12 ? phv_data_111 : _GEN_6950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6952 = 8'h70 == total_offset_12 ? phv_data_112 : _GEN_6951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6953 = 8'h71 == total_offset_12 ? phv_data_113 : _GEN_6952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6954 = 8'h72 == total_offset_12 ? phv_data_114 : _GEN_6953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6955 = 8'h73 == total_offset_12 ? phv_data_115 : _GEN_6954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6956 = 8'h74 == total_offset_12 ? phv_data_116 : _GEN_6955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6957 = 8'h75 == total_offset_12 ? phv_data_117 : _GEN_6956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6958 = 8'h76 == total_offset_12 ? phv_data_118 : _GEN_6957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6959 = 8'h77 == total_offset_12 ? phv_data_119 : _GEN_6958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6960 = 8'h78 == total_offset_12 ? phv_data_120 : _GEN_6959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6961 = 8'h79 == total_offset_12 ? phv_data_121 : _GEN_6960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6962 = 8'h7a == total_offset_12 ? phv_data_122 : _GEN_6961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6963 = 8'h7b == total_offset_12 ? phv_data_123 : _GEN_6962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6964 = 8'h7c == total_offset_12 ? phv_data_124 : _GEN_6963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6965 = 8'h7d == total_offset_12 ? phv_data_125 : _GEN_6964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6966 = 8'h7e == total_offset_12 ? phv_data_126 : _GEN_6965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6967 = 8'h7f == total_offset_12 ? phv_data_127 : _GEN_6966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6968 = 8'h80 == total_offset_12 ? phv_data_128 : _GEN_6967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6969 = 8'h81 == total_offset_12 ? phv_data_129 : _GEN_6968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6970 = 8'h82 == total_offset_12 ? phv_data_130 : _GEN_6969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6971 = 8'h83 == total_offset_12 ? phv_data_131 : _GEN_6970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6972 = 8'h84 == total_offset_12 ? phv_data_132 : _GEN_6971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6973 = 8'h85 == total_offset_12 ? phv_data_133 : _GEN_6972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6974 = 8'h86 == total_offset_12 ? phv_data_134 : _GEN_6973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6975 = 8'h87 == total_offset_12 ? phv_data_135 : _GEN_6974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6976 = 8'h88 == total_offset_12 ? phv_data_136 : _GEN_6975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6977 = 8'h89 == total_offset_12 ? phv_data_137 : _GEN_6976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6978 = 8'h8a == total_offset_12 ? phv_data_138 : _GEN_6977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6979 = 8'h8b == total_offset_12 ? phv_data_139 : _GEN_6978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6980 = 8'h8c == total_offset_12 ? phv_data_140 : _GEN_6979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6981 = 8'h8d == total_offset_12 ? phv_data_141 : _GEN_6980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6982 = 8'h8e == total_offset_12 ? phv_data_142 : _GEN_6981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6983 = 8'h8f == total_offset_12 ? phv_data_143 : _GEN_6982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6984 = 8'h90 == total_offset_12 ? phv_data_144 : _GEN_6983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6985 = 8'h91 == total_offset_12 ? phv_data_145 : _GEN_6984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6986 = 8'h92 == total_offset_12 ? phv_data_146 : _GEN_6985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6987 = 8'h93 == total_offset_12 ? phv_data_147 : _GEN_6986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6988 = 8'h94 == total_offset_12 ? phv_data_148 : _GEN_6987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6989 = 8'h95 == total_offset_12 ? phv_data_149 : _GEN_6988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6990 = 8'h96 == total_offset_12 ? phv_data_150 : _GEN_6989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6991 = 8'h97 == total_offset_12 ? phv_data_151 : _GEN_6990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6992 = 8'h98 == total_offset_12 ? phv_data_152 : _GEN_6991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6993 = 8'h99 == total_offset_12 ? phv_data_153 : _GEN_6992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6994 = 8'h9a == total_offset_12 ? phv_data_154 : _GEN_6993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6995 = 8'h9b == total_offset_12 ? phv_data_155 : _GEN_6994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6996 = 8'h9c == total_offset_12 ? phv_data_156 : _GEN_6995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6997 = 8'h9d == total_offset_12 ? phv_data_157 : _GEN_6996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6998 = 8'h9e == total_offset_12 ? phv_data_158 : _GEN_6997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_6999 = 8'h9f == total_offset_12 ? phv_data_159 : _GEN_6998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7000 = 8'ha0 == total_offset_12 ? phv_data_160 : _GEN_6999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7001 = 8'ha1 == total_offset_12 ? phv_data_161 : _GEN_7000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7002 = 8'ha2 == total_offset_12 ? phv_data_162 : _GEN_7001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7003 = 8'ha3 == total_offset_12 ? phv_data_163 : _GEN_7002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7004 = 8'ha4 == total_offset_12 ? phv_data_164 : _GEN_7003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7005 = 8'ha5 == total_offset_12 ? phv_data_165 : _GEN_7004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7006 = 8'ha6 == total_offset_12 ? phv_data_166 : _GEN_7005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7007 = 8'ha7 == total_offset_12 ? phv_data_167 : _GEN_7006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7008 = 8'ha8 == total_offset_12 ? phv_data_168 : _GEN_7007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7009 = 8'ha9 == total_offset_12 ? phv_data_169 : _GEN_7008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7010 = 8'haa == total_offset_12 ? phv_data_170 : _GEN_7009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7011 = 8'hab == total_offset_12 ? phv_data_171 : _GEN_7010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7012 = 8'hac == total_offset_12 ? phv_data_172 : _GEN_7011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7013 = 8'had == total_offset_12 ? phv_data_173 : _GEN_7012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7014 = 8'hae == total_offset_12 ? phv_data_174 : _GEN_7013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7015 = 8'haf == total_offset_12 ? phv_data_175 : _GEN_7014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7016 = 8'hb0 == total_offset_12 ? phv_data_176 : _GEN_7015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7017 = 8'hb1 == total_offset_12 ? phv_data_177 : _GEN_7016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7018 = 8'hb2 == total_offset_12 ? phv_data_178 : _GEN_7017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7019 = 8'hb3 == total_offset_12 ? phv_data_179 : _GEN_7018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7020 = 8'hb4 == total_offset_12 ? phv_data_180 : _GEN_7019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7021 = 8'hb5 == total_offset_12 ? phv_data_181 : _GEN_7020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7022 = 8'hb6 == total_offset_12 ? phv_data_182 : _GEN_7021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7023 = 8'hb7 == total_offset_12 ? phv_data_183 : _GEN_7022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7024 = 8'hb8 == total_offset_12 ? phv_data_184 : _GEN_7023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7025 = 8'hb9 == total_offset_12 ? phv_data_185 : _GEN_7024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7026 = 8'hba == total_offset_12 ? phv_data_186 : _GEN_7025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7027 = 8'hbb == total_offset_12 ? phv_data_187 : _GEN_7026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7028 = 8'hbc == total_offset_12 ? phv_data_188 : _GEN_7027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7029 = 8'hbd == total_offset_12 ? phv_data_189 : _GEN_7028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7030 = 8'hbe == total_offset_12 ? phv_data_190 : _GEN_7029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7031 = 8'hbf == total_offset_12 ? phv_data_191 : _GEN_7030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7032 = 8'hc0 == total_offset_12 ? phv_data_192 : _GEN_7031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7033 = 8'hc1 == total_offset_12 ? phv_data_193 : _GEN_7032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7034 = 8'hc2 == total_offset_12 ? phv_data_194 : _GEN_7033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7035 = 8'hc3 == total_offset_12 ? phv_data_195 : _GEN_7034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7036 = 8'hc4 == total_offset_12 ? phv_data_196 : _GEN_7035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7037 = 8'hc5 == total_offset_12 ? phv_data_197 : _GEN_7036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7038 = 8'hc6 == total_offset_12 ? phv_data_198 : _GEN_7037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7039 = 8'hc7 == total_offset_12 ? phv_data_199 : _GEN_7038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7040 = 8'hc8 == total_offset_12 ? phv_data_200 : _GEN_7039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7041 = 8'hc9 == total_offset_12 ? phv_data_201 : _GEN_7040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7042 = 8'hca == total_offset_12 ? phv_data_202 : _GEN_7041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7043 = 8'hcb == total_offset_12 ? phv_data_203 : _GEN_7042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7044 = 8'hcc == total_offset_12 ? phv_data_204 : _GEN_7043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7045 = 8'hcd == total_offset_12 ? phv_data_205 : _GEN_7044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7046 = 8'hce == total_offset_12 ? phv_data_206 : _GEN_7045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7047 = 8'hcf == total_offset_12 ? phv_data_207 : _GEN_7046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7048 = 8'hd0 == total_offset_12 ? phv_data_208 : _GEN_7047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7049 = 8'hd1 == total_offset_12 ? phv_data_209 : _GEN_7048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7050 = 8'hd2 == total_offset_12 ? phv_data_210 : _GEN_7049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7051 = 8'hd3 == total_offset_12 ? phv_data_211 : _GEN_7050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7052 = 8'hd4 == total_offset_12 ? phv_data_212 : _GEN_7051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7053 = 8'hd5 == total_offset_12 ? phv_data_213 : _GEN_7052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7054 = 8'hd6 == total_offset_12 ? phv_data_214 : _GEN_7053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7055 = 8'hd7 == total_offset_12 ? phv_data_215 : _GEN_7054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7056 = 8'hd8 == total_offset_12 ? phv_data_216 : _GEN_7055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7057 = 8'hd9 == total_offset_12 ? phv_data_217 : _GEN_7056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7058 = 8'hda == total_offset_12 ? phv_data_218 : _GEN_7057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7059 = 8'hdb == total_offset_12 ? phv_data_219 : _GEN_7058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7060 = 8'hdc == total_offset_12 ? phv_data_220 : _GEN_7059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7061 = 8'hdd == total_offset_12 ? phv_data_221 : _GEN_7060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7062 = 8'hde == total_offset_12 ? phv_data_222 : _GEN_7061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7063 = 8'hdf == total_offset_12 ? phv_data_223 : _GEN_7062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7064 = 8'he0 == total_offset_12 ? phv_data_224 : _GEN_7063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7065 = 8'he1 == total_offset_12 ? phv_data_225 : _GEN_7064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7066 = 8'he2 == total_offset_12 ? phv_data_226 : _GEN_7065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7067 = 8'he3 == total_offset_12 ? phv_data_227 : _GEN_7066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7068 = 8'he4 == total_offset_12 ? phv_data_228 : _GEN_7067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7069 = 8'he5 == total_offset_12 ? phv_data_229 : _GEN_7068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7070 = 8'he6 == total_offset_12 ? phv_data_230 : _GEN_7069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7071 = 8'he7 == total_offset_12 ? phv_data_231 : _GEN_7070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7072 = 8'he8 == total_offset_12 ? phv_data_232 : _GEN_7071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7073 = 8'he9 == total_offset_12 ? phv_data_233 : _GEN_7072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7074 = 8'hea == total_offset_12 ? phv_data_234 : _GEN_7073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7075 = 8'heb == total_offset_12 ? phv_data_235 : _GEN_7074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7076 = 8'hec == total_offset_12 ? phv_data_236 : _GEN_7075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7077 = 8'hed == total_offset_12 ? phv_data_237 : _GEN_7076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7078 = 8'hee == total_offset_12 ? phv_data_238 : _GEN_7077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7079 = 8'hef == total_offset_12 ? phv_data_239 : _GEN_7078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7080 = 8'hf0 == total_offset_12 ? phv_data_240 : _GEN_7079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7081 = 8'hf1 == total_offset_12 ? phv_data_241 : _GEN_7080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7082 = 8'hf2 == total_offset_12 ? phv_data_242 : _GEN_7081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7083 = 8'hf3 == total_offset_12 ? phv_data_243 : _GEN_7082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7084 = 8'hf4 == total_offset_12 ? phv_data_244 : _GEN_7083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7085 = 8'hf5 == total_offset_12 ? phv_data_245 : _GEN_7084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7086 = 8'hf6 == total_offset_12 ? phv_data_246 : _GEN_7085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7087 = 8'hf7 == total_offset_12 ? phv_data_247 : _GEN_7086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7088 = 8'hf8 == total_offset_12 ? phv_data_248 : _GEN_7087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7089 = 8'hf9 == total_offset_12 ? phv_data_249 : _GEN_7088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7090 = 8'hfa == total_offset_12 ? phv_data_250 : _GEN_7089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7091 = 8'hfb == total_offset_12 ? phv_data_251 : _GEN_7090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7092 = 8'hfc == total_offset_12 ? phv_data_252 : _GEN_7091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7093 = 8'hfd == total_offset_12 ? phv_data_253 : _GEN_7092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7094 = 8'hfe == total_offset_12 ? phv_data_254 : _GEN_7093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7095 = 8'hff == total_offset_12 ? phv_data_255 : _GEN_7094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_12214 = {{1'd0}, total_offset_12}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7096 = 9'h100 == _GEN_12214 ? phv_data_256 : _GEN_7095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7097 = 9'h101 == _GEN_12214 ? phv_data_257 : _GEN_7096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7098 = 9'h102 == _GEN_12214 ? phv_data_258 : _GEN_7097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7099 = 9'h103 == _GEN_12214 ? phv_data_259 : _GEN_7098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7100 = 9'h104 == _GEN_12214 ? phv_data_260 : _GEN_7099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7101 = 9'h105 == _GEN_12214 ? phv_data_261 : _GEN_7100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7102 = 9'h106 == _GEN_12214 ? phv_data_262 : _GEN_7101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7103 = 9'h107 == _GEN_12214 ? phv_data_263 : _GEN_7102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7104 = 9'h108 == _GEN_12214 ? phv_data_264 : _GEN_7103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7105 = 9'h109 == _GEN_12214 ? phv_data_265 : _GEN_7104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7106 = 9'h10a == _GEN_12214 ? phv_data_266 : _GEN_7105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7107 = 9'h10b == _GEN_12214 ? phv_data_267 : _GEN_7106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7108 = 9'h10c == _GEN_12214 ? phv_data_268 : _GEN_7107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7109 = 9'h10d == _GEN_12214 ? phv_data_269 : _GEN_7108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7110 = 9'h10e == _GEN_12214 ? phv_data_270 : _GEN_7109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7111 = 9'h10f == _GEN_12214 ? phv_data_271 : _GEN_7110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7112 = 9'h110 == _GEN_12214 ? phv_data_272 : _GEN_7111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7113 = 9'h111 == _GEN_12214 ? phv_data_273 : _GEN_7112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7114 = 9'h112 == _GEN_12214 ? phv_data_274 : _GEN_7113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7115 = 9'h113 == _GEN_12214 ? phv_data_275 : _GEN_7114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7116 = 9'h114 == _GEN_12214 ? phv_data_276 : _GEN_7115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7117 = 9'h115 == _GEN_12214 ? phv_data_277 : _GEN_7116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7118 = 9'h116 == _GEN_12214 ? phv_data_278 : _GEN_7117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7119 = 9'h117 == _GEN_12214 ? phv_data_279 : _GEN_7118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7120 = 9'h118 == _GEN_12214 ? phv_data_280 : _GEN_7119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7121 = 9'h119 == _GEN_12214 ? phv_data_281 : _GEN_7120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7122 = 9'h11a == _GEN_12214 ? phv_data_282 : _GEN_7121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7123 = 9'h11b == _GEN_12214 ? phv_data_283 : _GEN_7122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7124 = 9'h11c == _GEN_12214 ? phv_data_284 : _GEN_7123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7125 = 9'h11d == _GEN_12214 ? phv_data_285 : _GEN_7124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7126 = 9'h11e == _GEN_12214 ? phv_data_286 : _GEN_7125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7127 = 9'h11f == _GEN_12214 ? phv_data_287 : _GEN_7126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7128 = 9'h120 == _GEN_12214 ? phv_data_288 : _GEN_7127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7129 = 9'h121 == _GEN_12214 ? phv_data_289 : _GEN_7128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7130 = 9'h122 == _GEN_12214 ? phv_data_290 : _GEN_7129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7131 = 9'h123 == _GEN_12214 ? phv_data_291 : _GEN_7130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7132 = 9'h124 == _GEN_12214 ? phv_data_292 : _GEN_7131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7133 = 9'h125 == _GEN_12214 ? phv_data_293 : _GEN_7132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7134 = 9'h126 == _GEN_12214 ? phv_data_294 : _GEN_7133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7135 = 9'h127 == _GEN_12214 ? phv_data_295 : _GEN_7134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7136 = 9'h128 == _GEN_12214 ? phv_data_296 : _GEN_7135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7137 = 9'h129 == _GEN_12214 ? phv_data_297 : _GEN_7136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7138 = 9'h12a == _GEN_12214 ? phv_data_298 : _GEN_7137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7139 = 9'h12b == _GEN_12214 ? phv_data_299 : _GEN_7138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7140 = 9'h12c == _GEN_12214 ? phv_data_300 : _GEN_7139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7141 = 9'h12d == _GEN_12214 ? phv_data_301 : _GEN_7140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7142 = 9'h12e == _GEN_12214 ? phv_data_302 : _GEN_7141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7143 = 9'h12f == _GEN_12214 ? phv_data_303 : _GEN_7142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7144 = 9'h130 == _GEN_12214 ? phv_data_304 : _GEN_7143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7145 = 9'h131 == _GEN_12214 ? phv_data_305 : _GEN_7144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7146 = 9'h132 == _GEN_12214 ? phv_data_306 : _GEN_7145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7147 = 9'h133 == _GEN_12214 ? phv_data_307 : _GEN_7146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7148 = 9'h134 == _GEN_12214 ? phv_data_308 : _GEN_7147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7149 = 9'h135 == _GEN_12214 ? phv_data_309 : _GEN_7148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7150 = 9'h136 == _GEN_12214 ? phv_data_310 : _GEN_7149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7151 = 9'h137 == _GEN_12214 ? phv_data_311 : _GEN_7150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7152 = 9'h138 == _GEN_12214 ? phv_data_312 : _GEN_7151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7153 = 9'h139 == _GEN_12214 ? phv_data_313 : _GEN_7152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7154 = 9'h13a == _GEN_12214 ? phv_data_314 : _GEN_7153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7155 = 9'h13b == _GEN_12214 ? phv_data_315 : _GEN_7154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7156 = 9'h13c == _GEN_12214 ? phv_data_316 : _GEN_7155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7157 = 9'h13d == _GEN_12214 ? phv_data_317 : _GEN_7156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7158 = 9'h13e == _GEN_12214 ? phv_data_318 : _GEN_7157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7159 = 9'h13f == _GEN_12214 ? phv_data_319 : _GEN_7158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7160 = 9'h140 == _GEN_12214 ? phv_data_320 : _GEN_7159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7161 = 9'h141 == _GEN_12214 ? phv_data_321 : _GEN_7160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7162 = 9'h142 == _GEN_12214 ? phv_data_322 : _GEN_7161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7163 = 9'h143 == _GEN_12214 ? phv_data_323 : _GEN_7162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7164 = 9'h144 == _GEN_12214 ? phv_data_324 : _GEN_7163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7165 = 9'h145 == _GEN_12214 ? phv_data_325 : _GEN_7164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7166 = 9'h146 == _GEN_12214 ? phv_data_326 : _GEN_7165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7167 = 9'h147 == _GEN_12214 ? phv_data_327 : _GEN_7166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7168 = 9'h148 == _GEN_12214 ? phv_data_328 : _GEN_7167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7169 = 9'h149 == _GEN_12214 ? phv_data_329 : _GEN_7168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7170 = 9'h14a == _GEN_12214 ? phv_data_330 : _GEN_7169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7171 = 9'h14b == _GEN_12214 ? phv_data_331 : _GEN_7170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7172 = 9'h14c == _GEN_12214 ? phv_data_332 : _GEN_7171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7173 = 9'h14d == _GEN_12214 ? phv_data_333 : _GEN_7172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7174 = 9'h14e == _GEN_12214 ? phv_data_334 : _GEN_7173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7175 = 9'h14f == _GEN_12214 ? phv_data_335 : _GEN_7174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7176 = 9'h150 == _GEN_12214 ? phv_data_336 : _GEN_7175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7177 = 9'h151 == _GEN_12214 ? phv_data_337 : _GEN_7176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7178 = 9'h152 == _GEN_12214 ? phv_data_338 : _GEN_7177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7179 = 9'h153 == _GEN_12214 ? phv_data_339 : _GEN_7178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7180 = 9'h154 == _GEN_12214 ? phv_data_340 : _GEN_7179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7181 = 9'h155 == _GEN_12214 ? phv_data_341 : _GEN_7180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7182 = 9'h156 == _GEN_12214 ? phv_data_342 : _GEN_7181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7183 = 9'h157 == _GEN_12214 ? phv_data_343 : _GEN_7182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7184 = 9'h158 == _GEN_12214 ? phv_data_344 : _GEN_7183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7185 = 9'h159 == _GEN_12214 ? phv_data_345 : _GEN_7184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7186 = 9'h15a == _GEN_12214 ? phv_data_346 : _GEN_7185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7187 = 9'h15b == _GEN_12214 ? phv_data_347 : _GEN_7186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7188 = 9'h15c == _GEN_12214 ? phv_data_348 : _GEN_7187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7189 = 9'h15d == _GEN_12214 ? phv_data_349 : _GEN_7188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7190 = 9'h15e == _GEN_12214 ? phv_data_350 : _GEN_7189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7191 = 9'h15f == _GEN_12214 ? phv_data_351 : _GEN_7190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7192 = 9'h160 == _GEN_12214 ? phv_data_352 : _GEN_7191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7193 = 9'h161 == _GEN_12214 ? phv_data_353 : _GEN_7192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7194 = 9'h162 == _GEN_12214 ? phv_data_354 : _GEN_7193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7195 = 9'h163 == _GEN_12214 ? phv_data_355 : _GEN_7194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7196 = 9'h164 == _GEN_12214 ? phv_data_356 : _GEN_7195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7197 = 9'h165 == _GEN_12214 ? phv_data_357 : _GEN_7196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7198 = 9'h166 == _GEN_12214 ? phv_data_358 : _GEN_7197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7199 = 9'h167 == _GEN_12214 ? phv_data_359 : _GEN_7198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7200 = 9'h168 == _GEN_12214 ? phv_data_360 : _GEN_7199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7201 = 9'h169 == _GEN_12214 ? phv_data_361 : _GEN_7200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7202 = 9'h16a == _GEN_12214 ? phv_data_362 : _GEN_7201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7203 = 9'h16b == _GEN_12214 ? phv_data_363 : _GEN_7202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7204 = 9'h16c == _GEN_12214 ? phv_data_364 : _GEN_7203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7205 = 9'h16d == _GEN_12214 ? phv_data_365 : _GEN_7204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7206 = 9'h16e == _GEN_12214 ? phv_data_366 : _GEN_7205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7207 = 9'h16f == _GEN_12214 ? phv_data_367 : _GEN_7206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7208 = 9'h170 == _GEN_12214 ? phv_data_368 : _GEN_7207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7209 = 9'h171 == _GEN_12214 ? phv_data_369 : _GEN_7208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7210 = 9'h172 == _GEN_12214 ? phv_data_370 : _GEN_7209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7211 = 9'h173 == _GEN_12214 ? phv_data_371 : _GEN_7210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7212 = 9'h174 == _GEN_12214 ? phv_data_372 : _GEN_7211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7213 = 9'h175 == _GEN_12214 ? phv_data_373 : _GEN_7212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7214 = 9'h176 == _GEN_12214 ? phv_data_374 : _GEN_7213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7215 = 9'h177 == _GEN_12214 ? phv_data_375 : _GEN_7214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7216 = 9'h178 == _GEN_12214 ? phv_data_376 : _GEN_7215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7217 = 9'h179 == _GEN_12214 ? phv_data_377 : _GEN_7216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7218 = 9'h17a == _GEN_12214 ? phv_data_378 : _GEN_7217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7219 = 9'h17b == _GEN_12214 ? phv_data_379 : _GEN_7218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7220 = 9'h17c == _GEN_12214 ? phv_data_380 : _GEN_7219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7221 = 9'h17d == _GEN_12214 ? phv_data_381 : _GEN_7220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7222 = 9'h17e == _GEN_12214 ? phv_data_382 : _GEN_7221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7223 = 9'h17f == _GEN_12214 ? phv_data_383 : _GEN_7222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7224 = 9'h180 == _GEN_12214 ? phv_data_384 : _GEN_7223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7225 = 9'h181 == _GEN_12214 ? phv_data_385 : _GEN_7224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7226 = 9'h182 == _GEN_12214 ? phv_data_386 : _GEN_7225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7227 = 9'h183 == _GEN_12214 ? phv_data_387 : _GEN_7226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7228 = 9'h184 == _GEN_12214 ? phv_data_388 : _GEN_7227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7229 = 9'h185 == _GEN_12214 ? phv_data_389 : _GEN_7228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7230 = 9'h186 == _GEN_12214 ? phv_data_390 : _GEN_7229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7231 = 9'h187 == _GEN_12214 ? phv_data_391 : _GEN_7230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7232 = 9'h188 == _GEN_12214 ? phv_data_392 : _GEN_7231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7233 = 9'h189 == _GEN_12214 ? phv_data_393 : _GEN_7232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7234 = 9'h18a == _GEN_12214 ? phv_data_394 : _GEN_7233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7235 = 9'h18b == _GEN_12214 ? phv_data_395 : _GEN_7234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7236 = 9'h18c == _GEN_12214 ? phv_data_396 : _GEN_7235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7237 = 9'h18d == _GEN_12214 ? phv_data_397 : _GEN_7236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7238 = 9'h18e == _GEN_12214 ? phv_data_398 : _GEN_7237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7239 = 9'h18f == _GEN_12214 ? phv_data_399 : _GEN_7238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7240 = 9'h190 == _GEN_12214 ? phv_data_400 : _GEN_7239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7241 = 9'h191 == _GEN_12214 ? phv_data_401 : _GEN_7240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7242 = 9'h192 == _GEN_12214 ? phv_data_402 : _GEN_7241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7243 = 9'h193 == _GEN_12214 ? phv_data_403 : _GEN_7242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7244 = 9'h194 == _GEN_12214 ? phv_data_404 : _GEN_7243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7245 = 9'h195 == _GEN_12214 ? phv_data_405 : _GEN_7244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7246 = 9'h196 == _GEN_12214 ? phv_data_406 : _GEN_7245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7247 = 9'h197 == _GEN_12214 ? phv_data_407 : _GEN_7246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7248 = 9'h198 == _GEN_12214 ? phv_data_408 : _GEN_7247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7249 = 9'h199 == _GEN_12214 ? phv_data_409 : _GEN_7248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7250 = 9'h19a == _GEN_12214 ? phv_data_410 : _GEN_7249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7251 = 9'h19b == _GEN_12214 ? phv_data_411 : _GEN_7250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7252 = 9'h19c == _GEN_12214 ? phv_data_412 : _GEN_7251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7253 = 9'h19d == _GEN_12214 ? phv_data_413 : _GEN_7252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7254 = 9'h19e == _GEN_12214 ? phv_data_414 : _GEN_7253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7255 = 9'h19f == _GEN_12214 ? phv_data_415 : _GEN_7254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7256 = 9'h1a0 == _GEN_12214 ? phv_data_416 : _GEN_7255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7257 = 9'h1a1 == _GEN_12214 ? phv_data_417 : _GEN_7256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7258 = 9'h1a2 == _GEN_12214 ? phv_data_418 : _GEN_7257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7259 = 9'h1a3 == _GEN_12214 ? phv_data_419 : _GEN_7258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7260 = 9'h1a4 == _GEN_12214 ? phv_data_420 : _GEN_7259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7261 = 9'h1a5 == _GEN_12214 ? phv_data_421 : _GEN_7260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7262 = 9'h1a6 == _GEN_12214 ? phv_data_422 : _GEN_7261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7263 = 9'h1a7 == _GEN_12214 ? phv_data_423 : _GEN_7262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7264 = 9'h1a8 == _GEN_12214 ? phv_data_424 : _GEN_7263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7265 = 9'h1a9 == _GEN_12214 ? phv_data_425 : _GEN_7264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7266 = 9'h1aa == _GEN_12214 ? phv_data_426 : _GEN_7265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7267 = 9'h1ab == _GEN_12214 ? phv_data_427 : _GEN_7266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7268 = 9'h1ac == _GEN_12214 ? phv_data_428 : _GEN_7267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7269 = 9'h1ad == _GEN_12214 ? phv_data_429 : _GEN_7268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7270 = 9'h1ae == _GEN_12214 ? phv_data_430 : _GEN_7269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7271 = 9'h1af == _GEN_12214 ? phv_data_431 : _GEN_7270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7272 = 9'h1b0 == _GEN_12214 ? phv_data_432 : _GEN_7271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7273 = 9'h1b1 == _GEN_12214 ? phv_data_433 : _GEN_7272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7274 = 9'h1b2 == _GEN_12214 ? phv_data_434 : _GEN_7273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7275 = 9'h1b3 == _GEN_12214 ? phv_data_435 : _GEN_7274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7276 = 9'h1b4 == _GEN_12214 ? phv_data_436 : _GEN_7275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7277 = 9'h1b5 == _GEN_12214 ? phv_data_437 : _GEN_7276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7278 = 9'h1b6 == _GEN_12214 ? phv_data_438 : _GEN_7277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7279 = 9'h1b7 == _GEN_12214 ? phv_data_439 : _GEN_7278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7280 = 9'h1b8 == _GEN_12214 ? phv_data_440 : _GEN_7279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7281 = 9'h1b9 == _GEN_12214 ? phv_data_441 : _GEN_7280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7282 = 9'h1ba == _GEN_12214 ? phv_data_442 : _GEN_7281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7283 = 9'h1bb == _GEN_12214 ? phv_data_443 : _GEN_7282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7284 = 9'h1bc == _GEN_12214 ? phv_data_444 : _GEN_7283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7285 = 9'h1bd == _GEN_12214 ? phv_data_445 : _GEN_7284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7286 = 9'h1be == _GEN_12214 ? phv_data_446 : _GEN_7285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7287 = 9'h1bf == _GEN_12214 ? phv_data_447 : _GEN_7286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7288 = 9'h1c0 == _GEN_12214 ? phv_data_448 : _GEN_7287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7289 = 9'h1c1 == _GEN_12214 ? phv_data_449 : _GEN_7288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7290 = 9'h1c2 == _GEN_12214 ? phv_data_450 : _GEN_7289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7291 = 9'h1c3 == _GEN_12214 ? phv_data_451 : _GEN_7290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7292 = 9'h1c4 == _GEN_12214 ? phv_data_452 : _GEN_7291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7293 = 9'h1c5 == _GEN_12214 ? phv_data_453 : _GEN_7292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7294 = 9'h1c6 == _GEN_12214 ? phv_data_454 : _GEN_7293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7295 = 9'h1c7 == _GEN_12214 ? phv_data_455 : _GEN_7294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7296 = 9'h1c8 == _GEN_12214 ? phv_data_456 : _GEN_7295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7297 = 9'h1c9 == _GEN_12214 ? phv_data_457 : _GEN_7296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7298 = 9'h1ca == _GEN_12214 ? phv_data_458 : _GEN_7297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7299 = 9'h1cb == _GEN_12214 ? phv_data_459 : _GEN_7298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7300 = 9'h1cc == _GEN_12214 ? phv_data_460 : _GEN_7299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7301 = 9'h1cd == _GEN_12214 ? phv_data_461 : _GEN_7300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7302 = 9'h1ce == _GEN_12214 ? phv_data_462 : _GEN_7301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7303 = 9'h1cf == _GEN_12214 ? phv_data_463 : _GEN_7302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7304 = 9'h1d0 == _GEN_12214 ? phv_data_464 : _GEN_7303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7305 = 9'h1d1 == _GEN_12214 ? phv_data_465 : _GEN_7304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7306 = 9'h1d2 == _GEN_12214 ? phv_data_466 : _GEN_7305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7307 = 9'h1d3 == _GEN_12214 ? phv_data_467 : _GEN_7306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7308 = 9'h1d4 == _GEN_12214 ? phv_data_468 : _GEN_7307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7309 = 9'h1d5 == _GEN_12214 ? phv_data_469 : _GEN_7308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7310 = 9'h1d6 == _GEN_12214 ? phv_data_470 : _GEN_7309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7311 = 9'h1d7 == _GEN_12214 ? phv_data_471 : _GEN_7310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7312 = 9'h1d8 == _GEN_12214 ? phv_data_472 : _GEN_7311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7313 = 9'h1d9 == _GEN_12214 ? phv_data_473 : _GEN_7312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7314 = 9'h1da == _GEN_12214 ? phv_data_474 : _GEN_7313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7315 = 9'h1db == _GEN_12214 ? phv_data_475 : _GEN_7314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7316 = 9'h1dc == _GEN_12214 ? phv_data_476 : _GEN_7315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7317 = 9'h1dd == _GEN_12214 ? phv_data_477 : _GEN_7316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7318 = 9'h1de == _GEN_12214 ? phv_data_478 : _GEN_7317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7319 = 9'h1df == _GEN_12214 ? phv_data_479 : _GEN_7318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7320 = 9'h1e0 == _GEN_12214 ? phv_data_480 : _GEN_7319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7321 = 9'h1e1 == _GEN_12214 ? phv_data_481 : _GEN_7320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7322 = 9'h1e2 == _GEN_12214 ? phv_data_482 : _GEN_7321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7323 = 9'h1e3 == _GEN_12214 ? phv_data_483 : _GEN_7322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7324 = 9'h1e4 == _GEN_12214 ? phv_data_484 : _GEN_7323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7325 = 9'h1e5 == _GEN_12214 ? phv_data_485 : _GEN_7324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7326 = 9'h1e6 == _GEN_12214 ? phv_data_486 : _GEN_7325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7327 = 9'h1e7 == _GEN_12214 ? phv_data_487 : _GEN_7326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7328 = 9'h1e8 == _GEN_12214 ? phv_data_488 : _GEN_7327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7329 = 9'h1e9 == _GEN_12214 ? phv_data_489 : _GEN_7328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7330 = 9'h1ea == _GEN_12214 ? phv_data_490 : _GEN_7329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7331 = 9'h1eb == _GEN_12214 ? phv_data_491 : _GEN_7330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7332 = 9'h1ec == _GEN_12214 ? phv_data_492 : _GEN_7331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7333 = 9'h1ed == _GEN_12214 ? phv_data_493 : _GEN_7332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7334 = 9'h1ee == _GEN_12214 ? phv_data_494 : _GEN_7333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7335 = 9'h1ef == _GEN_12214 ? phv_data_495 : _GEN_7334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7336 = 9'h1f0 == _GEN_12214 ? phv_data_496 : _GEN_7335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7337 = 9'h1f1 == _GEN_12214 ? phv_data_497 : _GEN_7336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7338 = 9'h1f2 == _GEN_12214 ? phv_data_498 : _GEN_7337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7339 = 9'h1f3 == _GEN_12214 ? phv_data_499 : _GEN_7338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7340 = 9'h1f4 == _GEN_12214 ? phv_data_500 : _GEN_7339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7341 = 9'h1f5 == _GEN_12214 ? phv_data_501 : _GEN_7340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7342 = 9'h1f6 == _GEN_12214 ? phv_data_502 : _GEN_7341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7343 = 9'h1f7 == _GEN_12214 ? phv_data_503 : _GEN_7342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7344 = 9'h1f8 == _GEN_12214 ? phv_data_504 : _GEN_7343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7345 = 9'h1f9 == _GEN_12214 ? phv_data_505 : _GEN_7344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7346 = 9'h1fa == _GEN_12214 ? phv_data_506 : _GEN_7345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7347 = 9'h1fb == _GEN_12214 ? phv_data_507 : _GEN_7346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7348 = 9'h1fc == _GEN_12214 ? phv_data_508 : _GEN_7347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7349 = 9'h1fd == _GEN_12214 ? phv_data_509 : _GEN_7348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7350 = 9'h1fe == _GEN_12214 ? phv_data_510 : _GEN_7349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_3 = 9'h1ff == _GEN_12214 ? phv_data_511 : _GEN_7350; // @[executor.scala 197:66 executor.scala 197:66]
  wire  _mask_3_T_24 = ending_3 == 2'h0; // @[executor.scala 199:88]
  wire  mask_3_3 = 2'h0 >= offset_3[1:0] & (2'h0 < ending_3 | ending_3 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_13 = {total_offset_hi_3,2'h1}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_7353 = 8'h1 == total_offset_13 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7354 = 8'h2 == total_offset_13 ? phv_data_2 : _GEN_7353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7355 = 8'h3 == total_offset_13 ? phv_data_3 : _GEN_7354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7356 = 8'h4 == total_offset_13 ? phv_data_4 : _GEN_7355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7357 = 8'h5 == total_offset_13 ? phv_data_5 : _GEN_7356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7358 = 8'h6 == total_offset_13 ? phv_data_6 : _GEN_7357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7359 = 8'h7 == total_offset_13 ? phv_data_7 : _GEN_7358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7360 = 8'h8 == total_offset_13 ? phv_data_8 : _GEN_7359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7361 = 8'h9 == total_offset_13 ? phv_data_9 : _GEN_7360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7362 = 8'ha == total_offset_13 ? phv_data_10 : _GEN_7361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7363 = 8'hb == total_offset_13 ? phv_data_11 : _GEN_7362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7364 = 8'hc == total_offset_13 ? phv_data_12 : _GEN_7363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7365 = 8'hd == total_offset_13 ? phv_data_13 : _GEN_7364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7366 = 8'he == total_offset_13 ? phv_data_14 : _GEN_7365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7367 = 8'hf == total_offset_13 ? phv_data_15 : _GEN_7366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7368 = 8'h10 == total_offset_13 ? phv_data_16 : _GEN_7367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7369 = 8'h11 == total_offset_13 ? phv_data_17 : _GEN_7368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7370 = 8'h12 == total_offset_13 ? phv_data_18 : _GEN_7369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7371 = 8'h13 == total_offset_13 ? phv_data_19 : _GEN_7370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7372 = 8'h14 == total_offset_13 ? phv_data_20 : _GEN_7371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7373 = 8'h15 == total_offset_13 ? phv_data_21 : _GEN_7372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7374 = 8'h16 == total_offset_13 ? phv_data_22 : _GEN_7373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7375 = 8'h17 == total_offset_13 ? phv_data_23 : _GEN_7374; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7376 = 8'h18 == total_offset_13 ? phv_data_24 : _GEN_7375; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7377 = 8'h19 == total_offset_13 ? phv_data_25 : _GEN_7376; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7378 = 8'h1a == total_offset_13 ? phv_data_26 : _GEN_7377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7379 = 8'h1b == total_offset_13 ? phv_data_27 : _GEN_7378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7380 = 8'h1c == total_offset_13 ? phv_data_28 : _GEN_7379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7381 = 8'h1d == total_offset_13 ? phv_data_29 : _GEN_7380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7382 = 8'h1e == total_offset_13 ? phv_data_30 : _GEN_7381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7383 = 8'h1f == total_offset_13 ? phv_data_31 : _GEN_7382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7384 = 8'h20 == total_offset_13 ? phv_data_32 : _GEN_7383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7385 = 8'h21 == total_offset_13 ? phv_data_33 : _GEN_7384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7386 = 8'h22 == total_offset_13 ? phv_data_34 : _GEN_7385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7387 = 8'h23 == total_offset_13 ? phv_data_35 : _GEN_7386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7388 = 8'h24 == total_offset_13 ? phv_data_36 : _GEN_7387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7389 = 8'h25 == total_offset_13 ? phv_data_37 : _GEN_7388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7390 = 8'h26 == total_offset_13 ? phv_data_38 : _GEN_7389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7391 = 8'h27 == total_offset_13 ? phv_data_39 : _GEN_7390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7392 = 8'h28 == total_offset_13 ? phv_data_40 : _GEN_7391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7393 = 8'h29 == total_offset_13 ? phv_data_41 : _GEN_7392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7394 = 8'h2a == total_offset_13 ? phv_data_42 : _GEN_7393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7395 = 8'h2b == total_offset_13 ? phv_data_43 : _GEN_7394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7396 = 8'h2c == total_offset_13 ? phv_data_44 : _GEN_7395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7397 = 8'h2d == total_offset_13 ? phv_data_45 : _GEN_7396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7398 = 8'h2e == total_offset_13 ? phv_data_46 : _GEN_7397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7399 = 8'h2f == total_offset_13 ? phv_data_47 : _GEN_7398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7400 = 8'h30 == total_offset_13 ? phv_data_48 : _GEN_7399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7401 = 8'h31 == total_offset_13 ? phv_data_49 : _GEN_7400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7402 = 8'h32 == total_offset_13 ? phv_data_50 : _GEN_7401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7403 = 8'h33 == total_offset_13 ? phv_data_51 : _GEN_7402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7404 = 8'h34 == total_offset_13 ? phv_data_52 : _GEN_7403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7405 = 8'h35 == total_offset_13 ? phv_data_53 : _GEN_7404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7406 = 8'h36 == total_offset_13 ? phv_data_54 : _GEN_7405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7407 = 8'h37 == total_offset_13 ? phv_data_55 : _GEN_7406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7408 = 8'h38 == total_offset_13 ? phv_data_56 : _GEN_7407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7409 = 8'h39 == total_offset_13 ? phv_data_57 : _GEN_7408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7410 = 8'h3a == total_offset_13 ? phv_data_58 : _GEN_7409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7411 = 8'h3b == total_offset_13 ? phv_data_59 : _GEN_7410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7412 = 8'h3c == total_offset_13 ? phv_data_60 : _GEN_7411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7413 = 8'h3d == total_offset_13 ? phv_data_61 : _GEN_7412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7414 = 8'h3e == total_offset_13 ? phv_data_62 : _GEN_7413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7415 = 8'h3f == total_offset_13 ? phv_data_63 : _GEN_7414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7416 = 8'h40 == total_offset_13 ? phv_data_64 : _GEN_7415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7417 = 8'h41 == total_offset_13 ? phv_data_65 : _GEN_7416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7418 = 8'h42 == total_offset_13 ? phv_data_66 : _GEN_7417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7419 = 8'h43 == total_offset_13 ? phv_data_67 : _GEN_7418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7420 = 8'h44 == total_offset_13 ? phv_data_68 : _GEN_7419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7421 = 8'h45 == total_offset_13 ? phv_data_69 : _GEN_7420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7422 = 8'h46 == total_offset_13 ? phv_data_70 : _GEN_7421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7423 = 8'h47 == total_offset_13 ? phv_data_71 : _GEN_7422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7424 = 8'h48 == total_offset_13 ? phv_data_72 : _GEN_7423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7425 = 8'h49 == total_offset_13 ? phv_data_73 : _GEN_7424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7426 = 8'h4a == total_offset_13 ? phv_data_74 : _GEN_7425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7427 = 8'h4b == total_offset_13 ? phv_data_75 : _GEN_7426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7428 = 8'h4c == total_offset_13 ? phv_data_76 : _GEN_7427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7429 = 8'h4d == total_offset_13 ? phv_data_77 : _GEN_7428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7430 = 8'h4e == total_offset_13 ? phv_data_78 : _GEN_7429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7431 = 8'h4f == total_offset_13 ? phv_data_79 : _GEN_7430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7432 = 8'h50 == total_offset_13 ? phv_data_80 : _GEN_7431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7433 = 8'h51 == total_offset_13 ? phv_data_81 : _GEN_7432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7434 = 8'h52 == total_offset_13 ? phv_data_82 : _GEN_7433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7435 = 8'h53 == total_offset_13 ? phv_data_83 : _GEN_7434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7436 = 8'h54 == total_offset_13 ? phv_data_84 : _GEN_7435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7437 = 8'h55 == total_offset_13 ? phv_data_85 : _GEN_7436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7438 = 8'h56 == total_offset_13 ? phv_data_86 : _GEN_7437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7439 = 8'h57 == total_offset_13 ? phv_data_87 : _GEN_7438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7440 = 8'h58 == total_offset_13 ? phv_data_88 : _GEN_7439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7441 = 8'h59 == total_offset_13 ? phv_data_89 : _GEN_7440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7442 = 8'h5a == total_offset_13 ? phv_data_90 : _GEN_7441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7443 = 8'h5b == total_offset_13 ? phv_data_91 : _GEN_7442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7444 = 8'h5c == total_offset_13 ? phv_data_92 : _GEN_7443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7445 = 8'h5d == total_offset_13 ? phv_data_93 : _GEN_7444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7446 = 8'h5e == total_offset_13 ? phv_data_94 : _GEN_7445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7447 = 8'h5f == total_offset_13 ? phv_data_95 : _GEN_7446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7448 = 8'h60 == total_offset_13 ? phv_data_96 : _GEN_7447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7449 = 8'h61 == total_offset_13 ? phv_data_97 : _GEN_7448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7450 = 8'h62 == total_offset_13 ? phv_data_98 : _GEN_7449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7451 = 8'h63 == total_offset_13 ? phv_data_99 : _GEN_7450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7452 = 8'h64 == total_offset_13 ? phv_data_100 : _GEN_7451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7453 = 8'h65 == total_offset_13 ? phv_data_101 : _GEN_7452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7454 = 8'h66 == total_offset_13 ? phv_data_102 : _GEN_7453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7455 = 8'h67 == total_offset_13 ? phv_data_103 : _GEN_7454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7456 = 8'h68 == total_offset_13 ? phv_data_104 : _GEN_7455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7457 = 8'h69 == total_offset_13 ? phv_data_105 : _GEN_7456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7458 = 8'h6a == total_offset_13 ? phv_data_106 : _GEN_7457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7459 = 8'h6b == total_offset_13 ? phv_data_107 : _GEN_7458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7460 = 8'h6c == total_offset_13 ? phv_data_108 : _GEN_7459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7461 = 8'h6d == total_offset_13 ? phv_data_109 : _GEN_7460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7462 = 8'h6e == total_offset_13 ? phv_data_110 : _GEN_7461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7463 = 8'h6f == total_offset_13 ? phv_data_111 : _GEN_7462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7464 = 8'h70 == total_offset_13 ? phv_data_112 : _GEN_7463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7465 = 8'h71 == total_offset_13 ? phv_data_113 : _GEN_7464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7466 = 8'h72 == total_offset_13 ? phv_data_114 : _GEN_7465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7467 = 8'h73 == total_offset_13 ? phv_data_115 : _GEN_7466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7468 = 8'h74 == total_offset_13 ? phv_data_116 : _GEN_7467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7469 = 8'h75 == total_offset_13 ? phv_data_117 : _GEN_7468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7470 = 8'h76 == total_offset_13 ? phv_data_118 : _GEN_7469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7471 = 8'h77 == total_offset_13 ? phv_data_119 : _GEN_7470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7472 = 8'h78 == total_offset_13 ? phv_data_120 : _GEN_7471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7473 = 8'h79 == total_offset_13 ? phv_data_121 : _GEN_7472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7474 = 8'h7a == total_offset_13 ? phv_data_122 : _GEN_7473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7475 = 8'h7b == total_offset_13 ? phv_data_123 : _GEN_7474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7476 = 8'h7c == total_offset_13 ? phv_data_124 : _GEN_7475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7477 = 8'h7d == total_offset_13 ? phv_data_125 : _GEN_7476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7478 = 8'h7e == total_offset_13 ? phv_data_126 : _GEN_7477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7479 = 8'h7f == total_offset_13 ? phv_data_127 : _GEN_7478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7480 = 8'h80 == total_offset_13 ? phv_data_128 : _GEN_7479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7481 = 8'h81 == total_offset_13 ? phv_data_129 : _GEN_7480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7482 = 8'h82 == total_offset_13 ? phv_data_130 : _GEN_7481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7483 = 8'h83 == total_offset_13 ? phv_data_131 : _GEN_7482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7484 = 8'h84 == total_offset_13 ? phv_data_132 : _GEN_7483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7485 = 8'h85 == total_offset_13 ? phv_data_133 : _GEN_7484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7486 = 8'h86 == total_offset_13 ? phv_data_134 : _GEN_7485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7487 = 8'h87 == total_offset_13 ? phv_data_135 : _GEN_7486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7488 = 8'h88 == total_offset_13 ? phv_data_136 : _GEN_7487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7489 = 8'h89 == total_offset_13 ? phv_data_137 : _GEN_7488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7490 = 8'h8a == total_offset_13 ? phv_data_138 : _GEN_7489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7491 = 8'h8b == total_offset_13 ? phv_data_139 : _GEN_7490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7492 = 8'h8c == total_offset_13 ? phv_data_140 : _GEN_7491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7493 = 8'h8d == total_offset_13 ? phv_data_141 : _GEN_7492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7494 = 8'h8e == total_offset_13 ? phv_data_142 : _GEN_7493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7495 = 8'h8f == total_offset_13 ? phv_data_143 : _GEN_7494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7496 = 8'h90 == total_offset_13 ? phv_data_144 : _GEN_7495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7497 = 8'h91 == total_offset_13 ? phv_data_145 : _GEN_7496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7498 = 8'h92 == total_offset_13 ? phv_data_146 : _GEN_7497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7499 = 8'h93 == total_offset_13 ? phv_data_147 : _GEN_7498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7500 = 8'h94 == total_offset_13 ? phv_data_148 : _GEN_7499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7501 = 8'h95 == total_offset_13 ? phv_data_149 : _GEN_7500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7502 = 8'h96 == total_offset_13 ? phv_data_150 : _GEN_7501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7503 = 8'h97 == total_offset_13 ? phv_data_151 : _GEN_7502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7504 = 8'h98 == total_offset_13 ? phv_data_152 : _GEN_7503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7505 = 8'h99 == total_offset_13 ? phv_data_153 : _GEN_7504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7506 = 8'h9a == total_offset_13 ? phv_data_154 : _GEN_7505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7507 = 8'h9b == total_offset_13 ? phv_data_155 : _GEN_7506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7508 = 8'h9c == total_offset_13 ? phv_data_156 : _GEN_7507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7509 = 8'h9d == total_offset_13 ? phv_data_157 : _GEN_7508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7510 = 8'h9e == total_offset_13 ? phv_data_158 : _GEN_7509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7511 = 8'h9f == total_offset_13 ? phv_data_159 : _GEN_7510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7512 = 8'ha0 == total_offset_13 ? phv_data_160 : _GEN_7511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7513 = 8'ha1 == total_offset_13 ? phv_data_161 : _GEN_7512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7514 = 8'ha2 == total_offset_13 ? phv_data_162 : _GEN_7513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7515 = 8'ha3 == total_offset_13 ? phv_data_163 : _GEN_7514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7516 = 8'ha4 == total_offset_13 ? phv_data_164 : _GEN_7515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7517 = 8'ha5 == total_offset_13 ? phv_data_165 : _GEN_7516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7518 = 8'ha6 == total_offset_13 ? phv_data_166 : _GEN_7517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7519 = 8'ha7 == total_offset_13 ? phv_data_167 : _GEN_7518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7520 = 8'ha8 == total_offset_13 ? phv_data_168 : _GEN_7519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7521 = 8'ha9 == total_offset_13 ? phv_data_169 : _GEN_7520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7522 = 8'haa == total_offset_13 ? phv_data_170 : _GEN_7521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7523 = 8'hab == total_offset_13 ? phv_data_171 : _GEN_7522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7524 = 8'hac == total_offset_13 ? phv_data_172 : _GEN_7523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7525 = 8'had == total_offset_13 ? phv_data_173 : _GEN_7524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7526 = 8'hae == total_offset_13 ? phv_data_174 : _GEN_7525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7527 = 8'haf == total_offset_13 ? phv_data_175 : _GEN_7526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7528 = 8'hb0 == total_offset_13 ? phv_data_176 : _GEN_7527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7529 = 8'hb1 == total_offset_13 ? phv_data_177 : _GEN_7528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7530 = 8'hb2 == total_offset_13 ? phv_data_178 : _GEN_7529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7531 = 8'hb3 == total_offset_13 ? phv_data_179 : _GEN_7530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7532 = 8'hb4 == total_offset_13 ? phv_data_180 : _GEN_7531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7533 = 8'hb5 == total_offset_13 ? phv_data_181 : _GEN_7532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7534 = 8'hb6 == total_offset_13 ? phv_data_182 : _GEN_7533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7535 = 8'hb7 == total_offset_13 ? phv_data_183 : _GEN_7534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7536 = 8'hb8 == total_offset_13 ? phv_data_184 : _GEN_7535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7537 = 8'hb9 == total_offset_13 ? phv_data_185 : _GEN_7536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7538 = 8'hba == total_offset_13 ? phv_data_186 : _GEN_7537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7539 = 8'hbb == total_offset_13 ? phv_data_187 : _GEN_7538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7540 = 8'hbc == total_offset_13 ? phv_data_188 : _GEN_7539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7541 = 8'hbd == total_offset_13 ? phv_data_189 : _GEN_7540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7542 = 8'hbe == total_offset_13 ? phv_data_190 : _GEN_7541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7543 = 8'hbf == total_offset_13 ? phv_data_191 : _GEN_7542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7544 = 8'hc0 == total_offset_13 ? phv_data_192 : _GEN_7543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7545 = 8'hc1 == total_offset_13 ? phv_data_193 : _GEN_7544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7546 = 8'hc2 == total_offset_13 ? phv_data_194 : _GEN_7545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7547 = 8'hc3 == total_offset_13 ? phv_data_195 : _GEN_7546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7548 = 8'hc4 == total_offset_13 ? phv_data_196 : _GEN_7547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7549 = 8'hc5 == total_offset_13 ? phv_data_197 : _GEN_7548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7550 = 8'hc6 == total_offset_13 ? phv_data_198 : _GEN_7549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7551 = 8'hc7 == total_offset_13 ? phv_data_199 : _GEN_7550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7552 = 8'hc8 == total_offset_13 ? phv_data_200 : _GEN_7551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7553 = 8'hc9 == total_offset_13 ? phv_data_201 : _GEN_7552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7554 = 8'hca == total_offset_13 ? phv_data_202 : _GEN_7553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7555 = 8'hcb == total_offset_13 ? phv_data_203 : _GEN_7554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7556 = 8'hcc == total_offset_13 ? phv_data_204 : _GEN_7555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7557 = 8'hcd == total_offset_13 ? phv_data_205 : _GEN_7556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7558 = 8'hce == total_offset_13 ? phv_data_206 : _GEN_7557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7559 = 8'hcf == total_offset_13 ? phv_data_207 : _GEN_7558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7560 = 8'hd0 == total_offset_13 ? phv_data_208 : _GEN_7559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7561 = 8'hd1 == total_offset_13 ? phv_data_209 : _GEN_7560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7562 = 8'hd2 == total_offset_13 ? phv_data_210 : _GEN_7561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7563 = 8'hd3 == total_offset_13 ? phv_data_211 : _GEN_7562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7564 = 8'hd4 == total_offset_13 ? phv_data_212 : _GEN_7563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7565 = 8'hd5 == total_offset_13 ? phv_data_213 : _GEN_7564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7566 = 8'hd6 == total_offset_13 ? phv_data_214 : _GEN_7565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7567 = 8'hd7 == total_offset_13 ? phv_data_215 : _GEN_7566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7568 = 8'hd8 == total_offset_13 ? phv_data_216 : _GEN_7567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7569 = 8'hd9 == total_offset_13 ? phv_data_217 : _GEN_7568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7570 = 8'hda == total_offset_13 ? phv_data_218 : _GEN_7569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7571 = 8'hdb == total_offset_13 ? phv_data_219 : _GEN_7570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7572 = 8'hdc == total_offset_13 ? phv_data_220 : _GEN_7571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7573 = 8'hdd == total_offset_13 ? phv_data_221 : _GEN_7572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7574 = 8'hde == total_offset_13 ? phv_data_222 : _GEN_7573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7575 = 8'hdf == total_offset_13 ? phv_data_223 : _GEN_7574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7576 = 8'he0 == total_offset_13 ? phv_data_224 : _GEN_7575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7577 = 8'he1 == total_offset_13 ? phv_data_225 : _GEN_7576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7578 = 8'he2 == total_offset_13 ? phv_data_226 : _GEN_7577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7579 = 8'he3 == total_offset_13 ? phv_data_227 : _GEN_7578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7580 = 8'he4 == total_offset_13 ? phv_data_228 : _GEN_7579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7581 = 8'he5 == total_offset_13 ? phv_data_229 : _GEN_7580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7582 = 8'he6 == total_offset_13 ? phv_data_230 : _GEN_7581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7583 = 8'he7 == total_offset_13 ? phv_data_231 : _GEN_7582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7584 = 8'he8 == total_offset_13 ? phv_data_232 : _GEN_7583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7585 = 8'he9 == total_offset_13 ? phv_data_233 : _GEN_7584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7586 = 8'hea == total_offset_13 ? phv_data_234 : _GEN_7585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7587 = 8'heb == total_offset_13 ? phv_data_235 : _GEN_7586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7588 = 8'hec == total_offset_13 ? phv_data_236 : _GEN_7587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7589 = 8'hed == total_offset_13 ? phv_data_237 : _GEN_7588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7590 = 8'hee == total_offset_13 ? phv_data_238 : _GEN_7589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7591 = 8'hef == total_offset_13 ? phv_data_239 : _GEN_7590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7592 = 8'hf0 == total_offset_13 ? phv_data_240 : _GEN_7591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7593 = 8'hf1 == total_offset_13 ? phv_data_241 : _GEN_7592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7594 = 8'hf2 == total_offset_13 ? phv_data_242 : _GEN_7593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7595 = 8'hf3 == total_offset_13 ? phv_data_243 : _GEN_7594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7596 = 8'hf4 == total_offset_13 ? phv_data_244 : _GEN_7595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7597 = 8'hf5 == total_offset_13 ? phv_data_245 : _GEN_7596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7598 = 8'hf6 == total_offset_13 ? phv_data_246 : _GEN_7597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7599 = 8'hf7 == total_offset_13 ? phv_data_247 : _GEN_7598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7600 = 8'hf8 == total_offset_13 ? phv_data_248 : _GEN_7599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7601 = 8'hf9 == total_offset_13 ? phv_data_249 : _GEN_7600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7602 = 8'hfa == total_offset_13 ? phv_data_250 : _GEN_7601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7603 = 8'hfb == total_offset_13 ? phv_data_251 : _GEN_7602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7604 = 8'hfc == total_offset_13 ? phv_data_252 : _GEN_7603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7605 = 8'hfd == total_offset_13 ? phv_data_253 : _GEN_7604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7606 = 8'hfe == total_offset_13 ? phv_data_254 : _GEN_7605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7607 = 8'hff == total_offset_13 ? phv_data_255 : _GEN_7606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_12470 = {{1'd0}, total_offset_13}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7608 = 9'h100 == _GEN_12470 ? phv_data_256 : _GEN_7607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7609 = 9'h101 == _GEN_12470 ? phv_data_257 : _GEN_7608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7610 = 9'h102 == _GEN_12470 ? phv_data_258 : _GEN_7609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7611 = 9'h103 == _GEN_12470 ? phv_data_259 : _GEN_7610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7612 = 9'h104 == _GEN_12470 ? phv_data_260 : _GEN_7611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7613 = 9'h105 == _GEN_12470 ? phv_data_261 : _GEN_7612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7614 = 9'h106 == _GEN_12470 ? phv_data_262 : _GEN_7613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7615 = 9'h107 == _GEN_12470 ? phv_data_263 : _GEN_7614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7616 = 9'h108 == _GEN_12470 ? phv_data_264 : _GEN_7615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7617 = 9'h109 == _GEN_12470 ? phv_data_265 : _GEN_7616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7618 = 9'h10a == _GEN_12470 ? phv_data_266 : _GEN_7617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7619 = 9'h10b == _GEN_12470 ? phv_data_267 : _GEN_7618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7620 = 9'h10c == _GEN_12470 ? phv_data_268 : _GEN_7619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7621 = 9'h10d == _GEN_12470 ? phv_data_269 : _GEN_7620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7622 = 9'h10e == _GEN_12470 ? phv_data_270 : _GEN_7621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7623 = 9'h10f == _GEN_12470 ? phv_data_271 : _GEN_7622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7624 = 9'h110 == _GEN_12470 ? phv_data_272 : _GEN_7623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7625 = 9'h111 == _GEN_12470 ? phv_data_273 : _GEN_7624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7626 = 9'h112 == _GEN_12470 ? phv_data_274 : _GEN_7625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7627 = 9'h113 == _GEN_12470 ? phv_data_275 : _GEN_7626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7628 = 9'h114 == _GEN_12470 ? phv_data_276 : _GEN_7627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7629 = 9'h115 == _GEN_12470 ? phv_data_277 : _GEN_7628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7630 = 9'h116 == _GEN_12470 ? phv_data_278 : _GEN_7629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7631 = 9'h117 == _GEN_12470 ? phv_data_279 : _GEN_7630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7632 = 9'h118 == _GEN_12470 ? phv_data_280 : _GEN_7631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7633 = 9'h119 == _GEN_12470 ? phv_data_281 : _GEN_7632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7634 = 9'h11a == _GEN_12470 ? phv_data_282 : _GEN_7633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7635 = 9'h11b == _GEN_12470 ? phv_data_283 : _GEN_7634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7636 = 9'h11c == _GEN_12470 ? phv_data_284 : _GEN_7635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7637 = 9'h11d == _GEN_12470 ? phv_data_285 : _GEN_7636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7638 = 9'h11e == _GEN_12470 ? phv_data_286 : _GEN_7637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7639 = 9'h11f == _GEN_12470 ? phv_data_287 : _GEN_7638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7640 = 9'h120 == _GEN_12470 ? phv_data_288 : _GEN_7639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7641 = 9'h121 == _GEN_12470 ? phv_data_289 : _GEN_7640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7642 = 9'h122 == _GEN_12470 ? phv_data_290 : _GEN_7641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7643 = 9'h123 == _GEN_12470 ? phv_data_291 : _GEN_7642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7644 = 9'h124 == _GEN_12470 ? phv_data_292 : _GEN_7643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7645 = 9'h125 == _GEN_12470 ? phv_data_293 : _GEN_7644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7646 = 9'h126 == _GEN_12470 ? phv_data_294 : _GEN_7645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7647 = 9'h127 == _GEN_12470 ? phv_data_295 : _GEN_7646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7648 = 9'h128 == _GEN_12470 ? phv_data_296 : _GEN_7647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7649 = 9'h129 == _GEN_12470 ? phv_data_297 : _GEN_7648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7650 = 9'h12a == _GEN_12470 ? phv_data_298 : _GEN_7649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7651 = 9'h12b == _GEN_12470 ? phv_data_299 : _GEN_7650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7652 = 9'h12c == _GEN_12470 ? phv_data_300 : _GEN_7651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7653 = 9'h12d == _GEN_12470 ? phv_data_301 : _GEN_7652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7654 = 9'h12e == _GEN_12470 ? phv_data_302 : _GEN_7653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7655 = 9'h12f == _GEN_12470 ? phv_data_303 : _GEN_7654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7656 = 9'h130 == _GEN_12470 ? phv_data_304 : _GEN_7655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7657 = 9'h131 == _GEN_12470 ? phv_data_305 : _GEN_7656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7658 = 9'h132 == _GEN_12470 ? phv_data_306 : _GEN_7657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7659 = 9'h133 == _GEN_12470 ? phv_data_307 : _GEN_7658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7660 = 9'h134 == _GEN_12470 ? phv_data_308 : _GEN_7659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7661 = 9'h135 == _GEN_12470 ? phv_data_309 : _GEN_7660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7662 = 9'h136 == _GEN_12470 ? phv_data_310 : _GEN_7661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7663 = 9'h137 == _GEN_12470 ? phv_data_311 : _GEN_7662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7664 = 9'h138 == _GEN_12470 ? phv_data_312 : _GEN_7663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7665 = 9'h139 == _GEN_12470 ? phv_data_313 : _GEN_7664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7666 = 9'h13a == _GEN_12470 ? phv_data_314 : _GEN_7665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7667 = 9'h13b == _GEN_12470 ? phv_data_315 : _GEN_7666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7668 = 9'h13c == _GEN_12470 ? phv_data_316 : _GEN_7667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7669 = 9'h13d == _GEN_12470 ? phv_data_317 : _GEN_7668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7670 = 9'h13e == _GEN_12470 ? phv_data_318 : _GEN_7669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7671 = 9'h13f == _GEN_12470 ? phv_data_319 : _GEN_7670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7672 = 9'h140 == _GEN_12470 ? phv_data_320 : _GEN_7671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7673 = 9'h141 == _GEN_12470 ? phv_data_321 : _GEN_7672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7674 = 9'h142 == _GEN_12470 ? phv_data_322 : _GEN_7673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7675 = 9'h143 == _GEN_12470 ? phv_data_323 : _GEN_7674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7676 = 9'h144 == _GEN_12470 ? phv_data_324 : _GEN_7675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7677 = 9'h145 == _GEN_12470 ? phv_data_325 : _GEN_7676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7678 = 9'h146 == _GEN_12470 ? phv_data_326 : _GEN_7677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7679 = 9'h147 == _GEN_12470 ? phv_data_327 : _GEN_7678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7680 = 9'h148 == _GEN_12470 ? phv_data_328 : _GEN_7679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7681 = 9'h149 == _GEN_12470 ? phv_data_329 : _GEN_7680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7682 = 9'h14a == _GEN_12470 ? phv_data_330 : _GEN_7681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7683 = 9'h14b == _GEN_12470 ? phv_data_331 : _GEN_7682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7684 = 9'h14c == _GEN_12470 ? phv_data_332 : _GEN_7683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7685 = 9'h14d == _GEN_12470 ? phv_data_333 : _GEN_7684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7686 = 9'h14e == _GEN_12470 ? phv_data_334 : _GEN_7685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7687 = 9'h14f == _GEN_12470 ? phv_data_335 : _GEN_7686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7688 = 9'h150 == _GEN_12470 ? phv_data_336 : _GEN_7687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7689 = 9'h151 == _GEN_12470 ? phv_data_337 : _GEN_7688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7690 = 9'h152 == _GEN_12470 ? phv_data_338 : _GEN_7689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7691 = 9'h153 == _GEN_12470 ? phv_data_339 : _GEN_7690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7692 = 9'h154 == _GEN_12470 ? phv_data_340 : _GEN_7691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7693 = 9'h155 == _GEN_12470 ? phv_data_341 : _GEN_7692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7694 = 9'h156 == _GEN_12470 ? phv_data_342 : _GEN_7693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7695 = 9'h157 == _GEN_12470 ? phv_data_343 : _GEN_7694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7696 = 9'h158 == _GEN_12470 ? phv_data_344 : _GEN_7695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7697 = 9'h159 == _GEN_12470 ? phv_data_345 : _GEN_7696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7698 = 9'h15a == _GEN_12470 ? phv_data_346 : _GEN_7697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7699 = 9'h15b == _GEN_12470 ? phv_data_347 : _GEN_7698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7700 = 9'h15c == _GEN_12470 ? phv_data_348 : _GEN_7699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7701 = 9'h15d == _GEN_12470 ? phv_data_349 : _GEN_7700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7702 = 9'h15e == _GEN_12470 ? phv_data_350 : _GEN_7701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7703 = 9'h15f == _GEN_12470 ? phv_data_351 : _GEN_7702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7704 = 9'h160 == _GEN_12470 ? phv_data_352 : _GEN_7703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7705 = 9'h161 == _GEN_12470 ? phv_data_353 : _GEN_7704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7706 = 9'h162 == _GEN_12470 ? phv_data_354 : _GEN_7705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7707 = 9'h163 == _GEN_12470 ? phv_data_355 : _GEN_7706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7708 = 9'h164 == _GEN_12470 ? phv_data_356 : _GEN_7707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7709 = 9'h165 == _GEN_12470 ? phv_data_357 : _GEN_7708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7710 = 9'h166 == _GEN_12470 ? phv_data_358 : _GEN_7709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7711 = 9'h167 == _GEN_12470 ? phv_data_359 : _GEN_7710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7712 = 9'h168 == _GEN_12470 ? phv_data_360 : _GEN_7711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7713 = 9'h169 == _GEN_12470 ? phv_data_361 : _GEN_7712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7714 = 9'h16a == _GEN_12470 ? phv_data_362 : _GEN_7713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7715 = 9'h16b == _GEN_12470 ? phv_data_363 : _GEN_7714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7716 = 9'h16c == _GEN_12470 ? phv_data_364 : _GEN_7715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7717 = 9'h16d == _GEN_12470 ? phv_data_365 : _GEN_7716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7718 = 9'h16e == _GEN_12470 ? phv_data_366 : _GEN_7717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7719 = 9'h16f == _GEN_12470 ? phv_data_367 : _GEN_7718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7720 = 9'h170 == _GEN_12470 ? phv_data_368 : _GEN_7719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7721 = 9'h171 == _GEN_12470 ? phv_data_369 : _GEN_7720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7722 = 9'h172 == _GEN_12470 ? phv_data_370 : _GEN_7721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7723 = 9'h173 == _GEN_12470 ? phv_data_371 : _GEN_7722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7724 = 9'h174 == _GEN_12470 ? phv_data_372 : _GEN_7723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7725 = 9'h175 == _GEN_12470 ? phv_data_373 : _GEN_7724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7726 = 9'h176 == _GEN_12470 ? phv_data_374 : _GEN_7725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7727 = 9'h177 == _GEN_12470 ? phv_data_375 : _GEN_7726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7728 = 9'h178 == _GEN_12470 ? phv_data_376 : _GEN_7727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7729 = 9'h179 == _GEN_12470 ? phv_data_377 : _GEN_7728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7730 = 9'h17a == _GEN_12470 ? phv_data_378 : _GEN_7729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7731 = 9'h17b == _GEN_12470 ? phv_data_379 : _GEN_7730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7732 = 9'h17c == _GEN_12470 ? phv_data_380 : _GEN_7731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7733 = 9'h17d == _GEN_12470 ? phv_data_381 : _GEN_7732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7734 = 9'h17e == _GEN_12470 ? phv_data_382 : _GEN_7733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7735 = 9'h17f == _GEN_12470 ? phv_data_383 : _GEN_7734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7736 = 9'h180 == _GEN_12470 ? phv_data_384 : _GEN_7735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7737 = 9'h181 == _GEN_12470 ? phv_data_385 : _GEN_7736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7738 = 9'h182 == _GEN_12470 ? phv_data_386 : _GEN_7737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7739 = 9'h183 == _GEN_12470 ? phv_data_387 : _GEN_7738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7740 = 9'h184 == _GEN_12470 ? phv_data_388 : _GEN_7739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7741 = 9'h185 == _GEN_12470 ? phv_data_389 : _GEN_7740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7742 = 9'h186 == _GEN_12470 ? phv_data_390 : _GEN_7741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7743 = 9'h187 == _GEN_12470 ? phv_data_391 : _GEN_7742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7744 = 9'h188 == _GEN_12470 ? phv_data_392 : _GEN_7743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7745 = 9'h189 == _GEN_12470 ? phv_data_393 : _GEN_7744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7746 = 9'h18a == _GEN_12470 ? phv_data_394 : _GEN_7745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7747 = 9'h18b == _GEN_12470 ? phv_data_395 : _GEN_7746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7748 = 9'h18c == _GEN_12470 ? phv_data_396 : _GEN_7747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7749 = 9'h18d == _GEN_12470 ? phv_data_397 : _GEN_7748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7750 = 9'h18e == _GEN_12470 ? phv_data_398 : _GEN_7749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7751 = 9'h18f == _GEN_12470 ? phv_data_399 : _GEN_7750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7752 = 9'h190 == _GEN_12470 ? phv_data_400 : _GEN_7751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7753 = 9'h191 == _GEN_12470 ? phv_data_401 : _GEN_7752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7754 = 9'h192 == _GEN_12470 ? phv_data_402 : _GEN_7753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7755 = 9'h193 == _GEN_12470 ? phv_data_403 : _GEN_7754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7756 = 9'h194 == _GEN_12470 ? phv_data_404 : _GEN_7755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7757 = 9'h195 == _GEN_12470 ? phv_data_405 : _GEN_7756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7758 = 9'h196 == _GEN_12470 ? phv_data_406 : _GEN_7757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7759 = 9'h197 == _GEN_12470 ? phv_data_407 : _GEN_7758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7760 = 9'h198 == _GEN_12470 ? phv_data_408 : _GEN_7759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7761 = 9'h199 == _GEN_12470 ? phv_data_409 : _GEN_7760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7762 = 9'h19a == _GEN_12470 ? phv_data_410 : _GEN_7761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7763 = 9'h19b == _GEN_12470 ? phv_data_411 : _GEN_7762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7764 = 9'h19c == _GEN_12470 ? phv_data_412 : _GEN_7763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7765 = 9'h19d == _GEN_12470 ? phv_data_413 : _GEN_7764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7766 = 9'h19e == _GEN_12470 ? phv_data_414 : _GEN_7765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7767 = 9'h19f == _GEN_12470 ? phv_data_415 : _GEN_7766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7768 = 9'h1a0 == _GEN_12470 ? phv_data_416 : _GEN_7767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7769 = 9'h1a1 == _GEN_12470 ? phv_data_417 : _GEN_7768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7770 = 9'h1a2 == _GEN_12470 ? phv_data_418 : _GEN_7769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7771 = 9'h1a3 == _GEN_12470 ? phv_data_419 : _GEN_7770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7772 = 9'h1a4 == _GEN_12470 ? phv_data_420 : _GEN_7771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7773 = 9'h1a5 == _GEN_12470 ? phv_data_421 : _GEN_7772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7774 = 9'h1a6 == _GEN_12470 ? phv_data_422 : _GEN_7773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7775 = 9'h1a7 == _GEN_12470 ? phv_data_423 : _GEN_7774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7776 = 9'h1a8 == _GEN_12470 ? phv_data_424 : _GEN_7775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7777 = 9'h1a9 == _GEN_12470 ? phv_data_425 : _GEN_7776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7778 = 9'h1aa == _GEN_12470 ? phv_data_426 : _GEN_7777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7779 = 9'h1ab == _GEN_12470 ? phv_data_427 : _GEN_7778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7780 = 9'h1ac == _GEN_12470 ? phv_data_428 : _GEN_7779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7781 = 9'h1ad == _GEN_12470 ? phv_data_429 : _GEN_7780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7782 = 9'h1ae == _GEN_12470 ? phv_data_430 : _GEN_7781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7783 = 9'h1af == _GEN_12470 ? phv_data_431 : _GEN_7782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7784 = 9'h1b0 == _GEN_12470 ? phv_data_432 : _GEN_7783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7785 = 9'h1b1 == _GEN_12470 ? phv_data_433 : _GEN_7784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7786 = 9'h1b2 == _GEN_12470 ? phv_data_434 : _GEN_7785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7787 = 9'h1b3 == _GEN_12470 ? phv_data_435 : _GEN_7786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7788 = 9'h1b4 == _GEN_12470 ? phv_data_436 : _GEN_7787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7789 = 9'h1b5 == _GEN_12470 ? phv_data_437 : _GEN_7788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7790 = 9'h1b6 == _GEN_12470 ? phv_data_438 : _GEN_7789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7791 = 9'h1b7 == _GEN_12470 ? phv_data_439 : _GEN_7790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7792 = 9'h1b8 == _GEN_12470 ? phv_data_440 : _GEN_7791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7793 = 9'h1b9 == _GEN_12470 ? phv_data_441 : _GEN_7792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7794 = 9'h1ba == _GEN_12470 ? phv_data_442 : _GEN_7793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7795 = 9'h1bb == _GEN_12470 ? phv_data_443 : _GEN_7794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7796 = 9'h1bc == _GEN_12470 ? phv_data_444 : _GEN_7795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7797 = 9'h1bd == _GEN_12470 ? phv_data_445 : _GEN_7796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7798 = 9'h1be == _GEN_12470 ? phv_data_446 : _GEN_7797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7799 = 9'h1bf == _GEN_12470 ? phv_data_447 : _GEN_7798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7800 = 9'h1c0 == _GEN_12470 ? phv_data_448 : _GEN_7799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7801 = 9'h1c1 == _GEN_12470 ? phv_data_449 : _GEN_7800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7802 = 9'h1c2 == _GEN_12470 ? phv_data_450 : _GEN_7801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7803 = 9'h1c3 == _GEN_12470 ? phv_data_451 : _GEN_7802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7804 = 9'h1c4 == _GEN_12470 ? phv_data_452 : _GEN_7803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7805 = 9'h1c5 == _GEN_12470 ? phv_data_453 : _GEN_7804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7806 = 9'h1c6 == _GEN_12470 ? phv_data_454 : _GEN_7805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7807 = 9'h1c7 == _GEN_12470 ? phv_data_455 : _GEN_7806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7808 = 9'h1c8 == _GEN_12470 ? phv_data_456 : _GEN_7807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7809 = 9'h1c9 == _GEN_12470 ? phv_data_457 : _GEN_7808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7810 = 9'h1ca == _GEN_12470 ? phv_data_458 : _GEN_7809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7811 = 9'h1cb == _GEN_12470 ? phv_data_459 : _GEN_7810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7812 = 9'h1cc == _GEN_12470 ? phv_data_460 : _GEN_7811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7813 = 9'h1cd == _GEN_12470 ? phv_data_461 : _GEN_7812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7814 = 9'h1ce == _GEN_12470 ? phv_data_462 : _GEN_7813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7815 = 9'h1cf == _GEN_12470 ? phv_data_463 : _GEN_7814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7816 = 9'h1d0 == _GEN_12470 ? phv_data_464 : _GEN_7815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7817 = 9'h1d1 == _GEN_12470 ? phv_data_465 : _GEN_7816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7818 = 9'h1d2 == _GEN_12470 ? phv_data_466 : _GEN_7817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7819 = 9'h1d3 == _GEN_12470 ? phv_data_467 : _GEN_7818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7820 = 9'h1d4 == _GEN_12470 ? phv_data_468 : _GEN_7819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7821 = 9'h1d5 == _GEN_12470 ? phv_data_469 : _GEN_7820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7822 = 9'h1d6 == _GEN_12470 ? phv_data_470 : _GEN_7821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7823 = 9'h1d7 == _GEN_12470 ? phv_data_471 : _GEN_7822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7824 = 9'h1d8 == _GEN_12470 ? phv_data_472 : _GEN_7823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7825 = 9'h1d9 == _GEN_12470 ? phv_data_473 : _GEN_7824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7826 = 9'h1da == _GEN_12470 ? phv_data_474 : _GEN_7825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7827 = 9'h1db == _GEN_12470 ? phv_data_475 : _GEN_7826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7828 = 9'h1dc == _GEN_12470 ? phv_data_476 : _GEN_7827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7829 = 9'h1dd == _GEN_12470 ? phv_data_477 : _GEN_7828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7830 = 9'h1de == _GEN_12470 ? phv_data_478 : _GEN_7829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7831 = 9'h1df == _GEN_12470 ? phv_data_479 : _GEN_7830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7832 = 9'h1e0 == _GEN_12470 ? phv_data_480 : _GEN_7831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7833 = 9'h1e1 == _GEN_12470 ? phv_data_481 : _GEN_7832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7834 = 9'h1e2 == _GEN_12470 ? phv_data_482 : _GEN_7833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7835 = 9'h1e3 == _GEN_12470 ? phv_data_483 : _GEN_7834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7836 = 9'h1e4 == _GEN_12470 ? phv_data_484 : _GEN_7835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7837 = 9'h1e5 == _GEN_12470 ? phv_data_485 : _GEN_7836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7838 = 9'h1e6 == _GEN_12470 ? phv_data_486 : _GEN_7837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7839 = 9'h1e7 == _GEN_12470 ? phv_data_487 : _GEN_7838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7840 = 9'h1e8 == _GEN_12470 ? phv_data_488 : _GEN_7839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7841 = 9'h1e9 == _GEN_12470 ? phv_data_489 : _GEN_7840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7842 = 9'h1ea == _GEN_12470 ? phv_data_490 : _GEN_7841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7843 = 9'h1eb == _GEN_12470 ? phv_data_491 : _GEN_7842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7844 = 9'h1ec == _GEN_12470 ? phv_data_492 : _GEN_7843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7845 = 9'h1ed == _GEN_12470 ? phv_data_493 : _GEN_7844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7846 = 9'h1ee == _GEN_12470 ? phv_data_494 : _GEN_7845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7847 = 9'h1ef == _GEN_12470 ? phv_data_495 : _GEN_7846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7848 = 9'h1f0 == _GEN_12470 ? phv_data_496 : _GEN_7847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7849 = 9'h1f1 == _GEN_12470 ? phv_data_497 : _GEN_7848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7850 = 9'h1f2 == _GEN_12470 ? phv_data_498 : _GEN_7849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7851 = 9'h1f3 == _GEN_12470 ? phv_data_499 : _GEN_7850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7852 = 9'h1f4 == _GEN_12470 ? phv_data_500 : _GEN_7851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7853 = 9'h1f5 == _GEN_12470 ? phv_data_501 : _GEN_7852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7854 = 9'h1f6 == _GEN_12470 ? phv_data_502 : _GEN_7853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7855 = 9'h1f7 == _GEN_12470 ? phv_data_503 : _GEN_7854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7856 = 9'h1f8 == _GEN_12470 ? phv_data_504 : _GEN_7855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7857 = 9'h1f9 == _GEN_12470 ? phv_data_505 : _GEN_7856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7858 = 9'h1fa == _GEN_12470 ? phv_data_506 : _GEN_7857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7859 = 9'h1fb == _GEN_12470 ? phv_data_507 : _GEN_7858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7860 = 9'h1fc == _GEN_12470 ? phv_data_508 : _GEN_7859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7861 = 9'h1fd == _GEN_12470 ? phv_data_509 : _GEN_7860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7862 = 9'h1fe == _GEN_12470 ? phv_data_510 : _GEN_7861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_2 = 9'h1ff == _GEN_12470 ? phv_data_511 : _GEN_7862; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_3_2 = 2'h1 >= offset_3[1:0] & (2'h1 < ending_3 | ending_3 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_14 = {total_offset_hi_3,2'h2}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_7865 = 8'h1 == total_offset_14 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7866 = 8'h2 == total_offset_14 ? phv_data_2 : _GEN_7865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7867 = 8'h3 == total_offset_14 ? phv_data_3 : _GEN_7866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7868 = 8'h4 == total_offset_14 ? phv_data_4 : _GEN_7867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7869 = 8'h5 == total_offset_14 ? phv_data_5 : _GEN_7868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7870 = 8'h6 == total_offset_14 ? phv_data_6 : _GEN_7869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7871 = 8'h7 == total_offset_14 ? phv_data_7 : _GEN_7870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7872 = 8'h8 == total_offset_14 ? phv_data_8 : _GEN_7871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7873 = 8'h9 == total_offset_14 ? phv_data_9 : _GEN_7872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7874 = 8'ha == total_offset_14 ? phv_data_10 : _GEN_7873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7875 = 8'hb == total_offset_14 ? phv_data_11 : _GEN_7874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7876 = 8'hc == total_offset_14 ? phv_data_12 : _GEN_7875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7877 = 8'hd == total_offset_14 ? phv_data_13 : _GEN_7876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7878 = 8'he == total_offset_14 ? phv_data_14 : _GEN_7877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7879 = 8'hf == total_offset_14 ? phv_data_15 : _GEN_7878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7880 = 8'h10 == total_offset_14 ? phv_data_16 : _GEN_7879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7881 = 8'h11 == total_offset_14 ? phv_data_17 : _GEN_7880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7882 = 8'h12 == total_offset_14 ? phv_data_18 : _GEN_7881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7883 = 8'h13 == total_offset_14 ? phv_data_19 : _GEN_7882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7884 = 8'h14 == total_offset_14 ? phv_data_20 : _GEN_7883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7885 = 8'h15 == total_offset_14 ? phv_data_21 : _GEN_7884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7886 = 8'h16 == total_offset_14 ? phv_data_22 : _GEN_7885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7887 = 8'h17 == total_offset_14 ? phv_data_23 : _GEN_7886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7888 = 8'h18 == total_offset_14 ? phv_data_24 : _GEN_7887; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7889 = 8'h19 == total_offset_14 ? phv_data_25 : _GEN_7888; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7890 = 8'h1a == total_offset_14 ? phv_data_26 : _GEN_7889; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7891 = 8'h1b == total_offset_14 ? phv_data_27 : _GEN_7890; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7892 = 8'h1c == total_offset_14 ? phv_data_28 : _GEN_7891; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7893 = 8'h1d == total_offset_14 ? phv_data_29 : _GEN_7892; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7894 = 8'h1e == total_offset_14 ? phv_data_30 : _GEN_7893; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7895 = 8'h1f == total_offset_14 ? phv_data_31 : _GEN_7894; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7896 = 8'h20 == total_offset_14 ? phv_data_32 : _GEN_7895; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7897 = 8'h21 == total_offset_14 ? phv_data_33 : _GEN_7896; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7898 = 8'h22 == total_offset_14 ? phv_data_34 : _GEN_7897; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7899 = 8'h23 == total_offset_14 ? phv_data_35 : _GEN_7898; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7900 = 8'h24 == total_offset_14 ? phv_data_36 : _GEN_7899; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7901 = 8'h25 == total_offset_14 ? phv_data_37 : _GEN_7900; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7902 = 8'h26 == total_offset_14 ? phv_data_38 : _GEN_7901; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7903 = 8'h27 == total_offset_14 ? phv_data_39 : _GEN_7902; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7904 = 8'h28 == total_offset_14 ? phv_data_40 : _GEN_7903; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7905 = 8'h29 == total_offset_14 ? phv_data_41 : _GEN_7904; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7906 = 8'h2a == total_offset_14 ? phv_data_42 : _GEN_7905; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7907 = 8'h2b == total_offset_14 ? phv_data_43 : _GEN_7906; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7908 = 8'h2c == total_offset_14 ? phv_data_44 : _GEN_7907; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7909 = 8'h2d == total_offset_14 ? phv_data_45 : _GEN_7908; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7910 = 8'h2e == total_offset_14 ? phv_data_46 : _GEN_7909; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7911 = 8'h2f == total_offset_14 ? phv_data_47 : _GEN_7910; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7912 = 8'h30 == total_offset_14 ? phv_data_48 : _GEN_7911; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7913 = 8'h31 == total_offset_14 ? phv_data_49 : _GEN_7912; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7914 = 8'h32 == total_offset_14 ? phv_data_50 : _GEN_7913; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7915 = 8'h33 == total_offset_14 ? phv_data_51 : _GEN_7914; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7916 = 8'h34 == total_offset_14 ? phv_data_52 : _GEN_7915; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7917 = 8'h35 == total_offset_14 ? phv_data_53 : _GEN_7916; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7918 = 8'h36 == total_offset_14 ? phv_data_54 : _GEN_7917; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7919 = 8'h37 == total_offset_14 ? phv_data_55 : _GEN_7918; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7920 = 8'h38 == total_offset_14 ? phv_data_56 : _GEN_7919; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7921 = 8'h39 == total_offset_14 ? phv_data_57 : _GEN_7920; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7922 = 8'h3a == total_offset_14 ? phv_data_58 : _GEN_7921; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7923 = 8'h3b == total_offset_14 ? phv_data_59 : _GEN_7922; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7924 = 8'h3c == total_offset_14 ? phv_data_60 : _GEN_7923; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7925 = 8'h3d == total_offset_14 ? phv_data_61 : _GEN_7924; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7926 = 8'h3e == total_offset_14 ? phv_data_62 : _GEN_7925; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7927 = 8'h3f == total_offset_14 ? phv_data_63 : _GEN_7926; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7928 = 8'h40 == total_offset_14 ? phv_data_64 : _GEN_7927; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7929 = 8'h41 == total_offset_14 ? phv_data_65 : _GEN_7928; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7930 = 8'h42 == total_offset_14 ? phv_data_66 : _GEN_7929; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7931 = 8'h43 == total_offset_14 ? phv_data_67 : _GEN_7930; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7932 = 8'h44 == total_offset_14 ? phv_data_68 : _GEN_7931; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7933 = 8'h45 == total_offset_14 ? phv_data_69 : _GEN_7932; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7934 = 8'h46 == total_offset_14 ? phv_data_70 : _GEN_7933; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7935 = 8'h47 == total_offset_14 ? phv_data_71 : _GEN_7934; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7936 = 8'h48 == total_offset_14 ? phv_data_72 : _GEN_7935; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7937 = 8'h49 == total_offset_14 ? phv_data_73 : _GEN_7936; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7938 = 8'h4a == total_offset_14 ? phv_data_74 : _GEN_7937; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7939 = 8'h4b == total_offset_14 ? phv_data_75 : _GEN_7938; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7940 = 8'h4c == total_offset_14 ? phv_data_76 : _GEN_7939; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7941 = 8'h4d == total_offset_14 ? phv_data_77 : _GEN_7940; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7942 = 8'h4e == total_offset_14 ? phv_data_78 : _GEN_7941; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7943 = 8'h4f == total_offset_14 ? phv_data_79 : _GEN_7942; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7944 = 8'h50 == total_offset_14 ? phv_data_80 : _GEN_7943; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7945 = 8'h51 == total_offset_14 ? phv_data_81 : _GEN_7944; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7946 = 8'h52 == total_offset_14 ? phv_data_82 : _GEN_7945; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7947 = 8'h53 == total_offset_14 ? phv_data_83 : _GEN_7946; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7948 = 8'h54 == total_offset_14 ? phv_data_84 : _GEN_7947; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7949 = 8'h55 == total_offset_14 ? phv_data_85 : _GEN_7948; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7950 = 8'h56 == total_offset_14 ? phv_data_86 : _GEN_7949; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7951 = 8'h57 == total_offset_14 ? phv_data_87 : _GEN_7950; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7952 = 8'h58 == total_offset_14 ? phv_data_88 : _GEN_7951; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7953 = 8'h59 == total_offset_14 ? phv_data_89 : _GEN_7952; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7954 = 8'h5a == total_offset_14 ? phv_data_90 : _GEN_7953; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7955 = 8'h5b == total_offset_14 ? phv_data_91 : _GEN_7954; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7956 = 8'h5c == total_offset_14 ? phv_data_92 : _GEN_7955; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7957 = 8'h5d == total_offset_14 ? phv_data_93 : _GEN_7956; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7958 = 8'h5e == total_offset_14 ? phv_data_94 : _GEN_7957; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7959 = 8'h5f == total_offset_14 ? phv_data_95 : _GEN_7958; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7960 = 8'h60 == total_offset_14 ? phv_data_96 : _GEN_7959; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7961 = 8'h61 == total_offset_14 ? phv_data_97 : _GEN_7960; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7962 = 8'h62 == total_offset_14 ? phv_data_98 : _GEN_7961; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7963 = 8'h63 == total_offset_14 ? phv_data_99 : _GEN_7962; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7964 = 8'h64 == total_offset_14 ? phv_data_100 : _GEN_7963; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7965 = 8'h65 == total_offset_14 ? phv_data_101 : _GEN_7964; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7966 = 8'h66 == total_offset_14 ? phv_data_102 : _GEN_7965; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7967 = 8'h67 == total_offset_14 ? phv_data_103 : _GEN_7966; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7968 = 8'h68 == total_offset_14 ? phv_data_104 : _GEN_7967; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7969 = 8'h69 == total_offset_14 ? phv_data_105 : _GEN_7968; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7970 = 8'h6a == total_offset_14 ? phv_data_106 : _GEN_7969; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7971 = 8'h6b == total_offset_14 ? phv_data_107 : _GEN_7970; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7972 = 8'h6c == total_offset_14 ? phv_data_108 : _GEN_7971; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7973 = 8'h6d == total_offset_14 ? phv_data_109 : _GEN_7972; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7974 = 8'h6e == total_offset_14 ? phv_data_110 : _GEN_7973; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7975 = 8'h6f == total_offset_14 ? phv_data_111 : _GEN_7974; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7976 = 8'h70 == total_offset_14 ? phv_data_112 : _GEN_7975; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7977 = 8'h71 == total_offset_14 ? phv_data_113 : _GEN_7976; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7978 = 8'h72 == total_offset_14 ? phv_data_114 : _GEN_7977; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7979 = 8'h73 == total_offset_14 ? phv_data_115 : _GEN_7978; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7980 = 8'h74 == total_offset_14 ? phv_data_116 : _GEN_7979; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7981 = 8'h75 == total_offset_14 ? phv_data_117 : _GEN_7980; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7982 = 8'h76 == total_offset_14 ? phv_data_118 : _GEN_7981; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7983 = 8'h77 == total_offset_14 ? phv_data_119 : _GEN_7982; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7984 = 8'h78 == total_offset_14 ? phv_data_120 : _GEN_7983; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7985 = 8'h79 == total_offset_14 ? phv_data_121 : _GEN_7984; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7986 = 8'h7a == total_offset_14 ? phv_data_122 : _GEN_7985; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7987 = 8'h7b == total_offset_14 ? phv_data_123 : _GEN_7986; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7988 = 8'h7c == total_offset_14 ? phv_data_124 : _GEN_7987; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7989 = 8'h7d == total_offset_14 ? phv_data_125 : _GEN_7988; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7990 = 8'h7e == total_offset_14 ? phv_data_126 : _GEN_7989; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7991 = 8'h7f == total_offset_14 ? phv_data_127 : _GEN_7990; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7992 = 8'h80 == total_offset_14 ? phv_data_128 : _GEN_7991; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7993 = 8'h81 == total_offset_14 ? phv_data_129 : _GEN_7992; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7994 = 8'h82 == total_offset_14 ? phv_data_130 : _GEN_7993; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7995 = 8'h83 == total_offset_14 ? phv_data_131 : _GEN_7994; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7996 = 8'h84 == total_offset_14 ? phv_data_132 : _GEN_7995; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7997 = 8'h85 == total_offset_14 ? phv_data_133 : _GEN_7996; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7998 = 8'h86 == total_offset_14 ? phv_data_134 : _GEN_7997; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_7999 = 8'h87 == total_offset_14 ? phv_data_135 : _GEN_7998; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8000 = 8'h88 == total_offset_14 ? phv_data_136 : _GEN_7999; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8001 = 8'h89 == total_offset_14 ? phv_data_137 : _GEN_8000; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8002 = 8'h8a == total_offset_14 ? phv_data_138 : _GEN_8001; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8003 = 8'h8b == total_offset_14 ? phv_data_139 : _GEN_8002; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8004 = 8'h8c == total_offset_14 ? phv_data_140 : _GEN_8003; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8005 = 8'h8d == total_offset_14 ? phv_data_141 : _GEN_8004; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8006 = 8'h8e == total_offset_14 ? phv_data_142 : _GEN_8005; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8007 = 8'h8f == total_offset_14 ? phv_data_143 : _GEN_8006; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8008 = 8'h90 == total_offset_14 ? phv_data_144 : _GEN_8007; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8009 = 8'h91 == total_offset_14 ? phv_data_145 : _GEN_8008; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8010 = 8'h92 == total_offset_14 ? phv_data_146 : _GEN_8009; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8011 = 8'h93 == total_offset_14 ? phv_data_147 : _GEN_8010; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8012 = 8'h94 == total_offset_14 ? phv_data_148 : _GEN_8011; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8013 = 8'h95 == total_offset_14 ? phv_data_149 : _GEN_8012; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8014 = 8'h96 == total_offset_14 ? phv_data_150 : _GEN_8013; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8015 = 8'h97 == total_offset_14 ? phv_data_151 : _GEN_8014; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8016 = 8'h98 == total_offset_14 ? phv_data_152 : _GEN_8015; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8017 = 8'h99 == total_offset_14 ? phv_data_153 : _GEN_8016; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8018 = 8'h9a == total_offset_14 ? phv_data_154 : _GEN_8017; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8019 = 8'h9b == total_offset_14 ? phv_data_155 : _GEN_8018; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8020 = 8'h9c == total_offset_14 ? phv_data_156 : _GEN_8019; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8021 = 8'h9d == total_offset_14 ? phv_data_157 : _GEN_8020; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8022 = 8'h9e == total_offset_14 ? phv_data_158 : _GEN_8021; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8023 = 8'h9f == total_offset_14 ? phv_data_159 : _GEN_8022; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8024 = 8'ha0 == total_offset_14 ? phv_data_160 : _GEN_8023; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8025 = 8'ha1 == total_offset_14 ? phv_data_161 : _GEN_8024; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8026 = 8'ha2 == total_offset_14 ? phv_data_162 : _GEN_8025; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8027 = 8'ha3 == total_offset_14 ? phv_data_163 : _GEN_8026; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8028 = 8'ha4 == total_offset_14 ? phv_data_164 : _GEN_8027; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8029 = 8'ha5 == total_offset_14 ? phv_data_165 : _GEN_8028; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8030 = 8'ha6 == total_offset_14 ? phv_data_166 : _GEN_8029; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8031 = 8'ha7 == total_offset_14 ? phv_data_167 : _GEN_8030; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8032 = 8'ha8 == total_offset_14 ? phv_data_168 : _GEN_8031; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8033 = 8'ha9 == total_offset_14 ? phv_data_169 : _GEN_8032; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8034 = 8'haa == total_offset_14 ? phv_data_170 : _GEN_8033; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8035 = 8'hab == total_offset_14 ? phv_data_171 : _GEN_8034; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8036 = 8'hac == total_offset_14 ? phv_data_172 : _GEN_8035; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8037 = 8'had == total_offset_14 ? phv_data_173 : _GEN_8036; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8038 = 8'hae == total_offset_14 ? phv_data_174 : _GEN_8037; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8039 = 8'haf == total_offset_14 ? phv_data_175 : _GEN_8038; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8040 = 8'hb0 == total_offset_14 ? phv_data_176 : _GEN_8039; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8041 = 8'hb1 == total_offset_14 ? phv_data_177 : _GEN_8040; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8042 = 8'hb2 == total_offset_14 ? phv_data_178 : _GEN_8041; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8043 = 8'hb3 == total_offset_14 ? phv_data_179 : _GEN_8042; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8044 = 8'hb4 == total_offset_14 ? phv_data_180 : _GEN_8043; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8045 = 8'hb5 == total_offset_14 ? phv_data_181 : _GEN_8044; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8046 = 8'hb6 == total_offset_14 ? phv_data_182 : _GEN_8045; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8047 = 8'hb7 == total_offset_14 ? phv_data_183 : _GEN_8046; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8048 = 8'hb8 == total_offset_14 ? phv_data_184 : _GEN_8047; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8049 = 8'hb9 == total_offset_14 ? phv_data_185 : _GEN_8048; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8050 = 8'hba == total_offset_14 ? phv_data_186 : _GEN_8049; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8051 = 8'hbb == total_offset_14 ? phv_data_187 : _GEN_8050; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8052 = 8'hbc == total_offset_14 ? phv_data_188 : _GEN_8051; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8053 = 8'hbd == total_offset_14 ? phv_data_189 : _GEN_8052; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8054 = 8'hbe == total_offset_14 ? phv_data_190 : _GEN_8053; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8055 = 8'hbf == total_offset_14 ? phv_data_191 : _GEN_8054; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8056 = 8'hc0 == total_offset_14 ? phv_data_192 : _GEN_8055; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8057 = 8'hc1 == total_offset_14 ? phv_data_193 : _GEN_8056; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8058 = 8'hc2 == total_offset_14 ? phv_data_194 : _GEN_8057; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8059 = 8'hc3 == total_offset_14 ? phv_data_195 : _GEN_8058; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8060 = 8'hc4 == total_offset_14 ? phv_data_196 : _GEN_8059; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8061 = 8'hc5 == total_offset_14 ? phv_data_197 : _GEN_8060; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8062 = 8'hc6 == total_offset_14 ? phv_data_198 : _GEN_8061; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8063 = 8'hc7 == total_offset_14 ? phv_data_199 : _GEN_8062; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8064 = 8'hc8 == total_offset_14 ? phv_data_200 : _GEN_8063; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8065 = 8'hc9 == total_offset_14 ? phv_data_201 : _GEN_8064; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8066 = 8'hca == total_offset_14 ? phv_data_202 : _GEN_8065; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8067 = 8'hcb == total_offset_14 ? phv_data_203 : _GEN_8066; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8068 = 8'hcc == total_offset_14 ? phv_data_204 : _GEN_8067; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8069 = 8'hcd == total_offset_14 ? phv_data_205 : _GEN_8068; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8070 = 8'hce == total_offset_14 ? phv_data_206 : _GEN_8069; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8071 = 8'hcf == total_offset_14 ? phv_data_207 : _GEN_8070; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8072 = 8'hd0 == total_offset_14 ? phv_data_208 : _GEN_8071; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8073 = 8'hd1 == total_offset_14 ? phv_data_209 : _GEN_8072; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8074 = 8'hd2 == total_offset_14 ? phv_data_210 : _GEN_8073; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8075 = 8'hd3 == total_offset_14 ? phv_data_211 : _GEN_8074; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8076 = 8'hd4 == total_offset_14 ? phv_data_212 : _GEN_8075; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8077 = 8'hd5 == total_offset_14 ? phv_data_213 : _GEN_8076; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8078 = 8'hd6 == total_offset_14 ? phv_data_214 : _GEN_8077; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8079 = 8'hd7 == total_offset_14 ? phv_data_215 : _GEN_8078; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8080 = 8'hd8 == total_offset_14 ? phv_data_216 : _GEN_8079; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8081 = 8'hd9 == total_offset_14 ? phv_data_217 : _GEN_8080; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8082 = 8'hda == total_offset_14 ? phv_data_218 : _GEN_8081; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8083 = 8'hdb == total_offset_14 ? phv_data_219 : _GEN_8082; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8084 = 8'hdc == total_offset_14 ? phv_data_220 : _GEN_8083; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8085 = 8'hdd == total_offset_14 ? phv_data_221 : _GEN_8084; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8086 = 8'hde == total_offset_14 ? phv_data_222 : _GEN_8085; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8087 = 8'hdf == total_offset_14 ? phv_data_223 : _GEN_8086; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8088 = 8'he0 == total_offset_14 ? phv_data_224 : _GEN_8087; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8089 = 8'he1 == total_offset_14 ? phv_data_225 : _GEN_8088; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8090 = 8'he2 == total_offset_14 ? phv_data_226 : _GEN_8089; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8091 = 8'he3 == total_offset_14 ? phv_data_227 : _GEN_8090; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8092 = 8'he4 == total_offset_14 ? phv_data_228 : _GEN_8091; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8093 = 8'he5 == total_offset_14 ? phv_data_229 : _GEN_8092; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8094 = 8'he6 == total_offset_14 ? phv_data_230 : _GEN_8093; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8095 = 8'he7 == total_offset_14 ? phv_data_231 : _GEN_8094; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8096 = 8'he8 == total_offset_14 ? phv_data_232 : _GEN_8095; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8097 = 8'he9 == total_offset_14 ? phv_data_233 : _GEN_8096; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8098 = 8'hea == total_offset_14 ? phv_data_234 : _GEN_8097; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8099 = 8'heb == total_offset_14 ? phv_data_235 : _GEN_8098; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8100 = 8'hec == total_offset_14 ? phv_data_236 : _GEN_8099; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8101 = 8'hed == total_offset_14 ? phv_data_237 : _GEN_8100; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8102 = 8'hee == total_offset_14 ? phv_data_238 : _GEN_8101; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8103 = 8'hef == total_offset_14 ? phv_data_239 : _GEN_8102; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8104 = 8'hf0 == total_offset_14 ? phv_data_240 : _GEN_8103; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8105 = 8'hf1 == total_offset_14 ? phv_data_241 : _GEN_8104; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8106 = 8'hf2 == total_offset_14 ? phv_data_242 : _GEN_8105; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8107 = 8'hf3 == total_offset_14 ? phv_data_243 : _GEN_8106; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8108 = 8'hf4 == total_offset_14 ? phv_data_244 : _GEN_8107; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8109 = 8'hf5 == total_offset_14 ? phv_data_245 : _GEN_8108; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8110 = 8'hf6 == total_offset_14 ? phv_data_246 : _GEN_8109; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8111 = 8'hf7 == total_offset_14 ? phv_data_247 : _GEN_8110; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8112 = 8'hf8 == total_offset_14 ? phv_data_248 : _GEN_8111; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8113 = 8'hf9 == total_offset_14 ? phv_data_249 : _GEN_8112; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8114 = 8'hfa == total_offset_14 ? phv_data_250 : _GEN_8113; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8115 = 8'hfb == total_offset_14 ? phv_data_251 : _GEN_8114; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8116 = 8'hfc == total_offset_14 ? phv_data_252 : _GEN_8115; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8117 = 8'hfd == total_offset_14 ? phv_data_253 : _GEN_8116; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8118 = 8'hfe == total_offset_14 ? phv_data_254 : _GEN_8117; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8119 = 8'hff == total_offset_14 ? phv_data_255 : _GEN_8118; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_12726 = {{1'd0}, total_offset_14}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8120 = 9'h100 == _GEN_12726 ? phv_data_256 : _GEN_8119; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8121 = 9'h101 == _GEN_12726 ? phv_data_257 : _GEN_8120; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8122 = 9'h102 == _GEN_12726 ? phv_data_258 : _GEN_8121; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8123 = 9'h103 == _GEN_12726 ? phv_data_259 : _GEN_8122; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8124 = 9'h104 == _GEN_12726 ? phv_data_260 : _GEN_8123; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8125 = 9'h105 == _GEN_12726 ? phv_data_261 : _GEN_8124; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8126 = 9'h106 == _GEN_12726 ? phv_data_262 : _GEN_8125; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8127 = 9'h107 == _GEN_12726 ? phv_data_263 : _GEN_8126; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8128 = 9'h108 == _GEN_12726 ? phv_data_264 : _GEN_8127; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8129 = 9'h109 == _GEN_12726 ? phv_data_265 : _GEN_8128; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8130 = 9'h10a == _GEN_12726 ? phv_data_266 : _GEN_8129; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8131 = 9'h10b == _GEN_12726 ? phv_data_267 : _GEN_8130; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8132 = 9'h10c == _GEN_12726 ? phv_data_268 : _GEN_8131; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8133 = 9'h10d == _GEN_12726 ? phv_data_269 : _GEN_8132; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8134 = 9'h10e == _GEN_12726 ? phv_data_270 : _GEN_8133; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8135 = 9'h10f == _GEN_12726 ? phv_data_271 : _GEN_8134; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8136 = 9'h110 == _GEN_12726 ? phv_data_272 : _GEN_8135; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8137 = 9'h111 == _GEN_12726 ? phv_data_273 : _GEN_8136; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8138 = 9'h112 == _GEN_12726 ? phv_data_274 : _GEN_8137; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8139 = 9'h113 == _GEN_12726 ? phv_data_275 : _GEN_8138; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8140 = 9'h114 == _GEN_12726 ? phv_data_276 : _GEN_8139; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8141 = 9'h115 == _GEN_12726 ? phv_data_277 : _GEN_8140; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8142 = 9'h116 == _GEN_12726 ? phv_data_278 : _GEN_8141; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8143 = 9'h117 == _GEN_12726 ? phv_data_279 : _GEN_8142; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8144 = 9'h118 == _GEN_12726 ? phv_data_280 : _GEN_8143; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8145 = 9'h119 == _GEN_12726 ? phv_data_281 : _GEN_8144; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8146 = 9'h11a == _GEN_12726 ? phv_data_282 : _GEN_8145; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8147 = 9'h11b == _GEN_12726 ? phv_data_283 : _GEN_8146; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8148 = 9'h11c == _GEN_12726 ? phv_data_284 : _GEN_8147; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8149 = 9'h11d == _GEN_12726 ? phv_data_285 : _GEN_8148; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8150 = 9'h11e == _GEN_12726 ? phv_data_286 : _GEN_8149; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8151 = 9'h11f == _GEN_12726 ? phv_data_287 : _GEN_8150; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8152 = 9'h120 == _GEN_12726 ? phv_data_288 : _GEN_8151; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8153 = 9'h121 == _GEN_12726 ? phv_data_289 : _GEN_8152; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8154 = 9'h122 == _GEN_12726 ? phv_data_290 : _GEN_8153; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8155 = 9'h123 == _GEN_12726 ? phv_data_291 : _GEN_8154; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8156 = 9'h124 == _GEN_12726 ? phv_data_292 : _GEN_8155; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8157 = 9'h125 == _GEN_12726 ? phv_data_293 : _GEN_8156; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8158 = 9'h126 == _GEN_12726 ? phv_data_294 : _GEN_8157; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8159 = 9'h127 == _GEN_12726 ? phv_data_295 : _GEN_8158; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8160 = 9'h128 == _GEN_12726 ? phv_data_296 : _GEN_8159; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8161 = 9'h129 == _GEN_12726 ? phv_data_297 : _GEN_8160; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8162 = 9'h12a == _GEN_12726 ? phv_data_298 : _GEN_8161; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8163 = 9'h12b == _GEN_12726 ? phv_data_299 : _GEN_8162; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8164 = 9'h12c == _GEN_12726 ? phv_data_300 : _GEN_8163; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8165 = 9'h12d == _GEN_12726 ? phv_data_301 : _GEN_8164; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8166 = 9'h12e == _GEN_12726 ? phv_data_302 : _GEN_8165; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8167 = 9'h12f == _GEN_12726 ? phv_data_303 : _GEN_8166; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8168 = 9'h130 == _GEN_12726 ? phv_data_304 : _GEN_8167; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8169 = 9'h131 == _GEN_12726 ? phv_data_305 : _GEN_8168; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8170 = 9'h132 == _GEN_12726 ? phv_data_306 : _GEN_8169; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8171 = 9'h133 == _GEN_12726 ? phv_data_307 : _GEN_8170; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8172 = 9'h134 == _GEN_12726 ? phv_data_308 : _GEN_8171; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8173 = 9'h135 == _GEN_12726 ? phv_data_309 : _GEN_8172; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8174 = 9'h136 == _GEN_12726 ? phv_data_310 : _GEN_8173; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8175 = 9'h137 == _GEN_12726 ? phv_data_311 : _GEN_8174; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8176 = 9'h138 == _GEN_12726 ? phv_data_312 : _GEN_8175; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8177 = 9'h139 == _GEN_12726 ? phv_data_313 : _GEN_8176; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8178 = 9'h13a == _GEN_12726 ? phv_data_314 : _GEN_8177; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8179 = 9'h13b == _GEN_12726 ? phv_data_315 : _GEN_8178; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8180 = 9'h13c == _GEN_12726 ? phv_data_316 : _GEN_8179; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8181 = 9'h13d == _GEN_12726 ? phv_data_317 : _GEN_8180; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8182 = 9'h13e == _GEN_12726 ? phv_data_318 : _GEN_8181; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8183 = 9'h13f == _GEN_12726 ? phv_data_319 : _GEN_8182; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8184 = 9'h140 == _GEN_12726 ? phv_data_320 : _GEN_8183; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8185 = 9'h141 == _GEN_12726 ? phv_data_321 : _GEN_8184; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8186 = 9'h142 == _GEN_12726 ? phv_data_322 : _GEN_8185; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8187 = 9'h143 == _GEN_12726 ? phv_data_323 : _GEN_8186; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8188 = 9'h144 == _GEN_12726 ? phv_data_324 : _GEN_8187; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8189 = 9'h145 == _GEN_12726 ? phv_data_325 : _GEN_8188; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8190 = 9'h146 == _GEN_12726 ? phv_data_326 : _GEN_8189; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8191 = 9'h147 == _GEN_12726 ? phv_data_327 : _GEN_8190; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8192 = 9'h148 == _GEN_12726 ? phv_data_328 : _GEN_8191; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8193 = 9'h149 == _GEN_12726 ? phv_data_329 : _GEN_8192; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8194 = 9'h14a == _GEN_12726 ? phv_data_330 : _GEN_8193; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8195 = 9'h14b == _GEN_12726 ? phv_data_331 : _GEN_8194; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8196 = 9'h14c == _GEN_12726 ? phv_data_332 : _GEN_8195; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8197 = 9'h14d == _GEN_12726 ? phv_data_333 : _GEN_8196; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8198 = 9'h14e == _GEN_12726 ? phv_data_334 : _GEN_8197; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8199 = 9'h14f == _GEN_12726 ? phv_data_335 : _GEN_8198; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8200 = 9'h150 == _GEN_12726 ? phv_data_336 : _GEN_8199; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8201 = 9'h151 == _GEN_12726 ? phv_data_337 : _GEN_8200; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8202 = 9'h152 == _GEN_12726 ? phv_data_338 : _GEN_8201; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8203 = 9'h153 == _GEN_12726 ? phv_data_339 : _GEN_8202; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8204 = 9'h154 == _GEN_12726 ? phv_data_340 : _GEN_8203; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8205 = 9'h155 == _GEN_12726 ? phv_data_341 : _GEN_8204; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8206 = 9'h156 == _GEN_12726 ? phv_data_342 : _GEN_8205; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8207 = 9'h157 == _GEN_12726 ? phv_data_343 : _GEN_8206; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8208 = 9'h158 == _GEN_12726 ? phv_data_344 : _GEN_8207; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8209 = 9'h159 == _GEN_12726 ? phv_data_345 : _GEN_8208; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8210 = 9'h15a == _GEN_12726 ? phv_data_346 : _GEN_8209; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8211 = 9'h15b == _GEN_12726 ? phv_data_347 : _GEN_8210; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8212 = 9'h15c == _GEN_12726 ? phv_data_348 : _GEN_8211; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8213 = 9'h15d == _GEN_12726 ? phv_data_349 : _GEN_8212; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8214 = 9'h15e == _GEN_12726 ? phv_data_350 : _GEN_8213; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8215 = 9'h15f == _GEN_12726 ? phv_data_351 : _GEN_8214; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8216 = 9'h160 == _GEN_12726 ? phv_data_352 : _GEN_8215; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8217 = 9'h161 == _GEN_12726 ? phv_data_353 : _GEN_8216; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8218 = 9'h162 == _GEN_12726 ? phv_data_354 : _GEN_8217; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8219 = 9'h163 == _GEN_12726 ? phv_data_355 : _GEN_8218; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8220 = 9'h164 == _GEN_12726 ? phv_data_356 : _GEN_8219; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8221 = 9'h165 == _GEN_12726 ? phv_data_357 : _GEN_8220; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8222 = 9'h166 == _GEN_12726 ? phv_data_358 : _GEN_8221; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8223 = 9'h167 == _GEN_12726 ? phv_data_359 : _GEN_8222; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8224 = 9'h168 == _GEN_12726 ? phv_data_360 : _GEN_8223; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8225 = 9'h169 == _GEN_12726 ? phv_data_361 : _GEN_8224; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8226 = 9'h16a == _GEN_12726 ? phv_data_362 : _GEN_8225; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8227 = 9'h16b == _GEN_12726 ? phv_data_363 : _GEN_8226; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8228 = 9'h16c == _GEN_12726 ? phv_data_364 : _GEN_8227; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8229 = 9'h16d == _GEN_12726 ? phv_data_365 : _GEN_8228; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8230 = 9'h16e == _GEN_12726 ? phv_data_366 : _GEN_8229; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8231 = 9'h16f == _GEN_12726 ? phv_data_367 : _GEN_8230; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8232 = 9'h170 == _GEN_12726 ? phv_data_368 : _GEN_8231; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8233 = 9'h171 == _GEN_12726 ? phv_data_369 : _GEN_8232; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8234 = 9'h172 == _GEN_12726 ? phv_data_370 : _GEN_8233; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8235 = 9'h173 == _GEN_12726 ? phv_data_371 : _GEN_8234; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8236 = 9'h174 == _GEN_12726 ? phv_data_372 : _GEN_8235; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8237 = 9'h175 == _GEN_12726 ? phv_data_373 : _GEN_8236; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8238 = 9'h176 == _GEN_12726 ? phv_data_374 : _GEN_8237; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8239 = 9'h177 == _GEN_12726 ? phv_data_375 : _GEN_8238; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8240 = 9'h178 == _GEN_12726 ? phv_data_376 : _GEN_8239; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8241 = 9'h179 == _GEN_12726 ? phv_data_377 : _GEN_8240; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8242 = 9'h17a == _GEN_12726 ? phv_data_378 : _GEN_8241; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8243 = 9'h17b == _GEN_12726 ? phv_data_379 : _GEN_8242; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8244 = 9'h17c == _GEN_12726 ? phv_data_380 : _GEN_8243; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8245 = 9'h17d == _GEN_12726 ? phv_data_381 : _GEN_8244; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8246 = 9'h17e == _GEN_12726 ? phv_data_382 : _GEN_8245; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8247 = 9'h17f == _GEN_12726 ? phv_data_383 : _GEN_8246; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8248 = 9'h180 == _GEN_12726 ? phv_data_384 : _GEN_8247; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8249 = 9'h181 == _GEN_12726 ? phv_data_385 : _GEN_8248; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8250 = 9'h182 == _GEN_12726 ? phv_data_386 : _GEN_8249; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8251 = 9'h183 == _GEN_12726 ? phv_data_387 : _GEN_8250; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8252 = 9'h184 == _GEN_12726 ? phv_data_388 : _GEN_8251; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8253 = 9'h185 == _GEN_12726 ? phv_data_389 : _GEN_8252; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8254 = 9'h186 == _GEN_12726 ? phv_data_390 : _GEN_8253; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8255 = 9'h187 == _GEN_12726 ? phv_data_391 : _GEN_8254; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8256 = 9'h188 == _GEN_12726 ? phv_data_392 : _GEN_8255; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8257 = 9'h189 == _GEN_12726 ? phv_data_393 : _GEN_8256; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8258 = 9'h18a == _GEN_12726 ? phv_data_394 : _GEN_8257; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8259 = 9'h18b == _GEN_12726 ? phv_data_395 : _GEN_8258; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8260 = 9'h18c == _GEN_12726 ? phv_data_396 : _GEN_8259; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8261 = 9'h18d == _GEN_12726 ? phv_data_397 : _GEN_8260; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8262 = 9'h18e == _GEN_12726 ? phv_data_398 : _GEN_8261; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8263 = 9'h18f == _GEN_12726 ? phv_data_399 : _GEN_8262; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8264 = 9'h190 == _GEN_12726 ? phv_data_400 : _GEN_8263; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8265 = 9'h191 == _GEN_12726 ? phv_data_401 : _GEN_8264; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8266 = 9'h192 == _GEN_12726 ? phv_data_402 : _GEN_8265; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8267 = 9'h193 == _GEN_12726 ? phv_data_403 : _GEN_8266; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8268 = 9'h194 == _GEN_12726 ? phv_data_404 : _GEN_8267; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8269 = 9'h195 == _GEN_12726 ? phv_data_405 : _GEN_8268; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8270 = 9'h196 == _GEN_12726 ? phv_data_406 : _GEN_8269; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8271 = 9'h197 == _GEN_12726 ? phv_data_407 : _GEN_8270; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8272 = 9'h198 == _GEN_12726 ? phv_data_408 : _GEN_8271; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8273 = 9'h199 == _GEN_12726 ? phv_data_409 : _GEN_8272; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8274 = 9'h19a == _GEN_12726 ? phv_data_410 : _GEN_8273; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8275 = 9'h19b == _GEN_12726 ? phv_data_411 : _GEN_8274; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8276 = 9'h19c == _GEN_12726 ? phv_data_412 : _GEN_8275; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8277 = 9'h19d == _GEN_12726 ? phv_data_413 : _GEN_8276; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8278 = 9'h19e == _GEN_12726 ? phv_data_414 : _GEN_8277; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8279 = 9'h19f == _GEN_12726 ? phv_data_415 : _GEN_8278; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8280 = 9'h1a0 == _GEN_12726 ? phv_data_416 : _GEN_8279; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8281 = 9'h1a1 == _GEN_12726 ? phv_data_417 : _GEN_8280; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8282 = 9'h1a2 == _GEN_12726 ? phv_data_418 : _GEN_8281; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8283 = 9'h1a3 == _GEN_12726 ? phv_data_419 : _GEN_8282; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8284 = 9'h1a4 == _GEN_12726 ? phv_data_420 : _GEN_8283; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8285 = 9'h1a5 == _GEN_12726 ? phv_data_421 : _GEN_8284; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8286 = 9'h1a6 == _GEN_12726 ? phv_data_422 : _GEN_8285; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8287 = 9'h1a7 == _GEN_12726 ? phv_data_423 : _GEN_8286; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8288 = 9'h1a8 == _GEN_12726 ? phv_data_424 : _GEN_8287; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8289 = 9'h1a9 == _GEN_12726 ? phv_data_425 : _GEN_8288; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8290 = 9'h1aa == _GEN_12726 ? phv_data_426 : _GEN_8289; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8291 = 9'h1ab == _GEN_12726 ? phv_data_427 : _GEN_8290; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8292 = 9'h1ac == _GEN_12726 ? phv_data_428 : _GEN_8291; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8293 = 9'h1ad == _GEN_12726 ? phv_data_429 : _GEN_8292; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8294 = 9'h1ae == _GEN_12726 ? phv_data_430 : _GEN_8293; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8295 = 9'h1af == _GEN_12726 ? phv_data_431 : _GEN_8294; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8296 = 9'h1b0 == _GEN_12726 ? phv_data_432 : _GEN_8295; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8297 = 9'h1b1 == _GEN_12726 ? phv_data_433 : _GEN_8296; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8298 = 9'h1b2 == _GEN_12726 ? phv_data_434 : _GEN_8297; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8299 = 9'h1b3 == _GEN_12726 ? phv_data_435 : _GEN_8298; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8300 = 9'h1b4 == _GEN_12726 ? phv_data_436 : _GEN_8299; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8301 = 9'h1b5 == _GEN_12726 ? phv_data_437 : _GEN_8300; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8302 = 9'h1b6 == _GEN_12726 ? phv_data_438 : _GEN_8301; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8303 = 9'h1b7 == _GEN_12726 ? phv_data_439 : _GEN_8302; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8304 = 9'h1b8 == _GEN_12726 ? phv_data_440 : _GEN_8303; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8305 = 9'h1b9 == _GEN_12726 ? phv_data_441 : _GEN_8304; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8306 = 9'h1ba == _GEN_12726 ? phv_data_442 : _GEN_8305; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8307 = 9'h1bb == _GEN_12726 ? phv_data_443 : _GEN_8306; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8308 = 9'h1bc == _GEN_12726 ? phv_data_444 : _GEN_8307; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8309 = 9'h1bd == _GEN_12726 ? phv_data_445 : _GEN_8308; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8310 = 9'h1be == _GEN_12726 ? phv_data_446 : _GEN_8309; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8311 = 9'h1bf == _GEN_12726 ? phv_data_447 : _GEN_8310; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8312 = 9'h1c0 == _GEN_12726 ? phv_data_448 : _GEN_8311; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8313 = 9'h1c1 == _GEN_12726 ? phv_data_449 : _GEN_8312; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8314 = 9'h1c2 == _GEN_12726 ? phv_data_450 : _GEN_8313; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8315 = 9'h1c3 == _GEN_12726 ? phv_data_451 : _GEN_8314; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8316 = 9'h1c4 == _GEN_12726 ? phv_data_452 : _GEN_8315; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8317 = 9'h1c5 == _GEN_12726 ? phv_data_453 : _GEN_8316; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8318 = 9'h1c6 == _GEN_12726 ? phv_data_454 : _GEN_8317; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8319 = 9'h1c7 == _GEN_12726 ? phv_data_455 : _GEN_8318; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8320 = 9'h1c8 == _GEN_12726 ? phv_data_456 : _GEN_8319; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8321 = 9'h1c9 == _GEN_12726 ? phv_data_457 : _GEN_8320; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8322 = 9'h1ca == _GEN_12726 ? phv_data_458 : _GEN_8321; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8323 = 9'h1cb == _GEN_12726 ? phv_data_459 : _GEN_8322; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8324 = 9'h1cc == _GEN_12726 ? phv_data_460 : _GEN_8323; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8325 = 9'h1cd == _GEN_12726 ? phv_data_461 : _GEN_8324; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8326 = 9'h1ce == _GEN_12726 ? phv_data_462 : _GEN_8325; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8327 = 9'h1cf == _GEN_12726 ? phv_data_463 : _GEN_8326; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8328 = 9'h1d0 == _GEN_12726 ? phv_data_464 : _GEN_8327; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8329 = 9'h1d1 == _GEN_12726 ? phv_data_465 : _GEN_8328; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8330 = 9'h1d2 == _GEN_12726 ? phv_data_466 : _GEN_8329; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8331 = 9'h1d3 == _GEN_12726 ? phv_data_467 : _GEN_8330; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8332 = 9'h1d4 == _GEN_12726 ? phv_data_468 : _GEN_8331; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8333 = 9'h1d5 == _GEN_12726 ? phv_data_469 : _GEN_8332; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8334 = 9'h1d6 == _GEN_12726 ? phv_data_470 : _GEN_8333; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8335 = 9'h1d7 == _GEN_12726 ? phv_data_471 : _GEN_8334; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8336 = 9'h1d8 == _GEN_12726 ? phv_data_472 : _GEN_8335; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8337 = 9'h1d9 == _GEN_12726 ? phv_data_473 : _GEN_8336; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8338 = 9'h1da == _GEN_12726 ? phv_data_474 : _GEN_8337; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8339 = 9'h1db == _GEN_12726 ? phv_data_475 : _GEN_8338; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8340 = 9'h1dc == _GEN_12726 ? phv_data_476 : _GEN_8339; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8341 = 9'h1dd == _GEN_12726 ? phv_data_477 : _GEN_8340; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8342 = 9'h1de == _GEN_12726 ? phv_data_478 : _GEN_8341; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8343 = 9'h1df == _GEN_12726 ? phv_data_479 : _GEN_8342; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8344 = 9'h1e0 == _GEN_12726 ? phv_data_480 : _GEN_8343; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8345 = 9'h1e1 == _GEN_12726 ? phv_data_481 : _GEN_8344; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8346 = 9'h1e2 == _GEN_12726 ? phv_data_482 : _GEN_8345; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8347 = 9'h1e3 == _GEN_12726 ? phv_data_483 : _GEN_8346; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8348 = 9'h1e4 == _GEN_12726 ? phv_data_484 : _GEN_8347; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8349 = 9'h1e5 == _GEN_12726 ? phv_data_485 : _GEN_8348; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8350 = 9'h1e6 == _GEN_12726 ? phv_data_486 : _GEN_8349; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8351 = 9'h1e7 == _GEN_12726 ? phv_data_487 : _GEN_8350; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8352 = 9'h1e8 == _GEN_12726 ? phv_data_488 : _GEN_8351; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8353 = 9'h1e9 == _GEN_12726 ? phv_data_489 : _GEN_8352; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8354 = 9'h1ea == _GEN_12726 ? phv_data_490 : _GEN_8353; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8355 = 9'h1eb == _GEN_12726 ? phv_data_491 : _GEN_8354; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8356 = 9'h1ec == _GEN_12726 ? phv_data_492 : _GEN_8355; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8357 = 9'h1ed == _GEN_12726 ? phv_data_493 : _GEN_8356; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8358 = 9'h1ee == _GEN_12726 ? phv_data_494 : _GEN_8357; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8359 = 9'h1ef == _GEN_12726 ? phv_data_495 : _GEN_8358; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8360 = 9'h1f0 == _GEN_12726 ? phv_data_496 : _GEN_8359; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8361 = 9'h1f1 == _GEN_12726 ? phv_data_497 : _GEN_8360; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8362 = 9'h1f2 == _GEN_12726 ? phv_data_498 : _GEN_8361; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8363 = 9'h1f3 == _GEN_12726 ? phv_data_499 : _GEN_8362; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8364 = 9'h1f4 == _GEN_12726 ? phv_data_500 : _GEN_8363; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8365 = 9'h1f5 == _GEN_12726 ? phv_data_501 : _GEN_8364; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8366 = 9'h1f6 == _GEN_12726 ? phv_data_502 : _GEN_8365; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8367 = 9'h1f7 == _GEN_12726 ? phv_data_503 : _GEN_8366; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8368 = 9'h1f8 == _GEN_12726 ? phv_data_504 : _GEN_8367; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8369 = 9'h1f9 == _GEN_12726 ? phv_data_505 : _GEN_8368; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8370 = 9'h1fa == _GEN_12726 ? phv_data_506 : _GEN_8369; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8371 = 9'h1fb == _GEN_12726 ? phv_data_507 : _GEN_8370; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8372 = 9'h1fc == _GEN_12726 ? phv_data_508 : _GEN_8371; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8373 = 9'h1fd == _GEN_12726 ? phv_data_509 : _GEN_8372; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8374 = 9'h1fe == _GEN_12726 ? phv_data_510 : _GEN_8373; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_1 = 9'h1ff == _GEN_12726 ? phv_data_511 : _GEN_8374; // @[executor.scala 197:66 executor.scala 197:66]
  wire  mask_3_1 = 2'h2 >= offset_3[1:0] & (2'h2 < ending_3 | ending_3 == 2'h0); // @[executor.scala 199:56]
  wire [7:0] total_offset_15 = {total_offset_hi_3,2'h3}; // @[Cat.scala 30:58]
  wire [7:0] _GEN_8377 = 8'h1 == total_offset_15 ? phv_data_1 : phv_data_0; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8378 = 8'h2 == total_offset_15 ? phv_data_2 : _GEN_8377; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8379 = 8'h3 == total_offset_15 ? phv_data_3 : _GEN_8378; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8380 = 8'h4 == total_offset_15 ? phv_data_4 : _GEN_8379; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8381 = 8'h5 == total_offset_15 ? phv_data_5 : _GEN_8380; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8382 = 8'h6 == total_offset_15 ? phv_data_6 : _GEN_8381; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8383 = 8'h7 == total_offset_15 ? phv_data_7 : _GEN_8382; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8384 = 8'h8 == total_offset_15 ? phv_data_8 : _GEN_8383; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8385 = 8'h9 == total_offset_15 ? phv_data_9 : _GEN_8384; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8386 = 8'ha == total_offset_15 ? phv_data_10 : _GEN_8385; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8387 = 8'hb == total_offset_15 ? phv_data_11 : _GEN_8386; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8388 = 8'hc == total_offset_15 ? phv_data_12 : _GEN_8387; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8389 = 8'hd == total_offset_15 ? phv_data_13 : _GEN_8388; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8390 = 8'he == total_offset_15 ? phv_data_14 : _GEN_8389; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8391 = 8'hf == total_offset_15 ? phv_data_15 : _GEN_8390; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8392 = 8'h10 == total_offset_15 ? phv_data_16 : _GEN_8391; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8393 = 8'h11 == total_offset_15 ? phv_data_17 : _GEN_8392; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8394 = 8'h12 == total_offset_15 ? phv_data_18 : _GEN_8393; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8395 = 8'h13 == total_offset_15 ? phv_data_19 : _GEN_8394; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8396 = 8'h14 == total_offset_15 ? phv_data_20 : _GEN_8395; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8397 = 8'h15 == total_offset_15 ? phv_data_21 : _GEN_8396; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8398 = 8'h16 == total_offset_15 ? phv_data_22 : _GEN_8397; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8399 = 8'h17 == total_offset_15 ? phv_data_23 : _GEN_8398; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8400 = 8'h18 == total_offset_15 ? phv_data_24 : _GEN_8399; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8401 = 8'h19 == total_offset_15 ? phv_data_25 : _GEN_8400; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8402 = 8'h1a == total_offset_15 ? phv_data_26 : _GEN_8401; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8403 = 8'h1b == total_offset_15 ? phv_data_27 : _GEN_8402; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8404 = 8'h1c == total_offset_15 ? phv_data_28 : _GEN_8403; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8405 = 8'h1d == total_offset_15 ? phv_data_29 : _GEN_8404; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8406 = 8'h1e == total_offset_15 ? phv_data_30 : _GEN_8405; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8407 = 8'h1f == total_offset_15 ? phv_data_31 : _GEN_8406; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8408 = 8'h20 == total_offset_15 ? phv_data_32 : _GEN_8407; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8409 = 8'h21 == total_offset_15 ? phv_data_33 : _GEN_8408; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8410 = 8'h22 == total_offset_15 ? phv_data_34 : _GEN_8409; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8411 = 8'h23 == total_offset_15 ? phv_data_35 : _GEN_8410; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8412 = 8'h24 == total_offset_15 ? phv_data_36 : _GEN_8411; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8413 = 8'h25 == total_offset_15 ? phv_data_37 : _GEN_8412; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8414 = 8'h26 == total_offset_15 ? phv_data_38 : _GEN_8413; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8415 = 8'h27 == total_offset_15 ? phv_data_39 : _GEN_8414; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8416 = 8'h28 == total_offset_15 ? phv_data_40 : _GEN_8415; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8417 = 8'h29 == total_offset_15 ? phv_data_41 : _GEN_8416; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8418 = 8'h2a == total_offset_15 ? phv_data_42 : _GEN_8417; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8419 = 8'h2b == total_offset_15 ? phv_data_43 : _GEN_8418; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8420 = 8'h2c == total_offset_15 ? phv_data_44 : _GEN_8419; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8421 = 8'h2d == total_offset_15 ? phv_data_45 : _GEN_8420; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8422 = 8'h2e == total_offset_15 ? phv_data_46 : _GEN_8421; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8423 = 8'h2f == total_offset_15 ? phv_data_47 : _GEN_8422; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8424 = 8'h30 == total_offset_15 ? phv_data_48 : _GEN_8423; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8425 = 8'h31 == total_offset_15 ? phv_data_49 : _GEN_8424; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8426 = 8'h32 == total_offset_15 ? phv_data_50 : _GEN_8425; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8427 = 8'h33 == total_offset_15 ? phv_data_51 : _GEN_8426; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8428 = 8'h34 == total_offset_15 ? phv_data_52 : _GEN_8427; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8429 = 8'h35 == total_offset_15 ? phv_data_53 : _GEN_8428; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8430 = 8'h36 == total_offset_15 ? phv_data_54 : _GEN_8429; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8431 = 8'h37 == total_offset_15 ? phv_data_55 : _GEN_8430; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8432 = 8'h38 == total_offset_15 ? phv_data_56 : _GEN_8431; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8433 = 8'h39 == total_offset_15 ? phv_data_57 : _GEN_8432; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8434 = 8'h3a == total_offset_15 ? phv_data_58 : _GEN_8433; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8435 = 8'h3b == total_offset_15 ? phv_data_59 : _GEN_8434; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8436 = 8'h3c == total_offset_15 ? phv_data_60 : _GEN_8435; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8437 = 8'h3d == total_offset_15 ? phv_data_61 : _GEN_8436; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8438 = 8'h3e == total_offset_15 ? phv_data_62 : _GEN_8437; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8439 = 8'h3f == total_offset_15 ? phv_data_63 : _GEN_8438; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8440 = 8'h40 == total_offset_15 ? phv_data_64 : _GEN_8439; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8441 = 8'h41 == total_offset_15 ? phv_data_65 : _GEN_8440; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8442 = 8'h42 == total_offset_15 ? phv_data_66 : _GEN_8441; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8443 = 8'h43 == total_offset_15 ? phv_data_67 : _GEN_8442; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8444 = 8'h44 == total_offset_15 ? phv_data_68 : _GEN_8443; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8445 = 8'h45 == total_offset_15 ? phv_data_69 : _GEN_8444; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8446 = 8'h46 == total_offset_15 ? phv_data_70 : _GEN_8445; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8447 = 8'h47 == total_offset_15 ? phv_data_71 : _GEN_8446; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8448 = 8'h48 == total_offset_15 ? phv_data_72 : _GEN_8447; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8449 = 8'h49 == total_offset_15 ? phv_data_73 : _GEN_8448; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8450 = 8'h4a == total_offset_15 ? phv_data_74 : _GEN_8449; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8451 = 8'h4b == total_offset_15 ? phv_data_75 : _GEN_8450; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8452 = 8'h4c == total_offset_15 ? phv_data_76 : _GEN_8451; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8453 = 8'h4d == total_offset_15 ? phv_data_77 : _GEN_8452; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8454 = 8'h4e == total_offset_15 ? phv_data_78 : _GEN_8453; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8455 = 8'h4f == total_offset_15 ? phv_data_79 : _GEN_8454; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8456 = 8'h50 == total_offset_15 ? phv_data_80 : _GEN_8455; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8457 = 8'h51 == total_offset_15 ? phv_data_81 : _GEN_8456; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8458 = 8'h52 == total_offset_15 ? phv_data_82 : _GEN_8457; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8459 = 8'h53 == total_offset_15 ? phv_data_83 : _GEN_8458; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8460 = 8'h54 == total_offset_15 ? phv_data_84 : _GEN_8459; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8461 = 8'h55 == total_offset_15 ? phv_data_85 : _GEN_8460; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8462 = 8'h56 == total_offset_15 ? phv_data_86 : _GEN_8461; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8463 = 8'h57 == total_offset_15 ? phv_data_87 : _GEN_8462; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8464 = 8'h58 == total_offset_15 ? phv_data_88 : _GEN_8463; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8465 = 8'h59 == total_offset_15 ? phv_data_89 : _GEN_8464; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8466 = 8'h5a == total_offset_15 ? phv_data_90 : _GEN_8465; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8467 = 8'h5b == total_offset_15 ? phv_data_91 : _GEN_8466; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8468 = 8'h5c == total_offset_15 ? phv_data_92 : _GEN_8467; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8469 = 8'h5d == total_offset_15 ? phv_data_93 : _GEN_8468; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8470 = 8'h5e == total_offset_15 ? phv_data_94 : _GEN_8469; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8471 = 8'h5f == total_offset_15 ? phv_data_95 : _GEN_8470; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8472 = 8'h60 == total_offset_15 ? phv_data_96 : _GEN_8471; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8473 = 8'h61 == total_offset_15 ? phv_data_97 : _GEN_8472; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8474 = 8'h62 == total_offset_15 ? phv_data_98 : _GEN_8473; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8475 = 8'h63 == total_offset_15 ? phv_data_99 : _GEN_8474; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8476 = 8'h64 == total_offset_15 ? phv_data_100 : _GEN_8475; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8477 = 8'h65 == total_offset_15 ? phv_data_101 : _GEN_8476; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8478 = 8'h66 == total_offset_15 ? phv_data_102 : _GEN_8477; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8479 = 8'h67 == total_offset_15 ? phv_data_103 : _GEN_8478; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8480 = 8'h68 == total_offset_15 ? phv_data_104 : _GEN_8479; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8481 = 8'h69 == total_offset_15 ? phv_data_105 : _GEN_8480; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8482 = 8'h6a == total_offset_15 ? phv_data_106 : _GEN_8481; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8483 = 8'h6b == total_offset_15 ? phv_data_107 : _GEN_8482; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8484 = 8'h6c == total_offset_15 ? phv_data_108 : _GEN_8483; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8485 = 8'h6d == total_offset_15 ? phv_data_109 : _GEN_8484; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8486 = 8'h6e == total_offset_15 ? phv_data_110 : _GEN_8485; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8487 = 8'h6f == total_offset_15 ? phv_data_111 : _GEN_8486; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8488 = 8'h70 == total_offset_15 ? phv_data_112 : _GEN_8487; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8489 = 8'h71 == total_offset_15 ? phv_data_113 : _GEN_8488; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8490 = 8'h72 == total_offset_15 ? phv_data_114 : _GEN_8489; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8491 = 8'h73 == total_offset_15 ? phv_data_115 : _GEN_8490; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8492 = 8'h74 == total_offset_15 ? phv_data_116 : _GEN_8491; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8493 = 8'h75 == total_offset_15 ? phv_data_117 : _GEN_8492; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8494 = 8'h76 == total_offset_15 ? phv_data_118 : _GEN_8493; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8495 = 8'h77 == total_offset_15 ? phv_data_119 : _GEN_8494; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8496 = 8'h78 == total_offset_15 ? phv_data_120 : _GEN_8495; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8497 = 8'h79 == total_offset_15 ? phv_data_121 : _GEN_8496; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8498 = 8'h7a == total_offset_15 ? phv_data_122 : _GEN_8497; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8499 = 8'h7b == total_offset_15 ? phv_data_123 : _GEN_8498; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8500 = 8'h7c == total_offset_15 ? phv_data_124 : _GEN_8499; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8501 = 8'h7d == total_offset_15 ? phv_data_125 : _GEN_8500; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8502 = 8'h7e == total_offset_15 ? phv_data_126 : _GEN_8501; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8503 = 8'h7f == total_offset_15 ? phv_data_127 : _GEN_8502; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8504 = 8'h80 == total_offset_15 ? phv_data_128 : _GEN_8503; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8505 = 8'h81 == total_offset_15 ? phv_data_129 : _GEN_8504; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8506 = 8'h82 == total_offset_15 ? phv_data_130 : _GEN_8505; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8507 = 8'h83 == total_offset_15 ? phv_data_131 : _GEN_8506; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8508 = 8'h84 == total_offset_15 ? phv_data_132 : _GEN_8507; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8509 = 8'h85 == total_offset_15 ? phv_data_133 : _GEN_8508; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8510 = 8'h86 == total_offset_15 ? phv_data_134 : _GEN_8509; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8511 = 8'h87 == total_offset_15 ? phv_data_135 : _GEN_8510; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8512 = 8'h88 == total_offset_15 ? phv_data_136 : _GEN_8511; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8513 = 8'h89 == total_offset_15 ? phv_data_137 : _GEN_8512; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8514 = 8'h8a == total_offset_15 ? phv_data_138 : _GEN_8513; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8515 = 8'h8b == total_offset_15 ? phv_data_139 : _GEN_8514; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8516 = 8'h8c == total_offset_15 ? phv_data_140 : _GEN_8515; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8517 = 8'h8d == total_offset_15 ? phv_data_141 : _GEN_8516; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8518 = 8'h8e == total_offset_15 ? phv_data_142 : _GEN_8517; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8519 = 8'h8f == total_offset_15 ? phv_data_143 : _GEN_8518; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8520 = 8'h90 == total_offset_15 ? phv_data_144 : _GEN_8519; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8521 = 8'h91 == total_offset_15 ? phv_data_145 : _GEN_8520; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8522 = 8'h92 == total_offset_15 ? phv_data_146 : _GEN_8521; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8523 = 8'h93 == total_offset_15 ? phv_data_147 : _GEN_8522; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8524 = 8'h94 == total_offset_15 ? phv_data_148 : _GEN_8523; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8525 = 8'h95 == total_offset_15 ? phv_data_149 : _GEN_8524; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8526 = 8'h96 == total_offset_15 ? phv_data_150 : _GEN_8525; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8527 = 8'h97 == total_offset_15 ? phv_data_151 : _GEN_8526; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8528 = 8'h98 == total_offset_15 ? phv_data_152 : _GEN_8527; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8529 = 8'h99 == total_offset_15 ? phv_data_153 : _GEN_8528; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8530 = 8'h9a == total_offset_15 ? phv_data_154 : _GEN_8529; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8531 = 8'h9b == total_offset_15 ? phv_data_155 : _GEN_8530; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8532 = 8'h9c == total_offset_15 ? phv_data_156 : _GEN_8531; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8533 = 8'h9d == total_offset_15 ? phv_data_157 : _GEN_8532; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8534 = 8'h9e == total_offset_15 ? phv_data_158 : _GEN_8533; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8535 = 8'h9f == total_offset_15 ? phv_data_159 : _GEN_8534; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8536 = 8'ha0 == total_offset_15 ? phv_data_160 : _GEN_8535; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8537 = 8'ha1 == total_offset_15 ? phv_data_161 : _GEN_8536; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8538 = 8'ha2 == total_offset_15 ? phv_data_162 : _GEN_8537; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8539 = 8'ha3 == total_offset_15 ? phv_data_163 : _GEN_8538; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8540 = 8'ha4 == total_offset_15 ? phv_data_164 : _GEN_8539; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8541 = 8'ha5 == total_offset_15 ? phv_data_165 : _GEN_8540; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8542 = 8'ha6 == total_offset_15 ? phv_data_166 : _GEN_8541; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8543 = 8'ha7 == total_offset_15 ? phv_data_167 : _GEN_8542; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8544 = 8'ha8 == total_offset_15 ? phv_data_168 : _GEN_8543; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8545 = 8'ha9 == total_offset_15 ? phv_data_169 : _GEN_8544; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8546 = 8'haa == total_offset_15 ? phv_data_170 : _GEN_8545; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8547 = 8'hab == total_offset_15 ? phv_data_171 : _GEN_8546; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8548 = 8'hac == total_offset_15 ? phv_data_172 : _GEN_8547; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8549 = 8'had == total_offset_15 ? phv_data_173 : _GEN_8548; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8550 = 8'hae == total_offset_15 ? phv_data_174 : _GEN_8549; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8551 = 8'haf == total_offset_15 ? phv_data_175 : _GEN_8550; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8552 = 8'hb0 == total_offset_15 ? phv_data_176 : _GEN_8551; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8553 = 8'hb1 == total_offset_15 ? phv_data_177 : _GEN_8552; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8554 = 8'hb2 == total_offset_15 ? phv_data_178 : _GEN_8553; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8555 = 8'hb3 == total_offset_15 ? phv_data_179 : _GEN_8554; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8556 = 8'hb4 == total_offset_15 ? phv_data_180 : _GEN_8555; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8557 = 8'hb5 == total_offset_15 ? phv_data_181 : _GEN_8556; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8558 = 8'hb6 == total_offset_15 ? phv_data_182 : _GEN_8557; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8559 = 8'hb7 == total_offset_15 ? phv_data_183 : _GEN_8558; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8560 = 8'hb8 == total_offset_15 ? phv_data_184 : _GEN_8559; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8561 = 8'hb9 == total_offset_15 ? phv_data_185 : _GEN_8560; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8562 = 8'hba == total_offset_15 ? phv_data_186 : _GEN_8561; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8563 = 8'hbb == total_offset_15 ? phv_data_187 : _GEN_8562; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8564 = 8'hbc == total_offset_15 ? phv_data_188 : _GEN_8563; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8565 = 8'hbd == total_offset_15 ? phv_data_189 : _GEN_8564; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8566 = 8'hbe == total_offset_15 ? phv_data_190 : _GEN_8565; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8567 = 8'hbf == total_offset_15 ? phv_data_191 : _GEN_8566; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8568 = 8'hc0 == total_offset_15 ? phv_data_192 : _GEN_8567; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8569 = 8'hc1 == total_offset_15 ? phv_data_193 : _GEN_8568; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8570 = 8'hc2 == total_offset_15 ? phv_data_194 : _GEN_8569; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8571 = 8'hc3 == total_offset_15 ? phv_data_195 : _GEN_8570; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8572 = 8'hc4 == total_offset_15 ? phv_data_196 : _GEN_8571; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8573 = 8'hc5 == total_offset_15 ? phv_data_197 : _GEN_8572; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8574 = 8'hc6 == total_offset_15 ? phv_data_198 : _GEN_8573; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8575 = 8'hc7 == total_offset_15 ? phv_data_199 : _GEN_8574; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8576 = 8'hc8 == total_offset_15 ? phv_data_200 : _GEN_8575; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8577 = 8'hc9 == total_offset_15 ? phv_data_201 : _GEN_8576; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8578 = 8'hca == total_offset_15 ? phv_data_202 : _GEN_8577; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8579 = 8'hcb == total_offset_15 ? phv_data_203 : _GEN_8578; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8580 = 8'hcc == total_offset_15 ? phv_data_204 : _GEN_8579; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8581 = 8'hcd == total_offset_15 ? phv_data_205 : _GEN_8580; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8582 = 8'hce == total_offset_15 ? phv_data_206 : _GEN_8581; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8583 = 8'hcf == total_offset_15 ? phv_data_207 : _GEN_8582; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8584 = 8'hd0 == total_offset_15 ? phv_data_208 : _GEN_8583; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8585 = 8'hd1 == total_offset_15 ? phv_data_209 : _GEN_8584; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8586 = 8'hd2 == total_offset_15 ? phv_data_210 : _GEN_8585; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8587 = 8'hd3 == total_offset_15 ? phv_data_211 : _GEN_8586; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8588 = 8'hd4 == total_offset_15 ? phv_data_212 : _GEN_8587; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8589 = 8'hd5 == total_offset_15 ? phv_data_213 : _GEN_8588; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8590 = 8'hd6 == total_offset_15 ? phv_data_214 : _GEN_8589; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8591 = 8'hd7 == total_offset_15 ? phv_data_215 : _GEN_8590; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8592 = 8'hd8 == total_offset_15 ? phv_data_216 : _GEN_8591; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8593 = 8'hd9 == total_offset_15 ? phv_data_217 : _GEN_8592; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8594 = 8'hda == total_offset_15 ? phv_data_218 : _GEN_8593; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8595 = 8'hdb == total_offset_15 ? phv_data_219 : _GEN_8594; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8596 = 8'hdc == total_offset_15 ? phv_data_220 : _GEN_8595; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8597 = 8'hdd == total_offset_15 ? phv_data_221 : _GEN_8596; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8598 = 8'hde == total_offset_15 ? phv_data_222 : _GEN_8597; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8599 = 8'hdf == total_offset_15 ? phv_data_223 : _GEN_8598; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8600 = 8'he0 == total_offset_15 ? phv_data_224 : _GEN_8599; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8601 = 8'he1 == total_offset_15 ? phv_data_225 : _GEN_8600; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8602 = 8'he2 == total_offset_15 ? phv_data_226 : _GEN_8601; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8603 = 8'he3 == total_offset_15 ? phv_data_227 : _GEN_8602; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8604 = 8'he4 == total_offset_15 ? phv_data_228 : _GEN_8603; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8605 = 8'he5 == total_offset_15 ? phv_data_229 : _GEN_8604; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8606 = 8'he6 == total_offset_15 ? phv_data_230 : _GEN_8605; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8607 = 8'he7 == total_offset_15 ? phv_data_231 : _GEN_8606; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8608 = 8'he8 == total_offset_15 ? phv_data_232 : _GEN_8607; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8609 = 8'he9 == total_offset_15 ? phv_data_233 : _GEN_8608; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8610 = 8'hea == total_offset_15 ? phv_data_234 : _GEN_8609; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8611 = 8'heb == total_offset_15 ? phv_data_235 : _GEN_8610; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8612 = 8'hec == total_offset_15 ? phv_data_236 : _GEN_8611; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8613 = 8'hed == total_offset_15 ? phv_data_237 : _GEN_8612; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8614 = 8'hee == total_offset_15 ? phv_data_238 : _GEN_8613; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8615 = 8'hef == total_offset_15 ? phv_data_239 : _GEN_8614; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8616 = 8'hf0 == total_offset_15 ? phv_data_240 : _GEN_8615; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8617 = 8'hf1 == total_offset_15 ? phv_data_241 : _GEN_8616; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8618 = 8'hf2 == total_offset_15 ? phv_data_242 : _GEN_8617; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8619 = 8'hf3 == total_offset_15 ? phv_data_243 : _GEN_8618; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8620 = 8'hf4 == total_offset_15 ? phv_data_244 : _GEN_8619; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8621 = 8'hf5 == total_offset_15 ? phv_data_245 : _GEN_8620; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8622 = 8'hf6 == total_offset_15 ? phv_data_246 : _GEN_8621; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8623 = 8'hf7 == total_offset_15 ? phv_data_247 : _GEN_8622; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8624 = 8'hf8 == total_offset_15 ? phv_data_248 : _GEN_8623; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8625 = 8'hf9 == total_offset_15 ? phv_data_249 : _GEN_8624; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8626 = 8'hfa == total_offset_15 ? phv_data_250 : _GEN_8625; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8627 = 8'hfb == total_offset_15 ? phv_data_251 : _GEN_8626; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8628 = 8'hfc == total_offset_15 ? phv_data_252 : _GEN_8627; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8629 = 8'hfd == total_offset_15 ? phv_data_253 : _GEN_8628; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8630 = 8'hfe == total_offset_15 ? phv_data_254 : _GEN_8629; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8631 = 8'hff == total_offset_15 ? phv_data_255 : _GEN_8630; // @[executor.scala 197:66 executor.scala 197:66]
  wire [8:0] _GEN_12982 = {{1'd0}, total_offset_15}; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8632 = 9'h100 == _GEN_12982 ? phv_data_256 : _GEN_8631; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8633 = 9'h101 == _GEN_12982 ? phv_data_257 : _GEN_8632; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8634 = 9'h102 == _GEN_12982 ? phv_data_258 : _GEN_8633; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8635 = 9'h103 == _GEN_12982 ? phv_data_259 : _GEN_8634; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8636 = 9'h104 == _GEN_12982 ? phv_data_260 : _GEN_8635; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8637 = 9'h105 == _GEN_12982 ? phv_data_261 : _GEN_8636; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8638 = 9'h106 == _GEN_12982 ? phv_data_262 : _GEN_8637; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8639 = 9'h107 == _GEN_12982 ? phv_data_263 : _GEN_8638; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8640 = 9'h108 == _GEN_12982 ? phv_data_264 : _GEN_8639; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8641 = 9'h109 == _GEN_12982 ? phv_data_265 : _GEN_8640; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8642 = 9'h10a == _GEN_12982 ? phv_data_266 : _GEN_8641; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8643 = 9'h10b == _GEN_12982 ? phv_data_267 : _GEN_8642; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8644 = 9'h10c == _GEN_12982 ? phv_data_268 : _GEN_8643; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8645 = 9'h10d == _GEN_12982 ? phv_data_269 : _GEN_8644; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8646 = 9'h10e == _GEN_12982 ? phv_data_270 : _GEN_8645; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8647 = 9'h10f == _GEN_12982 ? phv_data_271 : _GEN_8646; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8648 = 9'h110 == _GEN_12982 ? phv_data_272 : _GEN_8647; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8649 = 9'h111 == _GEN_12982 ? phv_data_273 : _GEN_8648; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8650 = 9'h112 == _GEN_12982 ? phv_data_274 : _GEN_8649; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8651 = 9'h113 == _GEN_12982 ? phv_data_275 : _GEN_8650; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8652 = 9'h114 == _GEN_12982 ? phv_data_276 : _GEN_8651; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8653 = 9'h115 == _GEN_12982 ? phv_data_277 : _GEN_8652; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8654 = 9'h116 == _GEN_12982 ? phv_data_278 : _GEN_8653; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8655 = 9'h117 == _GEN_12982 ? phv_data_279 : _GEN_8654; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8656 = 9'h118 == _GEN_12982 ? phv_data_280 : _GEN_8655; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8657 = 9'h119 == _GEN_12982 ? phv_data_281 : _GEN_8656; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8658 = 9'h11a == _GEN_12982 ? phv_data_282 : _GEN_8657; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8659 = 9'h11b == _GEN_12982 ? phv_data_283 : _GEN_8658; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8660 = 9'h11c == _GEN_12982 ? phv_data_284 : _GEN_8659; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8661 = 9'h11d == _GEN_12982 ? phv_data_285 : _GEN_8660; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8662 = 9'h11e == _GEN_12982 ? phv_data_286 : _GEN_8661; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8663 = 9'h11f == _GEN_12982 ? phv_data_287 : _GEN_8662; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8664 = 9'h120 == _GEN_12982 ? phv_data_288 : _GEN_8663; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8665 = 9'h121 == _GEN_12982 ? phv_data_289 : _GEN_8664; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8666 = 9'h122 == _GEN_12982 ? phv_data_290 : _GEN_8665; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8667 = 9'h123 == _GEN_12982 ? phv_data_291 : _GEN_8666; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8668 = 9'h124 == _GEN_12982 ? phv_data_292 : _GEN_8667; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8669 = 9'h125 == _GEN_12982 ? phv_data_293 : _GEN_8668; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8670 = 9'h126 == _GEN_12982 ? phv_data_294 : _GEN_8669; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8671 = 9'h127 == _GEN_12982 ? phv_data_295 : _GEN_8670; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8672 = 9'h128 == _GEN_12982 ? phv_data_296 : _GEN_8671; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8673 = 9'h129 == _GEN_12982 ? phv_data_297 : _GEN_8672; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8674 = 9'h12a == _GEN_12982 ? phv_data_298 : _GEN_8673; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8675 = 9'h12b == _GEN_12982 ? phv_data_299 : _GEN_8674; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8676 = 9'h12c == _GEN_12982 ? phv_data_300 : _GEN_8675; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8677 = 9'h12d == _GEN_12982 ? phv_data_301 : _GEN_8676; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8678 = 9'h12e == _GEN_12982 ? phv_data_302 : _GEN_8677; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8679 = 9'h12f == _GEN_12982 ? phv_data_303 : _GEN_8678; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8680 = 9'h130 == _GEN_12982 ? phv_data_304 : _GEN_8679; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8681 = 9'h131 == _GEN_12982 ? phv_data_305 : _GEN_8680; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8682 = 9'h132 == _GEN_12982 ? phv_data_306 : _GEN_8681; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8683 = 9'h133 == _GEN_12982 ? phv_data_307 : _GEN_8682; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8684 = 9'h134 == _GEN_12982 ? phv_data_308 : _GEN_8683; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8685 = 9'h135 == _GEN_12982 ? phv_data_309 : _GEN_8684; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8686 = 9'h136 == _GEN_12982 ? phv_data_310 : _GEN_8685; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8687 = 9'h137 == _GEN_12982 ? phv_data_311 : _GEN_8686; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8688 = 9'h138 == _GEN_12982 ? phv_data_312 : _GEN_8687; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8689 = 9'h139 == _GEN_12982 ? phv_data_313 : _GEN_8688; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8690 = 9'h13a == _GEN_12982 ? phv_data_314 : _GEN_8689; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8691 = 9'h13b == _GEN_12982 ? phv_data_315 : _GEN_8690; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8692 = 9'h13c == _GEN_12982 ? phv_data_316 : _GEN_8691; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8693 = 9'h13d == _GEN_12982 ? phv_data_317 : _GEN_8692; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8694 = 9'h13e == _GEN_12982 ? phv_data_318 : _GEN_8693; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8695 = 9'h13f == _GEN_12982 ? phv_data_319 : _GEN_8694; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8696 = 9'h140 == _GEN_12982 ? phv_data_320 : _GEN_8695; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8697 = 9'h141 == _GEN_12982 ? phv_data_321 : _GEN_8696; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8698 = 9'h142 == _GEN_12982 ? phv_data_322 : _GEN_8697; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8699 = 9'h143 == _GEN_12982 ? phv_data_323 : _GEN_8698; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8700 = 9'h144 == _GEN_12982 ? phv_data_324 : _GEN_8699; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8701 = 9'h145 == _GEN_12982 ? phv_data_325 : _GEN_8700; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8702 = 9'h146 == _GEN_12982 ? phv_data_326 : _GEN_8701; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8703 = 9'h147 == _GEN_12982 ? phv_data_327 : _GEN_8702; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8704 = 9'h148 == _GEN_12982 ? phv_data_328 : _GEN_8703; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8705 = 9'h149 == _GEN_12982 ? phv_data_329 : _GEN_8704; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8706 = 9'h14a == _GEN_12982 ? phv_data_330 : _GEN_8705; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8707 = 9'h14b == _GEN_12982 ? phv_data_331 : _GEN_8706; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8708 = 9'h14c == _GEN_12982 ? phv_data_332 : _GEN_8707; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8709 = 9'h14d == _GEN_12982 ? phv_data_333 : _GEN_8708; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8710 = 9'h14e == _GEN_12982 ? phv_data_334 : _GEN_8709; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8711 = 9'h14f == _GEN_12982 ? phv_data_335 : _GEN_8710; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8712 = 9'h150 == _GEN_12982 ? phv_data_336 : _GEN_8711; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8713 = 9'h151 == _GEN_12982 ? phv_data_337 : _GEN_8712; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8714 = 9'h152 == _GEN_12982 ? phv_data_338 : _GEN_8713; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8715 = 9'h153 == _GEN_12982 ? phv_data_339 : _GEN_8714; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8716 = 9'h154 == _GEN_12982 ? phv_data_340 : _GEN_8715; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8717 = 9'h155 == _GEN_12982 ? phv_data_341 : _GEN_8716; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8718 = 9'h156 == _GEN_12982 ? phv_data_342 : _GEN_8717; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8719 = 9'h157 == _GEN_12982 ? phv_data_343 : _GEN_8718; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8720 = 9'h158 == _GEN_12982 ? phv_data_344 : _GEN_8719; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8721 = 9'h159 == _GEN_12982 ? phv_data_345 : _GEN_8720; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8722 = 9'h15a == _GEN_12982 ? phv_data_346 : _GEN_8721; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8723 = 9'h15b == _GEN_12982 ? phv_data_347 : _GEN_8722; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8724 = 9'h15c == _GEN_12982 ? phv_data_348 : _GEN_8723; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8725 = 9'h15d == _GEN_12982 ? phv_data_349 : _GEN_8724; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8726 = 9'h15e == _GEN_12982 ? phv_data_350 : _GEN_8725; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8727 = 9'h15f == _GEN_12982 ? phv_data_351 : _GEN_8726; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8728 = 9'h160 == _GEN_12982 ? phv_data_352 : _GEN_8727; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8729 = 9'h161 == _GEN_12982 ? phv_data_353 : _GEN_8728; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8730 = 9'h162 == _GEN_12982 ? phv_data_354 : _GEN_8729; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8731 = 9'h163 == _GEN_12982 ? phv_data_355 : _GEN_8730; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8732 = 9'h164 == _GEN_12982 ? phv_data_356 : _GEN_8731; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8733 = 9'h165 == _GEN_12982 ? phv_data_357 : _GEN_8732; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8734 = 9'h166 == _GEN_12982 ? phv_data_358 : _GEN_8733; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8735 = 9'h167 == _GEN_12982 ? phv_data_359 : _GEN_8734; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8736 = 9'h168 == _GEN_12982 ? phv_data_360 : _GEN_8735; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8737 = 9'h169 == _GEN_12982 ? phv_data_361 : _GEN_8736; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8738 = 9'h16a == _GEN_12982 ? phv_data_362 : _GEN_8737; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8739 = 9'h16b == _GEN_12982 ? phv_data_363 : _GEN_8738; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8740 = 9'h16c == _GEN_12982 ? phv_data_364 : _GEN_8739; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8741 = 9'h16d == _GEN_12982 ? phv_data_365 : _GEN_8740; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8742 = 9'h16e == _GEN_12982 ? phv_data_366 : _GEN_8741; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8743 = 9'h16f == _GEN_12982 ? phv_data_367 : _GEN_8742; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8744 = 9'h170 == _GEN_12982 ? phv_data_368 : _GEN_8743; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8745 = 9'h171 == _GEN_12982 ? phv_data_369 : _GEN_8744; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8746 = 9'h172 == _GEN_12982 ? phv_data_370 : _GEN_8745; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8747 = 9'h173 == _GEN_12982 ? phv_data_371 : _GEN_8746; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8748 = 9'h174 == _GEN_12982 ? phv_data_372 : _GEN_8747; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8749 = 9'h175 == _GEN_12982 ? phv_data_373 : _GEN_8748; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8750 = 9'h176 == _GEN_12982 ? phv_data_374 : _GEN_8749; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8751 = 9'h177 == _GEN_12982 ? phv_data_375 : _GEN_8750; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8752 = 9'h178 == _GEN_12982 ? phv_data_376 : _GEN_8751; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8753 = 9'h179 == _GEN_12982 ? phv_data_377 : _GEN_8752; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8754 = 9'h17a == _GEN_12982 ? phv_data_378 : _GEN_8753; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8755 = 9'h17b == _GEN_12982 ? phv_data_379 : _GEN_8754; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8756 = 9'h17c == _GEN_12982 ? phv_data_380 : _GEN_8755; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8757 = 9'h17d == _GEN_12982 ? phv_data_381 : _GEN_8756; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8758 = 9'h17e == _GEN_12982 ? phv_data_382 : _GEN_8757; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8759 = 9'h17f == _GEN_12982 ? phv_data_383 : _GEN_8758; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8760 = 9'h180 == _GEN_12982 ? phv_data_384 : _GEN_8759; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8761 = 9'h181 == _GEN_12982 ? phv_data_385 : _GEN_8760; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8762 = 9'h182 == _GEN_12982 ? phv_data_386 : _GEN_8761; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8763 = 9'h183 == _GEN_12982 ? phv_data_387 : _GEN_8762; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8764 = 9'h184 == _GEN_12982 ? phv_data_388 : _GEN_8763; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8765 = 9'h185 == _GEN_12982 ? phv_data_389 : _GEN_8764; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8766 = 9'h186 == _GEN_12982 ? phv_data_390 : _GEN_8765; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8767 = 9'h187 == _GEN_12982 ? phv_data_391 : _GEN_8766; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8768 = 9'h188 == _GEN_12982 ? phv_data_392 : _GEN_8767; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8769 = 9'h189 == _GEN_12982 ? phv_data_393 : _GEN_8768; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8770 = 9'h18a == _GEN_12982 ? phv_data_394 : _GEN_8769; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8771 = 9'h18b == _GEN_12982 ? phv_data_395 : _GEN_8770; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8772 = 9'h18c == _GEN_12982 ? phv_data_396 : _GEN_8771; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8773 = 9'h18d == _GEN_12982 ? phv_data_397 : _GEN_8772; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8774 = 9'h18e == _GEN_12982 ? phv_data_398 : _GEN_8773; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8775 = 9'h18f == _GEN_12982 ? phv_data_399 : _GEN_8774; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8776 = 9'h190 == _GEN_12982 ? phv_data_400 : _GEN_8775; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8777 = 9'h191 == _GEN_12982 ? phv_data_401 : _GEN_8776; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8778 = 9'h192 == _GEN_12982 ? phv_data_402 : _GEN_8777; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8779 = 9'h193 == _GEN_12982 ? phv_data_403 : _GEN_8778; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8780 = 9'h194 == _GEN_12982 ? phv_data_404 : _GEN_8779; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8781 = 9'h195 == _GEN_12982 ? phv_data_405 : _GEN_8780; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8782 = 9'h196 == _GEN_12982 ? phv_data_406 : _GEN_8781; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8783 = 9'h197 == _GEN_12982 ? phv_data_407 : _GEN_8782; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8784 = 9'h198 == _GEN_12982 ? phv_data_408 : _GEN_8783; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8785 = 9'h199 == _GEN_12982 ? phv_data_409 : _GEN_8784; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8786 = 9'h19a == _GEN_12982 ? phv_data_410 : _GEN_8785; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8787 = 9'h19b == _GEN_12982 ? phv_data_411 : _GEN_8786; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8788 = 9'h19c == _GEN_12982 ? phv_data_412 : _GEN_8787; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8789 = 9'h19d == _GEN_12982 ? phv_data_413 : _GEN_8788; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8790 = 9'h19e == _GEN_12982 ? phv_data_414 : _GEN_8789; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8791 = 9'h19f == _GEN_12982 ? phv_data_415 : _GEN_8790; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8792 = 9'h1a0 == _GEN_12982 ? phv_data_416 : _GEN_8791; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8793 = 9'h1a1 == _GEN_12982 ? phv_data_417 : _GEN_8792; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8794 = 9'h1a2 == _GEN_12982 ? phv_data_418 : _GEN_8793; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8795 = 9'h1a3 == _GEN_12982 ? phv_data_419 : _GEN_8794; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8796 = 9'h1a4 == _GEN_12982 ? phv_data_420 : _GEN_8795; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8797 = 9'h1a5 == _GEN_12982 ? phv_data_421 : _GEN_8796; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8798 = 9'h1a6 == _GEN_12982 ? phv_data_422 : _GEN_8797; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8799 = 9'h1a7 == _GEN_12982 ? phv_data_423 : _GEN_8798; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8800 = 9'h1a8 == _GEN_12982 ? phv_data_424 : _GEN_8799; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8801 = 9'h1a9 == _GEN_12982 ? phv_data_425 : _GEN_8800; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8802 = 9'h1aa == _GEN_12982 ? phv_data_426 : _GEN_8801; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8803 = 9'h1ab == _GEN_12982 ? phv_data_427 : _GEN_8802; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8804 = 9'h1ac == _GEN_12982 ? phv_data_428 : _GEN_8803; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8805 = 9'h1ad == _GEN_12982 ? phv_data_429 : _GEN_8804; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8806 = 9'h1ae == _GEN_12982 ? phv_data_430 : _GEN_8805; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8807 = 9'h1af == _GEN_12982 ? phv_data_431 : _GEN_8806; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8808 = 9'h1b0 == _GEN_12982 ? phv_data_432 : _GEN_8807; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8809 = 9'h1b1 == _GEN_12982 ? phv_data_433 : _GEN_8808; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8810 = 9'h1b2 == _GEN_12982 ? phv_data_434 : _GEN_8809; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8811 = 9'h1b3 == _GEN_12982 ? phv_data_435 : _GEN_8810; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8812 = 9'h1b4 == _GEN_12982 ? phv_data_436 : _GEN_8811; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8813 = 9'h1b5 == _GEN_12982 ? phv_data_437 : _GEN_8812; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8814 = 9'h1b6 == _GEN_12982 ? phv_data_438 : _GEN_8813; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8815 = 9'h1b7 == _GEN_12982 ? phv_data_439 : _GEN_8814; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8816 = 9'h1b8 == _GEN_12982 ? phv_data_440 : _GEN_8815; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8817 = 9'h1b9 == _GEN_12982 ? phv_data_441 : _GEN_8816; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8818 = 9'h1ba == _GEN_12982 ? phv_data_442 : _GEN_8817; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8819 = 9'h1bb == _GEN_12982 ? phv_data_443 : _GEN_8818; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8820 = 9'h1bc == _GEN_12982 ? phv_data_444 : _GEN_8819; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8821 = 9'h1bd == _GEN_12982 ? phv_data_445 : _GEN_8820; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8822 = 9'h1be == _GEN_12982 ? phv_data_446 : _GEN_8821; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8823 = 9'h1bf == _GEN_12982 ? phv_data_447 : _GEN_8822; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8824 = 9'h1c0 == _GEN_12982 ? phv_data_448 : _GEN_8823; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8825 = 9'h1c1 == _GEN_12982 ? phv_data_449 : _GEN_8824; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8826 = 9'h1c2 == _GEN_12982 ? phv_data_450 : _GEN_8825; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8827 = 9'h1c3 == _GEN_12982 ? phv_data_451 : _GEN_8826; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8828 = 9'h1c4 == _GEN_12982 ? phv_data_452 : _GEN_8827; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8829 = 9'h1c5 == _GEN_12982 ? phv_data_453 : _GEN_8828; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8830 = 9'h1c6 == _GEN_12982 ? phv_data_454 : _GEN_8829; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8831 = 9'h1c7 == _GEN_12982 ? phv_data_455 : _GEN_8830; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8832 = 9'h1c8 == _GEN_12982 ? phv_data_456 : _GEN_8831; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8833 = 9'h1c9 == _GEN_12982 ? phv_data_457 : _GEN_8832; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8834 = 9'h1ca == _GEN_12982 ? phv_data_458 : _GEN_8833; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8835 = 9'h1cb == _GEN_12982 ? phv_data_459 : _GEN_8834; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8836 = 9'h1cc == _GEN_12982 ? phv_data_460 : _GEN_8835; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8837 = 9'h1cd == _GEN_12982 ? phv_data_461 : _GEN_8836; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8838 = 9'h1ce == _GEN_12982 ? phv_data_462 : _GEN_8837; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8839 = 9'h1cf == _GEN_12982 ? phv_data_463 : _GEN_8838; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8840 = 9'h1d0 == _GEN_12982 ? phv_data_464 : _GEN_8839; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8841 = 9'h1d1 == _GEN_12982 ? phv_data_465 : _GEN_8840; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8842 = 9'h1d2 == _GEN_12982 ? phv_data_466 : _GEN_8841; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8843 = 9'h1d3 == _GEN_12982 ? phv_data_467 : _GEN_8842; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8844 = 9'h1d4 == _GEN_12982 ? phv_data_468 : _GEN_8843; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8845 = 9'h1d5 == _GEN_12982 ? phv_data_469 : _GEN_8844; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8846 = 9'h1d6 == _GEN_12982 ? phv_data_470 : _GEN_8845; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8847 = 9'h1d7 == _GEN_12982 ? phv_data_471 : _GEN_8846; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8848 = 9'h1d8 == _GEN_12982 ? phv_data_472 : _GEN_8847; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8849 = 9'h1d9 == _GEN_12982 ? phv_data_473 : _GEN_8848; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8850 = 9'h1da == _GEN_12982 ? phv_data_474 : _GEN_8849; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8851 = 9'h1db == _GEN_12982 ? phv_data_475 : _GEN_8850; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8852 = 9'h1dc == _GEN_12982 ? phv_data_476 : _GEN_8851; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8853 = 9'h1dd == _GEN_12982 ? phv_data_477 : _GEN_8852; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8854 = 9'h1de == _GEN_12982 ? phv_data_478 : _GEN_8853; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8855 = 9'h1df == _GEN_12982 ? phv_data_479 : _GEN_8854; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8856 = 9'h1e0 == _GEN_12982 ? phv_data_480 : _GEN_8855; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8857 = 9'h1e1 == _GEN_12982 ? phv_data_481 : _GEN_8856; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8858 = 9'h1e2 == _GEN_12982 ? phv_data_482 : _GEN_8857; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8859 = 9'h1e3 == _GEN_12982 ? phv_data_483 : _GEN_8858; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8860 = 9'h1e4 == _GEN_12982 ? phv_data_484 : _GEN_8859; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8861 = 9'h1e5 == _GEN_12982 ? phv_data_485 : _GEN_8860; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8862 = 9'h1e6 == _GEN_12982 ? phv_data_486 : _GEN_8861; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8863 = 9'h1e7 == _GEN_12982 ? phv_data_487 : _GEN_8862; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8864 = 9'h1e8 == _GEN_12982 ? phv_data_488 : _GEN_8863; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8865 = 9'h1e9 == _GEN_12982 ? phv_data_489 : _GEN_8864; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8866 = 9'h1ea == _GEN_12982 ? phv_data_490 : _GEN_8865; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8867 = 9'h1eb == _GEN_12982 ? phv_data_491 : _GEN_8866; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8868 = 9'h1ec == _GEN_12982 ? phv_data_492 : _GEN_8867; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8869 = 9'h1ed == _GEN_12982 ? phv_data_493 : _GEN_8868; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8870 = 9'h1ee == _GEN_12982 ? phv_data_494 : _GEN_8869; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8871 = 9'h1ef == _GEN_12982 ? phv_data_495 : _GEN_8870; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8872 = 9'h1f0 == _GEN_12982 ? phv_data_496 : _GEN_8871; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8873 = 9'h1f1 == _GEN_12982 ? phv_data_497 : _GEN_8872; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8874 = 9'h1f2 == _GEN_12982 ? phv_data_498 : _GEN_8873; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8875 = 9'h1f3 == _GEN_12982 ? phv_data_499 : _GEN_8874; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8876 = 9'h1f4 == _GEN_12982 ? phv_data_500 : _GEN_8875; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8877 = 9'h1f5 == _GEN_12982 ? phv_data_501 : _GEN_8876; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8878 = 9'h1f6 == _GEN_12982 ? phv_data_502 : _GEN_8877; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8879 = 9'h1f7 == _GEN_12982 ? phv_data_503 : _GEN_8878; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8880 = 9'h1f8 == _GEN_12982 ? phv_data_504 : _GEN_8879; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8881 = 9'h1f9 == _GEN_12982 ? phv_data_505 : _GEN_8880; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8882 = 9'h1fa == _GEN_12982 ? phv_data_506 : _GEN_8881; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8883 = 9'h1fb == _GEN_12982 ? phv_data_507 : _GEN_8882; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8884 = 9'h1fc == _GEN_12982 ? phv_data_508 : _GEN_8883; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8885 = 9'h1fd == _GEN_12982 ? phv_data_509 : _GEN_8884; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] _GEN_8886 = 9'h1fe == _GEN_12982 ? phv_data_510 : _GEN_8885; // @[executor.scala 197:66 executor.scala 197:66]
  wire [7:0] bytes_3_0 = 9'h1ff == _GEN_12982 ? phv_data_511 : _GEN_8886; // @[executor.scala 197:66 executor.scala 197:66]
  wire [31:0] _io_field_out_3_T = {bytes_3_0,bytes_3_1,bytes_3_2,bytes_3_3}; // @[Cat.scala 30:58]
  wire [3:0] _io_mask_out_3_T = {_mask_3_T_24,mask_3_1,mask_3_2,mask_3_3}; // @[Cat.scala 30:58]
  wire [2:0] args_offset_3 = io_field_out_3_lo[13:11]; // @[primitive.scala 35:52]
  wire [2:0] args_length_3 = io_field_out_3_lo[10:8]; // @[primitive.scala 36:52]
  wire [3:0] _local_offset_T_169 = {{1'd0}, args_offset_3}; // @[executor.scala 222:61]
  wire [2:0] local_offset_84 = _local_offset_T_169[2:0]; // @[executor.scala 222:61]
  wire [7:0] _GEN_8889 = 3'h1 == local_offset_84 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8890 = 3'h2 == local_offset_84 ? args_2 : _GEN_8889; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8891 = 3'h3 == local_offset_84 ? args_3 : _GEN_8890; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8892 = 3'h4 == local_offset_84 ? args_4 : _GEN_8891; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8893 = 3'h5 == local_offset_84 ? args_5 : _GEN_8892; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8894 = 3'h6 == local_offset_84 ? args_6 : _GEN_8893; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8895 = 3'h1 == args_length_3 ? _GEN_8894 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [2:0] local_offset_85 = 3'h1 + args_offset_3; // @[executor.scala 222:61]
  wire [7:0] _GEN_8897 = 3'h1 == local_offset_85 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8898 = 3'h2 == local_offset_85 ? args_2 : _GEN_8897; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8899 = 3'h3 == local_offset_85 ? args_3 : _GEN_8898; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8900 = 3'h4 == local_offset_85 ? args_4 : _GEN_8899; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8901 = 3'h5 == local_offset_85 ? args_5 : _GEN_8900; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8902 = 3'h6 == local_offset_85 ? args_6 : _GEN_8901; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8903 = 3'h2 == args_length_3 ? _GEN_8902 : _GEN_8895; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_86 = 3'h2 + args_offset_3; // @[executor.scala 222:61]
  wire [7:0] _GEN_8905 = 3'h1 == local_offset_86 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8906 = 3'h2 == local_offset_86 ? args_2 : _GEN_8905; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8907 = 3'h3 == local_offset_86 ? args_3 : _GEN_8906; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8908 = 3'h4 == local_offset_86 ? args_4 : _GEN_8907; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8909 = 3'h5 == local_offset_86 ? args_5 : _GEN_8908; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8910 = 3'h6 == local_offset_86 ? args_6 : _GEN_8909; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8911 = 3'h3 == args_length_3 ? _GEN_8910 : _GEN_8903; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_87 = 3'h3 + args_offset_3; // @[executor.scala 222:61]
  wire [7:0] _GEN_8913 = 3'h1 == local_offset_87 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8914 = 3'h2 == local_offset_87 ? args_2 : _GEN_8913; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8915 = 3'h3 == local_offset_87 ? args_3 : _GEN_8914; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8916 = 3'h4 == local_offset_87 ? args_4 : _GEN_8915; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8917 = 3'h5 == local_offset_87 ? args_5 : _GEN_8916; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8918 = 3'h6 == local_offset_87 ? args_6 : _GEN_8917; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8919 = 3'h4 == args_length_3 ? _GEN_8918 : _GEN_8911; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_88 = 3'h4 + args_offset_3; // @[executor.scala 222:61]
  wire [7:0] _GEN_8921 = 3'h1 == local_offset_88 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8922 = 3'h2 == local_offset_88 ? args_2 : _GEN_8921; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8923 = 3'h3 == local_offset_88 ? args_3 : _GEN_8922; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8924 = 3'h4 == local_offset_88 ? args_4 : _GEN_8923; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8925 = 3'h5 == local_offset_88 ? args_5 : _GEN_8924; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8926 = 3'h6 == local_offset_88 ? args_6 : _GEN_8925; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8927 = 3'h5 == args_length_3 ? _GEN_8926 : _GEN_8919; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_89 = 3'h5 + args_offset_3; // @[executor.scala 222:61]
  wire [7:0] _GEN_8929 = 3'h1 == local_offset_89 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8930 = 3'h2 == local_offset_89 ? args_2 : _GEN_8929; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8931 = 3'h3 == local_offset_89 ? args_3 : _GEN_8930; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8932 = 3'h4 == local_offset_89 ? args_4 : _GEN_8931; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8933 = 3'h5 == local_offset_89 ? args_5 : _GEN_8932; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8934 = 3'h6 == local_offset_89 ? args_6 : _GEN_8933; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8935 = 3'h6 == args_length_3 ? _GEN_8934 : _GEN_8927; // @[executor.scala 223:66 executor.scala 224:52]
  wire [2:0] local_offset_90 = 3'h6 + args_offset_3; // @[executor.scala 222:61]
  wire [7:0] _GEN_8937 = 3'h1 == local_offset_90 ? args_1 : args_0; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8938 = 3'h2 == local_offset_90 ? args_2 : _GEN_8937; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8939 = 3'h3 == local_offset_90 ? args_3 : _GEN_8938; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8940 = 3'h4 == local_offset_90 ? args_4 : _GEN_8939; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8941 = 3'h5 == local_offset_90 ? args_5 : _GEN_8940; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] _GEN_8942 = 3'h6 == local_offset_90 ? args_6 : _GEN_8941; // @[executor.scala 224:52 executor.scala 224:52]
  wire [7:0] field_bytes_7_0 = 3'h7 == args_length_3 ? _GEN_8942 : _GEN_8935; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_8951 = 3'h2 == args_length_3 ? _GEN_8894 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_8959 = 3'h3 == args_length_3 ? _GEN_8902 : _GEN_8951; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_8967 = 3'h4 == args_length_3 ? _GEN_8910 : _GEN_8959; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_8975 = 3'h5 == args_length_3 ? _GEN_8918 : _GEN_8967; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_8983 = 3'h6 == args_length_3 ? _GEN_8926 : _GEN_8975; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_8991 = 3'h7 == args_length_3 ? _GEN_8934 : _GEN_8983; // @[executor.scala 223:66 executor.scala 224:52]
  wire [3:0] _GEN_13238 = {{1'd0}, args_length_3}; // @[executor.scala 223:49]
  wire [7:0] field_bytes_7_1 = 4'h8 == _GEN_13238 ? _GEN_8942 : _GEN_8991; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9007 = 3'h3 == args_length_3 ? _GEN_8894 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_9015 = 3'h4 == args_length_3 ? _GEN_8902 : _GEN_9007; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9023 = 3'h5 == args_length_3 ? _GEN_8910 : _GEN_9015; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9031 = 3'h6 == args_length_3 ? _GEN_8918 : _GEN_9023; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9039 = 3'h7 == args_length_3 ? _GEN_8926 : _GEN_9031; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9047 = 4'h8 == _GEN_13238 ? _GEN_8934 : _GEN_9039; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_7_2 = 4'h9 == _GEN_13238 ? _GEN_8942 : _GEN_9047; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9063 = 3'h4 == args_length_3 ? _GEN_8894 : 8'h0; // @[executor.scala 223:66 executor.scala 224:52 executor.scala 220:44]
  wire [7:0] _GEN_9071 = 3'h5 == args_length_3 ? _GEN_8902 : _GEN_9063; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9079 = 3'h6 == args_length_3 ? _GEN_8910 : _GEN_9071; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9087 = 3'h7 == args_length_3 ? _GEN_8918 : _GEN_9079; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9095 = 4'h8 == _GEN_13238 ? _GEN_8926 : _GEN_9087; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] _GEN_9103 = 4'h9 == _GEN_13238 ? _GEN_8934 : _GEN_9095; // @[executor.scala 223:66 executor.scala 224:52]
  wire [7:0] field_bytes_7_3 = 4'ha == _GEN_13238 ? _GEN_8942 : _GEN_9103; // @[executor.scala 223:66 executor.scala 224:52]
  wire [31:0] _io_field_out_3_T_1 = {field_bytes_7_0,field_bytes_7_1,field_bytes_7_2,field_bytes_7_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_9112 = 4'ha == opcode_3 ? _io_field_out_3_T_1 : 32'h0; // @[executor.scala 207:55 executor.scala 228:41 executor.scala 172:29]
  wire [17:0] io_field_out_3_hi_4 = io_field_out_3_lo[13] ? 18'h3ffff : 18'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _io_field_out_3_T_4 = {io_field_out_3_hi_4,io_field_out_3_lo}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_9113 = 4'hb == opcode_3 ? _io_field_out_3_T_4 : _GEN_9112; // @[executor.scala 230:56 executor.scala 231:41]
  wire [1:0] _GEN_9114 = from_header_3 ? bias_3 : 2'h0; // @[executor.scala 178:36 executor.scala 203:36 executor.scala 174:29]
  wire [31:0] _GEN_9115 = from_header_3 ? _io_field_out_3_T : _GEN_9113; // @[executor.scala 178:36 executor.scala 204:37]
  wire [3:0] _GEN_9116 = from_header_3 ? _io_mask_out_3_T : 4'h0; // @[executor.scala 178:36 executor.scala 205:37 executor.scala 173:29]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_256 = phv_data_256; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_257 = phv_data_257; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_258 = phv_data_258; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_259 = phv_data_259; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_260 = phv_data_260; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_261 = phv_data_261; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_262 = phv_data_262; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_263 = phv_data_263; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_264 = phv_data_264; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_265 = phv_data_265; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_266 = phv_data_266; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_267 = phv_data_267; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_268 = phv_data_268; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_269 = phv_data_269; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_270 = phv_data_270; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_271 = phv_data_271; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_272 = phv_data_272; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_273 = phv_data_273; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_274 = phv_data_274; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_275 = phv_data_275; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_276 = phv_data_276; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_277 = phv_data_277; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_278 = phv_data_278; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_279 = phv_data_279; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_280 = phv_data_280; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_281 = phv_data_281; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_282 = phv_data_282; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_283 = phv_data_283; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_284 = phv_data_284; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_285 = phv_data_285; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_286 = phv_data_286; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_287 = phv_data_287; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_288 = phv_data_288; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_289 = phv_data_289; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_290 = phv_data_290; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_291 = phv_data_291; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_292 = phv_data_292; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_293 = phv_data_293; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_294 = phv_data_294; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_295 = phv_data_295; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_296 = phv_data_296; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_297 = phv_data_297; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_298 = phv_data_298; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_299 = phv_data_299; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_300 = phv_data_300; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_301 = phv_data_301; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_302 = phv_data_302; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_303 = phv_data_303; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_304 = phv_data_304; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_305 = phv_data_305; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_306 = phv_data_306; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_307 = phv_data_307; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_308 = phv_data_308; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_309 = phv_data_309; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_310 = phv_data_310; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_311 = phv_data_311; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_312 = phv_data_312; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_313 = phv_data_313; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_314 = phv_data_314; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_315 = phv_data_315; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_316 = phv_data_316; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_317 = phv_data_317; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_318 = phv_data_318; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_319 = phv_data_319; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_320 = phv_data_320; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_321 = phv_data_321; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_322 = phv_data_322; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_323 = phv_data_323; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_324 = phv_data_324; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_325 = phv_data_325; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_326 = phv_data_326; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_327 = phv_data_327; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_328 = phv_data_328; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_329 = phv_data_329; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_330 = phv_data_330; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_331 = phv_data_331; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_332 = phv_data_332; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_333 = phv_data_333; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_334 = phv_data_334; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_335 = phv_data_335; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_336 = phv_data_336; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_337 = phv_data_337; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_338 = phv_data_338; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_339 = phv_data_339; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_340 = phv_data_340; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_341 = phv_data_341; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_342 = phv_data_342; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_343 = phv_data_343; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_344 = phv_data_344; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_345 = phv_data_345; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_346 = phv_data_346; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_347 = phv_data_347; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_348 = phv_data_348; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_349 = phv_data_349; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_350 = phv_data_350; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_351 = phv_data_351; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_352 = phv_data_352; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_353 = phv_data_353; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_354 = phv_data_354; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_355 = phv_data_355; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_356 = phv_data_356; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_357 = phv_data_357; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_358 = phv_data_358; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_359 = phv_data_359; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_360 = phv_data_360; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_361 = phv_data_361; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_362 = phv_data_362; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_363 = phv_data_363; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_364 = phv_data_364; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_365 = phv_data_365; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_366 = phv_data_366; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_367 = phv_data_367; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_368 = phv_data_368; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_369 = phv_data_369; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_370 = phv_data_370; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_371 = phv_data_371; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_372 = phv_data_372; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_373 = phv_data_373; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_374 = phv_data_374; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_375 = phv_data_375; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_376 = phv_data_376; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_377 = phv_data_377; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_378 = phv_data_378; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_379 = phv_data_379; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_380 = phv_data_380; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_381 = phv_data_381; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_382 = phv_data_382; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_383 = phv_data_383; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_384 = phv_data_384; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_385 = phv_data_385; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_386 = phv_data_386; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_387 = phv_data_387; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_388 = phv_data_388; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_389 = phv_data_389; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_390 = phv_data_390; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_391 = phv_data_391; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_392 = phv_data_392; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_393 = phv_data_393; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_394 = phv_data_394; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_395 = phv_data_395; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_396 = phv_data_396; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_397 = phv_data_397; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_398 = phv_data_398; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_399 = phv_data_399; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_400 = phv_data_400; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_401 = phv_data_401; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_402 = phv_data_402; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_403 = phv_data_403; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_404 = phv_data_404; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_405 = phv_data_405; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_406 = phv_data_406; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_407 = phv_data_407; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_408 = phv_data_408; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_409 = phv_data_409; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_410 = phv_data_410; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_411 = phv_data_411; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_412 = phv_data_412; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_413 = phv_data_413; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_414 = phv_data_414; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_415 = phv_data_415; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_416 = phv_data_416; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_417 = phv_data_417; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_418 = phv_data_418; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_419 = phv_data_419; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_420 = phv_data_420; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_421 = phv_data_421; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_422 = phv_data_422; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_423 = phv_data_423; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_424 = phv_data_424; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_425 = phv_data_425; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_426 = phv_data_426; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_427 = phv_data_427; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_428 = phv_data_428; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_429 = phv_data_429; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_430 = phv_data_430; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_431 = phv_data_431; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_432 = phv_data_432; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_433 = phv_data_433; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_434 = phv_data_434; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_435 = phv_data_435; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_436 = phv_data_436; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_437 = phv_data_437; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_438 = phv_data_438; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_439 = phv_data_439; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_440 = phv_data_440; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_441 = phv_data_441; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_442 = phv_data_442; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_443 = phv_data_443; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_444 = phv_data_444; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_445 = phv_data_445; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_446 = phv_data_446; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_447 = phv_data_447; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_448 = phv_data_448; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_449 = phv_data_449; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_450 = phv_data_450; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_451 = phv_data_451; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_452 = phv_data_452; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_453 = phv_data_453; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_454 = phv_data_454; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_455 = phv_data_455; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_456 = phv_data_456; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_457 = phv_data_457; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_458 = phv_data_458; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_459 = phv_data_459; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_460 = phv_data_460; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_461 = phv_data_461; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_462 = phv_data_462; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_463 = phv_data_463; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_464 = phv_data_464; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_465 = phv_data_465; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_466 = phv_data_466; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_467 = phv_data_467; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_468 = phv_data_468; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_469 = phv_data_469; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_470 = phv_data_470; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_471 = phv_data_471; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_472 = phv_data_472; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_473 = phv_data_473; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_474 = phv_data_474; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_475 = phv_data_475; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_476 = phv_data_476; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_477 = phv_data_477; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_478 = phv_data_478; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_479 = phv_data_479; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_480 = phv_data_480; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_481 = phv_data_481; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_482 = phv_data_482; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_483 = phv_data_483; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_484 = phv_data_484; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_485 = phv_data_485; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_486 = phv_data_486; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_487 = phv_data_487; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_488 = phv_data_488; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_489 = phv_data_489; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_490 = phv_data_490; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_491 = phv_data_491; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_492 = phv_data_492; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_493 = phv_data_493; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_494 = phv_data_494; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_495 = phv_data_495; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_496 = phv_data_496; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_497 = phv_data_497; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_498 = phv_data_498; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_499 = phv_data_499; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_500 = phv_data_500; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_501 = phv_data_501; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_502 = phv_data_502; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_503 = phv_data_503; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_504 = phv_data_504; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_505 = phv_data_505; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_506 = phv_data_506; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_507 = phv_data_507; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_508 = phv_data_508; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_509 = phv_data_509; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_510 = phv_data_510; // @[executor.scala 153:25]
  assign io_pipe_phv_out_data_511 = phv_data_511; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[executor.scala 153:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[executor.scala 153:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[executor.scala 153:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[executor.scala 153:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[executor.scala 153:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor.scala 153:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[executor.scala 153:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[executor.scala 153:25]
  assign io_vliw_out_0 = vliw_0; // @[executor.scala 160:21]
  assign io_vliw_out_1 = vliw_1; // @[executor.scala 160:21]
  assign io_vliw_out_2 = vliw_2; // @[executor.scala 160:21]
  assign io_vliw_out_3 = vliw_3; // @[executor.scala 160:21]
  assign io_field_out_0 = phv_is_valid_processor ? _GEN_2275 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_field_out_1 = phv_is_valid_processor ? _GEN_4555 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_field_out_2 = phv_is_valid_processor ? _GEN_6835 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_field_out_3 = phv_is_valid_processor ? _GEN_9115 : 32'h0; // @[executor.scala 176:43 executor.scala 172:29]
  assign io_mask_out_0 = phv_is_valid_processor ? _GEN_2276 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_mask_out_1 = phv_is_valid_processor ? _GEN_4556 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_mask_out_2 = phv_is_valid_processor ? _GEN_6836 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_mask_out_3 = phv_is_valid_processor ? _GEN_9116 : 4'h0; // @[executor.scala 176:43 executor.scala 173:29]
  assign io_bias_out_0 = phv_is_valid_processor ? _GEN_2274 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  assign io_bias_out_1 = phv_is_valid_processor ? _GEN_4554 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  assign io_bias_out_2 = phv_is_valid_processor ? _GEN_6834 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  assign io_bias_out_3 = phv_is_valid_processor ? _GEN_9114 : 2'h0; // @[executor.scala 176:43 executor.scala 174:29]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor.scala 152:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor.scala 152:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor.scala 152:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor.scala 152:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor.scala 152:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor.scala 152:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor.scala 152:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor.scala 152:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor.scala 152:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor.scala 152:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor.scala 152:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor.scala 152:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor.scala 152:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor.scala 152:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor.scala 152:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor.scala 152:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor.scala 152:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor.scala 152:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor.scala 152:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor.scala 152:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor.scala 152:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor.scala 152:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor.scala 152:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor.scala 152:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor.scala 152:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor.scala 152:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor.scala 152:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor.scala 152:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor.scala 152:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor.scala 152:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor.scala 152:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor.scala 152:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor.scala 152:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor.scala 152:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor.scala 152:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor.scala 152:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor.scala 152:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor.scala 152:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor.scala 152:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor.scala 152:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor.scala 152:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor.scala 152:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor.scala 152:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor.scala 152:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor.scala 152:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor.scala 152:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor.scala 152:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor.scala 152:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor.scala 152:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor.scala 152:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor.scala 152:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor.scala 152:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor.scala 152:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor.scala 152:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor.scala 152:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor.scala 152:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor.scala 152:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor.scala 152:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor.scala 152:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor.scala 152:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor.scala 152:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor.scala 152:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor.scala 152:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor.scala 152:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor.scala 152:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor.scala 152:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor.scala 152:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor.scala 152:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor.scala 152:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor.scala 152:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor.scala 152:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor.scala 152:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor.scala 152:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor.scala 152:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor.scala 152:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor.scala 152:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor.scala 152:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor.scala 152:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor.scala 152:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor.scala 152:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor.scala 152:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor.scala 152:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor.scala 152:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor.scala 152:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor.scala 152:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor.scala 152:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor.scala 152:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor.scala 152:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor.scala 152:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor.scala 152:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor.scala 152:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor.scala 152:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor.scala 152:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor.scala 152:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor.scala 152:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor.scala 152:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor.scala 152:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor.scala 152:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor.scala 152:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor.scala 152:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor.scala 152:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor.scala 152:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor.scala 152:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor.scala 152:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor.scala 152:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor.scala 152:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor.scala 152:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor.scala 152:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor.scala 152:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor.scala 152:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor.scala 152:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor.scala 152:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor.scala 152:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor.scala 152:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor.scala 152:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor.scala 152:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor.scala 152:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor.scala 152:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor.scala 152:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor.scala 152:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor.scala 152:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor.scala 152:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor.scala 152:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor.scala 152:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor.scala 152:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor.scala 152:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor.scala 152:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor.scala 152:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor.scala 152:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor.scala 152:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor.scala 152:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor.scala 152:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor.scala 152:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor.scala 152:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor.scala 152:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor.scala 152:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor.scala 152:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor.scala 152:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor.scala 152:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor.scala 152:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor.scala 152:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor.scala 152:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor.scala 152:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor.scala 152:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor.scala 152:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor.scala 152:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor.scala 152:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor.scala 152:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor.scala 152:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor.scala 152:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor.scala 152:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor.scala 152:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor.scala 152:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor.scala 152:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor.scala 152:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor.scala 152:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor.scala 152:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor.scala 152:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor.scala 152:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor.scala 152:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor.scala 152:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor.scala 152:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor.scala 152:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor.scala 152:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor.scala 152:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor.scala 152:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor.scala 152:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor.scala 152:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor.scala 152:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor.scala 152:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor.scala 152:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor.scala 152:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor.scala 152:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor.scala 152:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor.scala 152:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor.scala 152:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor.scala 152:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor.scala 152:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor.scala 152:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor.scala 152:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor.scala 152:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor.scala 152:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor.scala 152:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor.scala 152:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor.scala 152:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor.scala 152:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor.scala 152:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor.scala 152:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor.scala 152:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor.scala 152:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor.scala 152:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor.scala 152:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor.scala 152:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor.scala 152:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor.scala 152:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor.scala 152:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor.scala 152:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor.scala 152:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor.scala 152:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor.scala 152:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor.scala 152:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor.scala 152:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor.scala 152:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor.scala 152:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor.scala 152:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor.scala 152:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor.scala 152:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor.scala 152:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor.scala 152:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor.scala 152:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor.scala 152:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor.scala 152:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor.scala 152:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor.scala 152:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor.scala 152:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor.scala 152:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor.scala 152:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor.scala 152:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor.scala 152:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor.scala 152:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor.scala 152:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor.scala 152:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor.scala 152:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor.scala 152:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor.scala 152:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor.scala 152:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor.scala 152:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor.scala 152:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor.scala 152:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor.scala 152:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor.scala 152:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor.scala 152:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor.scala 152:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor.scala 152:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor.scala 152:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor.scala 152:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor.scala 152:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor.scala 152:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor.scala 152:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor.scala 152:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor.scala 152:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor.scala 152:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor.scala 152:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor.scala 152:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor.scala 152:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor.scala 152:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor.scala 152:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor.scala 152:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor.scala 152:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor.scala 152:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor.scala 152:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor.scala 152:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor.scala 152:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor.scala 152:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor.scala 152:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor.scala 152:13]
    phv_data_256 <= io_pipe_phv_in_data_256; // @[executor.scala 152:13]
    phv_data_257 <= io_pipe_phv_in_data_257; // @[executor.scala 152:13]
    phv_data_258 <= io_pipe_phv_in_data_258; // @[executor.scala 152:13]
    phv_data_259 <= io_pipe_phv_in_data_259; // @[executor.scala 152:13]
    phv_data_260 <= io_pipe_phv_in_data_260; // @[executor.scala 152:13]
    phv_data_261 <= io_pipe_phv_in_data_261; // @[executor.scala 152:13]
    phv_data_262 <= io_pipe_phv_in_data_262; // @[executor.scala 152:13]
    phv_data_263 <= io_pipe_phv_in_data_263; // @[executor.scala 152:13]
    phv_data_264 <= io_pipe_phv_in_data_264; // @[executor.scala 152:13]
    phv_data_265 <= io_pipe_phv_in_data_265; // @[executor.scala 152:13]
    phv_data_266 <= io_pipe_phv_in_data_266; // @[executor.scala 152:13]
    phv_data_267 <= io_pipe_phv_in_data_267; // @[executor.scala 152:13]
    phv_data_268 <= io_pipe_phv_in_data_268; // @[executor.scala 152:13]
    phv_data_269 <= io_pipe_phv_in_data_269; // @[executor.scala 152:13]
    phv_data_270 <= io_pipe_phv_in_data_270; // @[executor.scala 152:13]
    phv_data_271 <= io_pipe_phv_in_data_271; // @[executor.scala 152:13]
    phv_data_272 <= io_pipe_phv_in_data_272; // @[executor.scala 152:13]
    phv_data_273 <= io_pipe_phv_in_data_273; // @[executor.scala 152:13]
    phv_data_274 <= io_pipe_phv_in_data_274; // @[executor.scala 152:13]
    phv_data_275 <= io_pipe_phv_in_data_275; // @[executor.scala 152:13]
    phv_data_276 <= io_pipe_phv_in_data_276; // @[executor.scala 152:13]
    phv_data_277 <= io_pipe_phv_in_data_277; // @[executor.scala 152:13]
    phv_data_278 <= io_pipe_phv_in_data_278; // @[executor.scala 152:13]
    phv_data_279 <= io_pipe_phv_in_data_279; // @[executor.scala 152:13]
    phv_data_280 <= io_pipe_phv_in_data_280; // @[executor.scala 152:13]
    phv_data_281 <= io_pipe_phv_in_data_281; // @[executor.scala 152:13]
    phv_data_282 <= io_pipe_phv_in_data_282; // @[executor.scala 152:13]
    phv_data_283 <= io_pipe_phv_in_data_283; // @[executor.scala 152:13]
    phv_data_284 <= io_pipe_phv_in_data_284; // @[executor.scala 152:13]
    phv_data_285 <= io_pipe_phv_in_data_285; // @[executor.scala 152:13]
    phv_data_286 <= io_pipe_phv_in_data_286; // @[executor.scala 152:13]
    phv_data_287 <= io_pipe_phv_in_data_287; // @[executor.scala 152:13]
    phv_data_288 <= io_pipe_phv_in_data_288; // @[executor.scala 152:13]
    phv_data_289 <= io_pipe_phv_in_data_289; // @[executor.scala 152:13]
    phv_data_290 <= io_pipe_phv_in_data_290; // @[executor.scala 152:13]
    phv_data_291 <= io_pipe_phv_in_data_291; // @[executor.scala 152:13]
    phv_data_292 <= io_pipe_phv_in_data_292; // @[executor.scala 152:13]
    phv_data_293 <= io_pipe_phv_in_data_293; // @[executor.scala 152:13]
    phv_data_294 <= io_pipe_phv_in_data_294; // @[executor.scala 152:13]
    phv_data_295 <= io_pipe_phv_in_data_295; // @[executor.scala 152:13]
    phv_data_296 <= io_pipe_phv_in_data_296; // @[executor.scala 152:13]
    phv_data_297 <= io_pipe_phv_in_data_297; // @[executor.scala 152:13]
    phv_data_298 <= io_pipe_phv_in_data_298; // @[executor.scala 152:13]
    phv_data_299 <= io_pipe_phv_in_data_299; // @[executor.scala 152:13]
    phv_data_300 <= io_pipe_phv_in_data_300; // @[executor.scala 152:13]
    phv_data_301 <= io_pipe_phv_in_data_301; // @[executor.scala 152:13]
    phv_data_302 <= io_pipe_phv_in_data_302; // @[executor.scala 152:13]
    phv_data_303 <= io_pipe_phv_in_data_303; // @[executor.scala 152:13]
    phv_data_304 <= io_pipe_phv_in_data_304; // @[executor.scala 152:13]
    phv_data_305 <= io_pipe_phv_in_data_305; // @[executor.scala 152:13]
    phv_data_306 <= io_pipe_phv_in_data_306; // @[executor.scala 152:13]
    phv_data_307 <= io_pipe_phv_in_data_307; // @[executor.scala 152:13]
    phv_data_308 <= io_pipe_phv_in_data_308; // @[executor.scala 152:13]
    phv_data_309 <= io_pipe_phv_in_data_309; // @[executor.scala 152:13]
    phv_data_310 <= io_pipe_phv_in_data_310; // @[executor.scala 152:13]
    phv_data_311 <= io_pipe_phv_in_data_311; // @[executor.scala 152:13]
    phv_data_312 <= io_pipe_phv_in_data_312; // @[executor.scala 152:13]
    phv_data_313 <= io_pipe_phv_in_data_313; // @[executor.scala 152:13]
    phv_data_314 <= io_pipe_phv_in_data_314; // @[executor.scala 152:13]
    phv_data_315 <= io_pipe_phv_in_data_315; // @[executor.scala 152:13]
    phv_data_316 <= io_pipe_phv_in_data_316; // @[executor.scala 152:13]
    phv_data_317 <= io_pipe_phv_in_data_317; // @[executor.scala 152:13]
    phv_data_318 <= io_pipe_phv_in_data_318; // @[executor.scala 152:13]
    phv_data_319 <= io_pipe_phv_in_data_319; // @[executor.scala 152:13]
    phv_data_320 <= io_pipe_phv_in_data_320; // @[executor.scala 152:13]
    phv_data_321 <= io_pipe_phv_in_data_321; // @[executor.scala 152:13]
    phv_data_322 <= io_pipe_phv_in_data_322; // @[executor.scala 152:13]
    phv_data_323 <= io_pipe_phv_in_data_323; // @[executor.scala 152:13]
    phv_data_324 <= io_pipe_phv_in_data_324; // @[executor.scala 152:13]
    phv_data_325 <= io_pipe_phv_in_data_325; // @[executor.scala 152:13]
    phv_data_326 <= io_pipe_phv_in_data_326; // @[executor.scala 152:13]
    phv_data_327 <= io_pipe_phv_in_data_327; // @[executor.scala 152:13]
    phv_data_328 <= io_pipe_phv_in_data_328; // @[executor.scala 152:13]
    phv_data_329 <= io_pipe_phv_in_data_329; // @[executor.scala 152:13]
    phv_data_330 <= io_pipe_phv_in_data_330; // @[executor.scala 152:13]
    phv_data_331 <= io_pipe_phv_in_data_331; // @[executor.scala 152:13]
    phv_data_332 <= io_pipe_phv_in_data_332; // @[executor.scala 152:13]
    phv_data_333 <= io_pipe_phv_in_data_333; // @[executor.scala 152:13]
    phv_data_334 <= io_pipe_phv_in_data_334; // @[executor.scala 152:13]
    phv_data_335 <= io_pipe_phv_in_data_335; // @[executor.scala 152:13]
    phv_data_336 <= io_pipe_phv_in_data_336; // @[executor.scala 152:13]
    phv_data_337 <= io_pipe_phv_in_data_337; // @[executor.scala 152:13]
    phv_data_338 <= io_pipe_phv_in_data_338; // @[executor.scala 152:13]
    phv_data_339 <= io_pipe_phv_in_data_339; // @[executor.scala 152:13]
    phv_data_340 <= io_pipe_phv_in_data_340; // @[executor.scala 152:13]
    phv_data_341 <= io_pipe_phv_in_data_341; // @[executor.scala 152:13]
    phv_data_342 <= io_pipe_phv_in_data_342; // @[executor.scala 152:13]
    phv_data_343 <= io_pipe_phv_in_data_343; // @[executor.scala 152:13]
    phv_data_344 <= io_pipe_phv_in_data_344; // @[executor.scala 152:13]
    phv_data_345 <= io_pipe_phv_in_data_345; // @[executor.scala 152:13]
    phv_data_346 <= io_pipe_phv_in_data_346; // @[executor.scala 152:13]
    phv_data_347 <= io_pipe_phv_in_data_347; // @[executor.scala 152:13]
    phv_data_348 <= io_pipe_phv_in_data_348; // @[executor.scala 152:13]
    phv_data_349 <= io_pipe_phv_in_data_349; // @[executor.scala 152:13]
    phv_data_350 <= io_pipe_phv_in_data_350; // @[executor.scala 152:13]
    phv_data_351 <= io_pipe_phv_in_data_351; // @[executor.scala 152:13]
    phv_data_352 <= io_pipe_phv_in_data_352; // @[executor.scala 152:13]
    phv_data_353 <= io_pipe_phv_in_data_353; // @[executor.scala 152:13]
    phv_data_354 <= io_pipe_phv_in_data_354; // @[executor.scala 152:13]
    phv_data_355 <= io_pipe_phv_in_data_355; // @[executor.scala 152:13]
    phv_data_356 <= io_pipe_phv_in_data_356; // @[executor.scala 152:13]
    phv_data_357 <= io_pipe_phv_in_data_357; // @[executor.scala 152:13]
    phv_data_358 <= io_pipe_phv_in_data_358; // @[executor.scala 152:13]
    phv_data_359 <= io_pipe_phv_in_data_359; // @[executor.scala 152:13]
    phv_data_360 <= io_pipe_phv_in_data_360; // @[executor.scala 152:13]
    phv_data_361 <= io_pipe_phv_in_data_361; // @[executor.scala 152:13]
    phv_data_362 <= io_pipe_phv_in_data_362; // @[executor.scala 152:13]
    phv_data_363 <= io_pipe_phv_in_data_363; // @[executor.scala 152:13]
    phv_data_364 <= io_pipe_phv_in_data_364; // @[executor.scala 152:13]
    phv_data_365 <= io_pipe_phv_in_data_365; // @[executor.scala 152:13]
    phv_data_366 <= io_pipe_phv_in_data_366; // @[executor.scala 152:13]
    phv_data_367 <= io_pipe_phv_in_data_367; // @[executor.scala 152:13]
    phv_data_368 <= io_pipe_phv_in_data_368; // @[executor.scala 152:13]
    phv_data_369 <= io_pipe_phv_in_data_369; // @[executor.scala 152:13]
    phv_data_370 <= io_pipe_phv_in_data_370; // @[executor.scala 152:13]
    phv_data_371 <= io_pipe_phv_in_data_371; // @[executor.scala 152:13]
    phv_data_372 <= io_pipe_phv_in_data_372; // @[executor.scala 152:13]
    phv_data_373 <= io_pipe_phv_in_data_373; // @[executor.scala 152:13]
    phv_data_374 <= io_pipe_phv_in_data_374; // @[executor.scala 152:13]
    phv_data_375 <= io_pipe_phv_in_data_375; // @[executor.scala 152:13]
    phv_data_376 <= io_pipe_phv_in_data_376; // @[executor.scala 152:13]
    phv_data_377 <= io_pipe_phv_in_data_377; // @[executor.scala 152:13]
    phv_data_378 <= io_pipe_phv_in_data_378; // @[executor.scala 152:13]
    phv_data_379 <= io_pipe_phv_in_data_379; // @[executor.scala 152:13]
    phv_data_380 <= io_pipe_phv_in_data_380; // @[executor.scala 152:13]
    phv_data_381 <= io_pipe_phv_in_data_381; // @[executor.scala 152:13]
    phv_data_382 <= io_pipe_phv_in_data_382; // @[executor.scala 152:13]
    phv_data_383 <= io_pipe_phv_in_data_383; // @[executor.scala 152:13]
    phv_data_384 <= io_pipe_phv_in_data_384; // @[executor.scala 152:13]
    phv_data_385 <= io_pipe_phv_in_data_385; // @[executor.scala 152:13]
    phv_data_386 <= io_pipe_phv_in_data_386; // @[executor.scala 152:13]
    phv_data_387 <= io_pipe_phv_in_data_387; // @[executor.scala 152:13]
    phv_data_388 <= io_pipe_phv_in_data_388; // @[executor.scala 152:13]
    phv_data_389 <= io_pipe_phv_in_data_389; // @[executor.scala 152:13]
    phv_data_390 <= io_pipe_phv_in_data_390; // @[executor.scala 152:13]
    phv_data_391 <= io_pipe_phv_in_data_391; // @[executor.scala 152:13]
    phv_data_392 <= io_pipe_phv_in_data_392; // @[executor.scala 152:13]
    phv_data_393 <= io_pipe_phv_in_data_393; // @[executor.scala 152:13]
    phv_data_394 <= io_pipe_phv_in_data_394; // @[executor.scala 152:13]
    phv_data_395 <= io_pipe_phv_in_data_395; // @[executor.scala 152:13]
    phv_data_396 <= io_pipe_phv_in_data_396; // @[executor.scala 152:13]
    phv_data_397 <= io_pipe_phv_in_data_397; // @[executor.scala 152:13]
    phv_data_398 <= io_pipe_phv_in_data_398; // @[executor.scala 152:13]
    phv_data_399 <= io_pipe_phv_in_data_399; // @[executor.scala 152:13]
    phv_data_400 <= io_pipe_phv_in_data_400; // @[executor.scala 152:13]
    phv_data_401 <= io_pipe_phv_in_data_401; // @[executor.scala 152:13]
    phv_data_402 <= io_pipe_phv_in_data_402; // @[executor.scala 152:13]
    phv_data_403 <= io_pipe_phv_in_data_403; // @[executor.scala 152:13]
    phv_data_404 <= io_pipe_phv_in_data_404; // @[executor.scala 152:13]
    phv_data_405 <= io_pipe_phv_in_data_405; // @[executor.scala 152:13]
    phv_data_406 <= io_pipe_phv_in_data_406; // @[executor.scala 152:13]
    phv_data_407 <= io_pipe_phv_in_data_407; // @[executor.scala 152:13]
    phv_data_408 <= io_pipe_phv_in_data_408; // @[executor.scala 152:13]
    phv_data_409 <= io_pipe_phv_in_data_409; // @[executor.scala 152:13]
    phv_data_410 <= io_pipe_phv_in_data_410; // @[executor.scala 152:13]
    phv_data_411 <= io_pipe_phv_in_data_411; // @[executor.scala 152:13]
    phv_data_412 <= io_pipe_phv_in_data_412; // @[executor.scala 152:13]
    phv_data_413 <= io_pipe_phv_in_data_413; // @[executor.scala 152:13]
    phv_data_414 <= io_pipe_phv_in_data_414; // @[executor.scala 152:13]
    phv_data_415 <= io_pipe_phv_in_data_415; // @[executor.scala 152:13]
    phv_data_416 <= io_pipe_phv_in_data_416; // @[executor.scala 152:13]
    phv_data_417 <= io_pipe_phv_in_data_417; // @[executor.scala 152:13]
    phv_data_418 <= io_pipe_phv_in_data_418; // @[executor.scala 152:13]
    phv_data_419 <= io_pipe_phv_in_data_419; // @[executor.scala 152:13]
    phv_data_420 <= io_pipe_phv_in_data_420; // @[executor.scala 152:13]
    phv_data_421 <= io_pipe_phv_in_data_421; // @[executor.scala 152:13]
    phv_data_422 <= io_pipe_phv_in_data_422; // @[executor.scala 152:13]
    phv_data_423 <= io_pipe_phv_in_data_423; // @[executor.scala 152:13]
    phv_data_424 <= io_pipe_phv_in_data_424; // @[executor.scala 152:13]
    phv_data_425 <= io_pipe_phv_in_data_425; // @[executor.scala 152:13]
    phv_data_426 <= io_pipe_phv_in_data_426; // @[executor.scala 152:13]
    phv_data_427 <= io_pipe_phv_in_data_427; // @[executor.scala 152:13]
    phv_data_428 <= io_pipe_phv_in_data_428; // @[executor.scala 152:13]
    phv_data_429 <= io_pipe_phv_in_data_429; // @[executor.scala 152:13]
    phv_data_430 <= io_pipe_phv_in_data_430; // @[executor.scala 152:13]
    phv_data_431 <= io_pipe_phv_in_data_431; // @[executor.scala 152:13]
    phv_data_432 <= io_pipe_phv_in_data_432; // @[executor.scala 152:13]
    phv_data_433 <= io_pipe_phv_in_data_433; // @[executor.scala 152:13]
    phv_data_434 <= io_pipe_phv_in_data_434; // @[executor.scala 152:13]
    phv_data_435 <= io_pipe_phv_in_data_435; // @[executor.scala 152:13]
    phv_data_436 <= io_pipe_phv_in_data_436; // @[executor.scala 152:13]
    phv_data_437 <= io_pipe_phv_in_data_437; // @[executor.scala 152:13]
    phv_data_438 <= io_pipe_phv_in_data_438; // @[executor.scala 152:13]
    phv_data_439 <= io_pipe_phv_in_data_439; // @[executor.scala 152:13]
    phv_data_440 <= io_pipe_phv_in_data_440; // @[executor.scala 152:13]
    phv_data_441 <= io_pipe_phv_in_data_441; // @[executor.scala 152:13]
    phv_data_442 <= io_pipe_phv_in_data_442; // @[executor.scala 152:13]
    phv_data_443 <= io_pipe_phv_in_data_443; // @[executor.scala 152:13]
    phv_data_444 <= io_pipe_phv_in_data_444; // @[executor.scala 152:13]
    phv_data_445 <= io_pipe_phv_in_data_445; // @[executor.scala 152:13]
    phv_data_446 <= io_pipe_phv_in_data_446; // @[executor.scala 152:13]
    phv_data_447 <= io_pipe_phv_in_data_447; // @[executor.scala 152:13]
    phv_data_448 <= io_pipe_phv_in_data_448; // @[executor.scala 152:13]
    phv_data_449 <= io_pipe_phv_in_data_449; // @[executor.scala 152:13]
    phv_data_450 <= io_pipe_phv_in_data_450; // @[executor.scala 152:13]
    phv_data_451 <= io_pipe_phv_in_data_451; // @[executor.scala 152:13]
    phv_data_452 <= io_pipe_phv_in_data_452; // @[executor.scala 152:13]
    phv_data_453 <= io_pipe_phv_in_data_453; // @[executor.scala 152:13]
    phv_data_454 <= io_pipe_phv_in_data_454; // @[executor.scala 152:13]
    phv_data_455 <= io_pipe_phv_in_data_455; // @[executor.scala 152:13]
    phv_data_456 <= io_pipe_phv_in_data_456; // @[executor.scala 152:13]
    phv_data_457 <= io_pipe_phv_in_data_457; // @[executor.scala 152:13]
    phv_data_458 <= io_pipe_phv_in_data_458; // @[executor.scala 152:13]
    phv_data_459 <= io_pipe_phv_in_data_459; // @[executor.scala 152:13]
    phv_data_460 <= io_pipe_phv_in_data_460; // @[executor.scala 152:13]
    phv_data_461 <= io_pipe_phv_in_data_461; // @[executor.scala 152:13]
    phv_data_462 <= io_pipe_phv_in_data_462; // @[executor.scala 152:13]
    phv_data_463 <= io_pipe_phv_in_data_463; // @[executor.scala 152:13]
    phv_data_464 <= io_pipe_phv_in_data_464; // @[executor.scala 152:13]
    phv_data_465 <= io_pipe_phv_in_data_465; // @[executor.scala 152:13]
    phv_data_466 <= io_pipe_phv_in_data_466; // @[executor.scala 152:13]
    phv_data_467 <= io_pipe_phv_in_data_467; // @[executor.scala 152:13]
    phv_data_468 <= io_pipe_phv_in_data_468; // @[executor.scala 152:13]
    phv_data_469 <= io_pipe_phv_in_data_469; // @[executor.scala 152:13]
    phv_data_470 <= io_pipe_phv_in_data_470; // @[executor.scala 152:13]
    phv_data_471 <= io_pipe_phv_in_data_471; // @[executor.scala 152:13]
    phv_data_472 <= io_pipe_phv_in_data_472; // @[executor.scala 152:13]
    phv_data_473 <= io_pipe_phv_in_data_473; // @[executor.scala 152:13]
    phv_data_474 <= io_pipe_phv_in_data_474; // @[executor.scala 152:13]
    phv_data_475 <= io_pipe_phv_in_data_475; // @[executor.scala 152:13]
    phv_data_476 <= io_pipe_phv_in_data_476; // @[executor.scala 152:13]
    phv_data_477 <= io_pipe_phv_in_data_477; // @[executor.scala 152:13]
    phv_data_478 <= io_pipe_phv_in_data_478; // @[executor.scala 152:13]
    phv_data_479 <= io_pipe_phv_in_data_479; // @[executor.scala 152:13]
    phv_data_480 <= io_pipe_phv_in_data_480; // @[executor.scala 152:13]
    phv_data_481 <= io_pipe_phv_in_data_481; // @[executor.scala 152:13]
    phv_data_482 <= io_pipe_phv_in_data_482; // @[executor.scala 152:13]
    phv_data_483 <= io_pipe_phv_in_data_483; // @[executor.scala 152:13]
    phv_data_484 <= io_pipe_phv_in_data_484; // @[executor.scala 152:13]
    phv_data_485 <= io_pipe_phv_in_data_485; // @[executor.scala 152:13]
    phv_data_486 <= io_pipe_phv_in_data_486; // @[executor.scala 152:13]
    phv_data_487 <= io_pipe_phv_in_data_487; // @[executor.scala 152:13]
    phv_data_488 <= io_pipe_phv_in_data_488; // @[executor.scala 152:13]
    phv_data_489 <= io_pipe_phv_in_data_489; // @[executor.scala 152:13]
    phv_data_490 <= io_pipe_phv_in_data_490; // @[executor.scala 152:13]
    phv_data_491 <= io_pipe_phv_in_data_491; // @[executor.scala 152:13]
    phv_data_492 <= io_pipe_phv_in_data_492; // @[executor.scala 152:13]
    phv_data_493 <= io_pipe_phv_in_data_493; // @[executor.scala 152:13]
    phv_data_494 <= io_pipe_phv_in_data_494; // @[executor.scala 152:13]
    phv_data_495 <= io_pipe_phv_in_data_495; // @[executor.scala 152:13]
    phv_data_496 <= io_pipe_phv_in_data_496; // @[executor.scala 152:13]
    phv_data_497 <= io_pipe_phv_in_data_497; // @[executor.scala 152:13]
    phv_data_498 <= io_pipe_phv_in_data_498; // @[executor.scala 152:13]
    phv_data_499 <= io_pipe_phv_in_data_499; // @[executor.scala 152:13]
    phv_data_500 <= io_pipe_phv_in_data_500; // @[executor.scala 152:13]
    phv_data_501 <= io_pipe_phv_in_data_501; // @[executor.scala 152:13]
    phv_data_502 <= io_pipe_phv_in_data_502; // @[executor.scala 152:13]
    phv_data_503 <= io_pipe_phv_in_data_503; // @[executor.scala 152:13]
    phv_data_504 <= io_pipe_phv_in_data_504; // @[executor.scala 152:13]
    phv_data_505 <= io_pipe_phv_in_data_505; // @[executor.scala 152:13]
    phv_data_506 <= io_pipe_phv_in_data_506; // @[executor.scala 152:13]
    phv_data_507 <= io_pipe_phv_in_data_507; // @[executor.scala 152:13]
    phv_data_508 <= io_pipe_phv_in_data_508; // @[executor.scala 152:13]
    phv_data_509 <= io_pipe_phv_in_data_509; // @[executor.scala 152:13]
    phv_data_510 <= io_pipe_phv_in_data_510; // @[executor.scala 152:13]
    phv_data_511 <= io_pipe_phv_in_data_511; // @[executor.scala 152:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[executor.scala 152:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[executor.scala 152:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[executor.scala 152:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[executor.scala 152:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[executor.scala 152:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[executor.scala 152:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[executor.scala 152:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[executor.scala 152:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[executor.scala 152:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[executor.scala 152:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[executor.scala 152:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[executor.scala 152:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[executor.scala 152:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[executor.scala 152:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[executor.scala 152:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[executor.scala 152:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[executor.scala 152:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[executor.scala 152:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[executor.scala 152:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor.scala 152:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor.scala 152:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor.scala 152:13]
    args_0 <= io_args_in_0; // @[executor.scala 156:14]
    args_1 <= io_args_in_1; // @[executor.scala 156:14]
    args_2 <= io_args_in_2; // @[executor.scala 156:14]
    args_3 <= io_args_in_3; // @[executor.scala 156:14]
    args_4 <= io_args_in_4; // @[executor.scala 156:14]
    args_5 <= io_args_in_5; // @[executor.scala 156:14]
    args_6 <= io_args_in_6; // @[executor.scala 156:14]
    vliw_0 <= io_vliw_in_0; // @[executor.scala 159:14]
    vliw_1 <= io_vliw_in_1; // @[executor.scala 159:14]
    vliw_2 <= io_vliw_in_2; // @[executor.scala 159:14]
    vliw_3 <= io_vliw_in_3; // @[executor.scala 159:14]
    offset_0 <= io_offset_in_0; // @[executor.scala 164:16]
    offset_1 <= io_offset_in_1; // @[executor.scala 164:16]
    offset_2 <= io_offset_in_2; // @[executor.scala 164:16]
    offset_3 <= io_offset_in_3; // @[executor.scala 164:16]
    length_0 <= io_length_in_0; // @[executor.scala 165:16]
    length_1 <= io_length_in_1; // @[executor.scala 165:16]
    length_2 <= io_length_in_2; // @[executor.scala 165:16]
    length_3 <= io_length_in_3; // @[executor.scala 165:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_data_256 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  phv_data_257 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  phv_data_258 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  phv_data_259 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  phv_data_260 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  phv_data_261 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  phv_data_262 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  phv_data_263 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  phv_data_264 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  phv_data_265 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  phv_data_266 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  phv_data_267 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  phv_data_268 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  phv_data_269 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  phv_data_270 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  phv_data_271 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  phv_data_272 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_data_273 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_data_274 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  phv_data_275 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  phv_data_276 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  phv_data_277 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  phv_data_278 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  phv_data_279 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  phv_data_280 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  phv_data_281 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  phv_data_282 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  phv_data_283 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  phv_data_284 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  phv_data_285 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  phv_data_286 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  phv_data_287 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  phv_data_288 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  phv_data_289 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  phv_data_290 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  phv_data_291 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  phv_data_292 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  phv_data_293 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  phv_data_294 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  phv_data_295 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  phv_data_296 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  phv_data_297 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  phv_data_298 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  phv_data_299 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  phv_data_300 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  phv_data_301 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  phv_data_302 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  phv_data_303 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  phv_data_304 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  phv_data_305 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  phv_data_306 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  phv_data_307 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  phv_data_308 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  phv_data_309 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  phv_data_310 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  phv_data_311 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  phv_data_312 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  phv_data_313 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  phv_data_314 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  phv_data_315 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  phv_data_316 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  phv_data_317 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  phv_data_318 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  phv_data_319 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  phv_data_320 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  phv_data_321 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  phv_data_322 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  phv_data_323 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  phv_data_324 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  phv_data_325 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  phv_data_326 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  phv_data_327 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  phv_data_328 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  phv_data_329 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  phv_data_330 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  phv_data_331 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  phv_data_332 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  phv_data_333 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  phv_data_334 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  phv_data_335 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  phv_data_336 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  phv_data_337 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  phv_data_338 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  phv_data_339 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  phv_data_340 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  phv_data_341 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  phv_data_342 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  phv_data_343 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  phv_data_344 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  phv_data_345 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  phv_data_346 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  phv_data_347 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  phv_data_348 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  phv_data_349 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  phv_data_350 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  phv_data_351 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  phv_data_352 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  phv_data_353 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  phv_data_354 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  phv_data_355 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  phv_data_356 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  phv_data_357 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  phv_data_358 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  phv_data_359 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  phv_data_360 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  phv_data_361 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  phv_data_362 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  phv_data_363 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  phv_data_364 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  phv_data_365 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  phv_data_366 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  phv_data_367 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  phv_data_368 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  phv_data_369 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  phv_data_370 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  phv_data_371 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  phv_data_372 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  phv_data_373 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  phv_data_374 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  phv_data_375 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  phv_data_376 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  phv_data_377 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  phv_data_378 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  phv_data_379 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  phv_data_380 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  phv_data_381 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  phv_data_382 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  phv_data_383 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  phv_data_384 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  phv_data_385 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  phv_data_386 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  phv_data_387 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  phv_data_388 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  phv_data_389 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  phv_data_390 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  phv_data_391 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  phv_data_392 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  phv_data_393 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  phv_data_394 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  phv_data_395 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  phv_data_396 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  phv_data_397 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  phv_data_398 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  phv_data_399 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  phv_data_400 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  phv_data_401 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  phv_data_402 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  phv_data_403 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  phv_data_404 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  phv_data_405 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  phv_data_406 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  phv_data_407 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  phv_data_408 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  phv_data_409 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  phv_data_410 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  phv_data_411 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  phv_data_412 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  phv_data_413 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  phv_data_414 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  phv_data_415 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  phv_data_416 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  phv_data_417 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  phv_data_418 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  phv_data_419 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  phv_data_420 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  phv_data_421 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  phv_data_422 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  phv_data_423 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  phv_data_424 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  phv_data_425 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  phv_data_426 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  phv_data_427 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  phv_data_428 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  phv_data_429 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  phv_data_430 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  phv_data_431 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  phv_data_432 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  phv_data_433 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  phv_data_434 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  phv_data_435 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  phv_data_436 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  phv_data_437 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  phv_data_438 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  phv_data_439 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  phv_data_440 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  phv_data_441 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  phv_data_442 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  phv_data_443 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  phv_data_444 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  phv_data_445 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  phv_data_446 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  phv_data_447 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  phv_data_448 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  phv_data_449 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  phv_data_450 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  phv_data_451 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  phv_data_452 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  phv_data_453 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  phv_data_454 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  phv_data_455 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  phv_data_456 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  phv_data_457 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  phv_data_458 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  phv_data_459 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  phv_data_460 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  phv_data_461 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  phv_data_462 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  phv_data_463 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  phv_data_464 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  phv_data_465 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  phv_data_466 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  phv_data_467 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  phv_data_468 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  phv_data_469 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  phv_data_470 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  phv_data_471 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  phv_data_472 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  phv_data_473 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  phv_data_474 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  phv_data_475 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  phv_data_476 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  phv_data_477 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  phv_data_478 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  phv_data_479 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  phv_data_480 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  phv_data_481 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  phv_data_482 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  phv_data_483 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  phv_data_484 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  phv_data_485 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  phv_data_486 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  phv_data_487 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  phv_data_488 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  phv_data_489 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  phv_data_490 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  phv_data_491 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  phv_data_492 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  phv_data_493 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  phv_data_494 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  phv_data_495 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  phv_data_496 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  phv_data_497 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  phv_data_498 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  phv_data_499 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  phv_data_500 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  phv_data_501 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  phv_data_502 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  phv_data_503 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  phv_data_504 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  phv_data_505 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  phv_data_506 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  phv_data_507 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  phv_data_508 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  phv_data_509 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  phv_data_510 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  phv_data_511 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  phv_header_0 = _RAND_512[15:0];
  _RAND_513 = {1{`RANDOM}};
  phv_header_1 = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  phv_header_2 = _RAND_514[15:0];
  _RAND_515 = {1{`RANDOM}};
  phv_header_3 = _RAND_515[15:0];
  _RAND_516 = {1{`RANDOM}};
  phv_header_4 = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  phv_header_5 = _RAND_517[15:0];
  _RAND_518 = {1{`RANDOM}};
  phv_header_6 = _RAND_518[15:0];
  _RAND_519 = {1{`RANDOM}};
  phv_header_7 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  phv_header_8 = _RAND_520[15:0];
  _RAND_521 = {1{`RANDOM}};
  phv_header_9 = _RAND_521[15:0];
  _RAND_522 = {1{`RANDOM}};
  phv_header_10 = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  phv_header_11 = _RAND_523[15:0];
  _RAND_524 = {1{`RANDOM}};
  phv_header_12 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  phv_header_13 = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  phv_header_14 = _RAND_526[15:0];
  _RAND_527 = {1{`RANDOM}};
  phv_header_15 = _RAND_527[15:0];
  _RAND_528 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_530[15:0];
  _RAND_531 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  phv_next_config_id = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  args_0 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  args_1 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  args_2 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  args_3 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  args_4 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  args_5 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  args_6 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  vliw_0 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  vliw_1 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  vliw_2 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  vliw_3 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  offset_0 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  offset_1 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  offset_2 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  offset_3 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  length_0 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  length_1 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  length_2 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  length_3 = _RAND_552[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
