module Processor(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  input         io_pipe_phv_in_valid,
  input         io_pipe_phv_in_last,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_valid,
  output        io_pipe_phv_out_last
);
  wire  PAR_clock; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_0; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_1; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_2; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_3; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_4; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_5; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_6; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_7; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_8; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_9; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_10; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_11; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_12; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_13; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_14; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_16; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_17; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_18; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_19; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_20; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_21; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_22; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_23; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_24; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_25; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_26; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_27; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_28; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_29; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_30; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_31; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_32; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_33; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_34; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_35; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_36; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_37; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_38; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_39; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_40; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_41; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_42; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_43; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_44; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_45; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_46; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_47; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_48; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_49; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_50; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_51; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_52; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_53; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_54; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_55; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_56; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_57; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_58; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_59; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_60; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_61; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_62; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_63; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_64; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_65; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_66; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_67; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_68; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_69; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_70; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_71; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_72; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_73; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_74; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_75; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_76; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_77; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_78; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_79; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_80; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_81; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_82; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_83; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_84; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_85; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_86; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_87; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_88; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_89; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_90; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_91; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_92; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_93; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_94; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_95; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_96; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_97; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_98; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_99; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_100; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_101; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_102; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_103; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_104; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_105; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_106; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_107; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_108; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_109; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_110; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_111; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_112; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_113; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_114; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_115; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_116; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_117; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_118; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_119; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_120; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_121; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_122; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_123; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_124; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_125; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_126; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_127; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_128; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_129; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_130; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_131; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_132; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_133; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_134; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_135; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_136; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_137; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_138; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_139; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_140; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_141; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_142; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_143; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_144; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_145; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_146; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_147; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_148; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_149; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_150; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_151; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_152; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_153; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_154; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_155; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_156; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_157; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_158; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_data_159; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_0; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_1; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_2; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_3; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_4; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_5; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_6; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_7; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_8; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_9; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_10; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_11; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_12; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_13; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_14; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_header_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_parse_current_state; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_in_parse_current_offset; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_in_parse_transition_field; // @[processor.scala 13:21]
  wire [3:0] PAR_io_pipe_phv_in_next_processor_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_next_config_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_is_valid_processor; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_valid; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_in_last; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_0; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_1; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_2; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_3; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_4; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_5; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_6; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_7; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_8; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_9; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_10; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_11; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_12; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_13; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_14; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_16; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_17; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_18; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_19; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_20; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_21; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_22; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_23; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_24; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_25; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_26; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_27; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_28; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_29; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_30; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_31; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_32; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_33; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_34; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_35; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_36; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_37; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_38; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_39; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_40; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_41; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_42; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_43; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_44; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_45; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_46; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_47; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_48; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_49; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_50; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_51; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_52; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_53; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_54; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_55; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_56; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_57; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_58; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_59; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_60; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_61; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_62; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_63; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_64; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_65; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_66; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_67; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_68; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_69; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_70; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_71; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_72; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_73; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_74; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_75; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_76; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_77; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_78; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_79; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_80; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_81; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_82; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_83; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_84; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_85; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_86; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_87; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_88; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_89; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_90; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_91; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_92; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_93; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_94; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_95; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_96; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_97; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_98; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_99; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_100; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_101; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_102; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_103; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_104; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_105; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_106; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_107; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_108; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_109; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_110; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_111; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_112; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_113; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_114; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_115; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_116; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_117; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_118; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_119; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_120; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_121; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_122; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_123; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_124; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_125; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_126; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_127; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_128; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_129; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_130; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_131; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_132; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_133; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_134; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_135; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_136; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_137; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_138; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_139; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_140; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_141; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_142; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_143; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_144; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_145; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_146; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_147; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_148; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_149; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_150; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_151; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_152; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_153; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_154; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_155; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_156; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_157; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_158; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_data_159; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_0; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_1; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_2; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_3; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_4; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_5; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_6; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_7; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_8; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_9; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_10; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_11; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_12; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_13; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_14; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_header_15; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_parse_current_state; // @[processor.scala 13:21]
  wire [7:0] PAR_io_pipe_phv_out_parse_current_offset; // @[processor.scala 13:21]
  wire [15:0] PAR_io_pipe_phv_out_parse_transition_field; // @[processor.scala 13:21]
  wire [3:0] PAR_io_pipe_phv_out_next_processor_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_next_config_id; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_is_valid_processor; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_valid; // @[processor.scala 13:21]
  wire  PAR_io_pipe_phv_out_last; // @[processor.scala 13:21]
  wire  MAT_clock; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_0; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_1; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_2; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_3; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_4; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_5; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_6; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_7; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_8; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_9; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_10; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_11; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_12; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_13; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_14; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_16; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_17; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_18; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_19; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_20; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_21; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_22; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_23; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_24; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_25; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_26; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_27; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_28; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_29; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_30; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_31; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_32; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_33; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_34; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_35; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_36; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_37; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_38; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_39; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_40; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_41; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_42; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_43; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_44; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_45; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_46; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_47; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_48; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_49; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_50; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_51; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_52; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_53; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_54; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_55; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_56; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_57; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_58; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_59; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_60; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_61; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_62; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_63; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_64; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_65; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_66; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_67; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_68; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_69; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_70; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_71; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_72; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_73; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_74; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_75; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_76; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_77; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_78; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_79; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_80; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_81; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_82; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_83; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_84; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_85; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_86; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_87; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_88; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_89; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_90; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_91; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_92; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_93; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_94; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_95; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_96; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_97; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_98; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_99; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_100; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_101; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_102; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_103; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_104; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_105; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_106; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_107; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_108; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_109; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_110; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_111; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_112; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_113; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_114; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_115; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_116; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_117; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_118; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_119; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_120; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_121; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_122; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_123; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_124; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_125; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_126; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_127; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_128; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_129; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_130; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_131; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_132; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_133; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_134; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_135; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_136; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_137; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_138; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_139; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_140; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_141; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_142; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_143; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_144; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_145; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_146; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_147; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_148; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_149; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_150; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_151; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_152; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_153; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_154; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_155; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_156; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_157; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_158; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_data_159; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_0; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_1; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_2; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_3; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_4; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_5; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_6; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_7; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_8; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_9; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_10; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_11; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_12; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_13; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_14; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_header_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_parse_current_state; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_in_parse_current_offset; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_in_parse_transition_field; // @[processor.scala 14:21]
  wire [3:0] MAT_io_pipe_phv_in_next_processor_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_next_config_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_is_valid_processor; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_valid; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_in_last; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_0; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_1; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_2; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_3; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_4; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_5; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_6; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_7; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_8; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_9; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_10; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_11; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_12; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_13; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_14; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_16; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_17; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_18; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_19; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_20; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_21; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_22; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_23; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_24; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_25; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_26; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_27; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_28; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_29; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_30; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_31; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_32; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_33; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_34; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_35; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_36; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_37; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_38; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_39; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_40; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_41; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_42; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_43; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_44; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_45; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_46; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_47; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_48; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_49; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_50; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_51; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_52; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_53; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_54; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_55; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_56; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_57; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_58; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_59; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_60; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_61; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_62; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_63; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_64; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_65; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_66; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_67; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_68; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_69; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_70; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_71; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_72; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_73; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_74; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_75; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_76; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_77; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_78; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_79; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_80; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_81; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_82; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_83; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_84; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_85; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_86; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_87; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_88; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_89; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_90; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_91; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_92; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_93; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_94; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_95; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_96; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_97; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_98; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_99; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_100; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_101; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_102; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_103; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_104; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_105; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_106; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_107; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_108; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_109; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_110; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_111; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_112; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_113; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_114; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_115; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_116; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_117; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_118; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_119; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_120; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_121; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_122; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_123; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_124; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_125; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_126; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_127; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_128; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_129; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_130; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_131; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_132; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_133; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_134; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_135; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_136; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_137; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_138; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_139; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_140; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_141; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_142; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_143; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_144; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_145; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_146; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_147; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_148; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_149; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_150; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_151; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_152; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_153; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_154; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_155; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_156; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_157; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_158; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_data_159; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_0; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_1; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_2; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_3; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_4; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_5; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_6; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_7; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_8; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_9; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_10; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_11; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_12; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_13; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_14; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_header_15; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_parse_current_state; // @[processor.scala 14:21]
  wire [7:0] MAT_io_pipe_phv_out_parse_current_offset; // @[processor.scala 14:21]
  wire [15:0] MAT_io_pipe_phv_out_parse_transition_field; // @[processor.scala 14:21]
  wire [3:0] MAT_io_pipe_phv_out_next_processor_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_next_config_id; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_is_valid_processor; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_valid; // @[processor.scala 14:21]
  wire  MAT_io_pipe_phv_out_last; // @[processor.scala 14:21]
  wire  EXE_clock; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_0; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_2; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_3; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_4; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_5; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_6; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_7; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_8; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_9; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_10; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_11; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_12; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_13; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_14; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_16; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_17; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_18; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_19; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_20; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_21; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_22; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_23; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_24; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_25; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_26; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_27; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_28; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_29; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_30; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_31; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_32; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_33; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_34; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_35; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_36; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_37; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_38; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_39; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_40; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_41; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_42; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_43; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_44; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_45; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_46; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_47; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_48; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_49; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_50; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_51; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_52; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_53; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_54; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_55; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_56; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_57; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_58; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_59; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_60; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_61; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_62; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_63; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_64; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_65; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_66; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_67; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_68; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_69; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_70; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_71; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_72; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_73; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_74; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_75; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_76; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_77; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_78; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_79; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_80; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_81; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_82; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_83; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_84; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_85; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_86; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_87; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_88; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_89; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_90; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_91; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_92; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_93; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_94; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_95; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_96; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_97; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_98; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_99; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_100; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_101; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_102; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_103; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_104; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_105; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_106; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_107; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_108; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_109; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_110; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_111; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_112; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_113; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_114; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_115; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_116; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_117; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_118; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_119; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_120; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_121; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_122; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_123; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_124; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_125; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_126; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_127; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_128; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_129; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_130; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_131; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_132; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_133; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_134; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_135; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_136; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_137; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_138; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_139; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_140; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_141; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_142; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_143; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_144; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_145; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_146; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_147; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_148; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_149; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_150; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_151; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_152; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_153; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_154; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_155; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_156; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_157; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_158; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_data_159; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_0; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_1; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_2; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_3; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_4; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_5; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_6; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_7; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_8; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_9; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_10; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_11; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_12; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_13; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_14; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_header_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_parse_current_state; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_in_parse_current_offset; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_in_parse_transition_field; // @[processor.scala 15:21]
  wire [3:0] EXE_io_pipe_phv_in_next_processor_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_next_config_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_is_valid_processor; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_valid; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_in_last; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_0; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_1; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_2; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_3; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_4; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_5; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_6; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_7; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_8; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_9; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_10; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_11; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_12; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_13; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_14; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_16; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_17; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_18; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_19; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_20; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_21; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_22; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_23; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_24; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_25; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_26; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_27; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_28; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_29; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_30; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_31; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_32; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_33; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_34; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_35; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_36; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_37; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_38; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_39; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_40; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_41; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_42; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_43; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_44; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_45; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_46; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_47; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_48; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_49; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_50; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_51; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_52; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_53; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_54; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_55; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_56; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_57; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_58; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_59; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_60; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_61; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_62; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_63; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_64; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_65; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_66; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_67; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_68; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_69; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_70; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_71; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_72; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_73; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_74; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_75; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_76; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_77; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_78; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_79; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_80; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_81; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_82; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_83; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_84; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_85; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_86; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_87; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_88; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_89; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_90; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_91; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_92; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_93; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_94; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_95; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_96; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_97; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_98; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_99; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_100; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_101; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_102; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_103; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_104; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_105; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_106; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_107; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_108; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_109; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_110; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_111; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_112; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_113; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_114; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_115; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_116; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_117; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_118; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_119; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_120; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_121; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_122; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_123; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_124; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_125; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_126; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_127; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_128; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_129; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_130; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_131; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_132; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_133; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_134; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_135; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_136; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_137; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_138; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_139; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_140; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_141; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_142; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_143; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_144; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_145; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_146; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_147; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_148; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_149; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_150; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_151; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_152; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_153; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_154; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_155; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_156; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_157; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_158; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_data_159; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_0; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_1; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_2; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_3; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_4; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_5; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_6; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_7; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_8; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_9; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_10; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_11; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_12; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_13; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_14; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_header_15; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_parse_current_state; // @[processor.scala 15:21]
  wire [7:0] EXE_io_pipe_phv_out_parse_current_offset; // @[processor.scala 15:21]
  wire [15:0] EXE_io_pipe_phv_out_parse_transition_field; // @[processor.scala 15:21]
  wire [3:0] EXE_io_pipe_phv_out_next_processor_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_out_next_config_id; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_out_valid; // @[processor.scala 15:21]
  wire  EXE_io_pipe_phv_out_last; // @[processor.scala 15:21]
  Parser PAR ( // @[processor.scala 13:21]
    .clock(PAR_clock),
    .io_pipe_phv_in_data_0(PAR_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(PAR_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(PAR_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(PAR_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(PAR_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(PAR_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(PAR_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(PAR_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(PAR_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(PAR_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(PAR_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(PAR_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(PAR_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(PAR_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(PAR_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(PAR_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(PAR_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(PAR_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(PAR_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(PAR_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(PAR_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(PAR_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(PAR_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(PAR_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(PAR_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(PAR_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(PAR_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(PAR_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(PAR_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(PAR_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(PAR_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(PAR_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(PAR_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(PAR_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(PAR_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(PAR_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(PAR_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(PAR_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(PAR_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(PAR_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(PAR_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(PAR_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(PAR_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(PAR_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(PAR_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(PAR_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(PAR_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(PAR_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(PAR_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(PAR_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(PAR_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(PAR_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(PAR_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(PAR_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(PAR_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(PAR_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(PAR_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(PAR_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(PAR_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(PAR_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(PAR_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(PAR_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(PAR_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(PAR_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(PAR_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(PAR_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(PAR_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(PAR_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(PAR_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(PAR_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(PAR_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(PAR_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(PAR_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(PAR_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(PAR_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(PAR_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(PAR_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(PAR_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(PAR_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(PAR_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(PAR_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(PAR_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(PAR_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(PAR_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(PAR_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(PAR_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(PAR_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(PAR_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(PAR_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(PAR_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(PAR_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(PAR_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(PAR_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(PAR_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(PAR_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(PAR_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(PAR_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(PAR_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(PAR_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(PAR_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(PAR_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(PAR_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(PAR_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(PAR_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(PAR_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(PAR_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(PAR_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(PAR_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(PAR_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(PAR_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(PAR_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(PAR_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(PAR_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(PAR_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(PAR_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(PAR_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(PAR_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(PAR_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(PAR_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(PAR_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(PAR_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(PAR_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(PAR_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(PAR_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(PAR_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(PAR_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(PAR_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(PAR_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(PAR_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(PAR_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(PAR_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(PAR_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(PAR_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(PAR_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(PAR_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(PAR_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(PAR_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(PAR_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(PAR_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(PAR_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(PAR_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(PAR_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(PAR_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(PAR_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(PAR_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(PAR_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(PAR_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(PAR_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(PAR_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(PAR_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(PAR_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(PAR_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(PAR_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(PAR_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(PAR_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(PAR_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(PAR_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(PAR_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(PAR_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(PAR_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(PAR_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(PAR_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(PAR_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(PAR_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(PAR_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(PAR_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(PAR_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(PAR_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(PAR_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(PAR_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(PAR_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(PAR_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(PAR_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(PAR_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(PAR_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(PAR_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(PAR_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(PAR_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(PAR_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(PAR_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(PAR_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(PAR_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(PAR_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(PAR_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(PAR_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(PAR_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(PAR_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(PAR_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(PAR_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(PAR_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(PAR_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(PAR_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(PAR_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(PAR_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(PAR_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(PAR_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(PAR_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(PAR_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(PAR_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(PAR_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(PAR_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(PAR_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(PAR_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(PAR_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(PAR_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(PAR_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(PAR_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(PAR_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(PAR_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(PAR_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(PAR_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(PAR_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(PAR_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(PAR_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(PAR_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(PAR_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(PAR_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(PAR_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(PAR_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(PAR_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(PAR_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(PAR_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(PAR_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(PAR_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(PAR_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(PAR_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(PAR_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(PAR_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(PAR_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(PAR_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(PAR_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(PAR_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(PAR_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(PAR_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(PAR_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(PAR_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(PAR_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(PAR_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(PAR_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(PAR_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(PAR_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(PAR_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(PAR_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(PAR_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(PAR_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(PAR_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(PAR_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(PAR_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(PAR_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(PAR_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(PAR_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(PAR_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(PAR_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(PAR_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(PAR_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(PAR_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(PAR_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(PAR_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(PAR_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(PAR_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(PAR_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(PAR_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(PAR_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(PAR_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(PAR_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(PAR_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(PAR_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(PAR_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(PAR_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(PAR_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(PAR_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(PAR_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(PAR_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(PAR_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(PAR_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(PAR_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(PAR_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(PAR_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(PAR_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(PAR_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(PAR_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(PAR_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(PAR_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(PAR_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(PAR_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(PAR_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(PAR_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(PAR_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(PAR_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(PAR_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(PAR_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(PAR_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(PAR_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(PAR_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(PAR_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(PAR_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(PAR_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(PAR_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(PAR_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(PAR_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(PAR_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(PAR_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(PAR_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(PAR_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(PAR_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(PAR_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(PAR_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(PAR_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(PAR_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(PAR_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(PAR_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(PAR_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(PAR_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(PAR_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(PAR_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(PAR_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(PAR_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(PAR_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(PAR_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(PAR_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(PAR_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(PAR_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(PAR_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(PAR_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(PAR_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(PAR_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(PAR_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(PAR_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(PAR_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(PAR_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(PAR_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(PAR_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(PAR_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(PAR_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(PAR_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(PAR_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(PAR_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(PAR_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(PAR_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(PAR_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(PAR_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(PAR_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(PAR_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(PAR_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(PAR_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(PAR_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(PAR_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(PAR_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(PAR_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(PAR_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(PAR_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(PAR_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(PAR_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(PAR_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(PAR_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(PAR_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(PAR_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(PAR_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(PAR_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(PAR_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(PAR_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(PAR_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(PAR_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(PAR_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(PAR_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(PAR_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(PAR_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(PAR_io_pipe_phv_out_last)
  );
  Matcher MAT ( // @[processor.scala 14:21]
    .clock(MAT_clock),
    .io_pipe_phv_in_data_0(MAT_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(MAT_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(MAT_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(MAT_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(MAT_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(MAT_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(MAT_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(MAT_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(MAT_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(MAT_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(MAT_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(MAT_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(MAT_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(MAT_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(MAT_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(MAT_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(MAT_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(MAT_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(MAT_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(MAT_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(MAT_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(MAT_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(MAT_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(MAT_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(MAT_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(MAT_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(MAT_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(MAT_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(MAT_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(MAT_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(MAT_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(MAT_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(MAT_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(MAT_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(MAT_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(MAT_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(MAT_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(MAT_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(MAT_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(MAT_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(MAT_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(MAT_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(MAT_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(MAT_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(MAT_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(MAT_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(MAT_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(MAT_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(MAT_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(MAT_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(MAT_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(MAT_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(MAT_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(MAT_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(MAT_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(MAT_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(MAT_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(MAT_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(MAT_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(MAT_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(MAT_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(MAT_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(MAT_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(MAT_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(MAT_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(MAT_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(MAT_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(MAT_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(MAT_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(MAT_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(MAT_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(MAT_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(MAT_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(MAT_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(MAT_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(MAT_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(MAT_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(MAT_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(MAT_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(MAT_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(MAT_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(MAT_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(MAT_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(MAT_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(MAT_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(MAT_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(MAT_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(MAT_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(MAT_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(MAT_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(MAT_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(MAT_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(MAT_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(MAT_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(MAT_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(MAT_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(MAT_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(MAT_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(MAT_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(MAT_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(MAT_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(MAT_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(MAT_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(MAT_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(MAT_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(MAT_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(MAT_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(MAT_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(MAT_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(MAT_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(MAT_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(MAT_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(MAT_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(MAT_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(MAT_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(MAT_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(MAT_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(MAT_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(MAT_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(MAT_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(MAT_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(MAT_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(MAT_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(MAT_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(MAT_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(MAT_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(MAT_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(MAT_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(MAT_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(MAT_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(MAT_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(MAT_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(MAT_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(MAT_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(MAT_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(MAT_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(MAT_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(MAT_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(MAT_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(MAT_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(MAT_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(MAT_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(MAT_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(MAT_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(MAT_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(MAT_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(MAT_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(MAT_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(MAT_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(MAT_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(MAT_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(MAT_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(MAT_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(MAT_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(MAT_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(MAT_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(MAT_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(MAT_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(MAT_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(MAT_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(MAT_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(MAT_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(MAT_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(MAT_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(MAT_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(MAT_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(MAT_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(MAT_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(MAT_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(MAT_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(MAT_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(MAT_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(MAT_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(MAT_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(MAT_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(MAT_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(MAT_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(MAT_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(MAT_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(MAT_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(MAT_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(MAT_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(MAT_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(MAT_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(MAT_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(MAT_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(MAT_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(MAT_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(MAT_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(MAT_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(MAT_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(MAT_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(MAT_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(MAT_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(MAT_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(MAT_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(MAT_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(MAT_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(MAT_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(MAT_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(MAT_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(MAT_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(MAT_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(MAT_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(MAT_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(MAT_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(MAT_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(MAT_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(MAT_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(MAT_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(MAT_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(MAT_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(MAT_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(MAT_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(MAT_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(MAT_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(MAT_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(MAT_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(MAT_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(MAT_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(MAT_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(MAT_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(MAT_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(MAT_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(MAT_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(MAT_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(MAT_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(MAT_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(MAT_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(MAT_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(MAT_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(MAT_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(MAT_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(MAT_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(MAT_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(MAT_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(MAT_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(MAT_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(MAT_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(MAT_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(MAT_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(MAT_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(MAT_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(MAT_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(MAT_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(MAT_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(MAT_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(MAT_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(MAT_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(MAT_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(MAT_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(MAT_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(MAT_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(MAT_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(MAT_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(MAT_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(MAT_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(MAT_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(MAT_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(MAT_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(MAT_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(MAT_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(MAT_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(MAT_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(MAT_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(MAT_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(MAT_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(MAT_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(MAT_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(MAT_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(MAT_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(MAT_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(MAT_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(MAT_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(MAT_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(MAT_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(MAT_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(MAT_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(MAT_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(MAT_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(MAT_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(MAT_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(MAT_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(MAT_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(MAT_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(MAT_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(MAT_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(MAT_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(MAT_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(MAT_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(MAT_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(MAT_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(MAT_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(MAT_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(MAT_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(MAT_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(MAT_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(MAT_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(MAT_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(MAT_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(MAT_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(MAT_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(MAT_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(MAT_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(MAT_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(MAT_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(MAT_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(MAT_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(MAT_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(MAT_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(MAT_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(MAT_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(MAT_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(MAT_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(MAT_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(MAT_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(MAT_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(MAT_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(MAT_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(MAT_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(MAT_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(MAT_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(MAT_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(MAT_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(MAT_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(MAT_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(MAT_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(MAT_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(MAT_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(MAT_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(MAT_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(MAT_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(MAT_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(MAT_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(MAT_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(MAT_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(MAT_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(MAT_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(MAT_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(MAT_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(MAT_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(MAT_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(MAT_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(MAT_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(MAT_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(MAT_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(MAT_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(MAT_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(MAT_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(MAT_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(MAT_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(MAT_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(MAT_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(MAT_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(MAT_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(MAT_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(MAT_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(MAT_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(MAT_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(MAT_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(MAT_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(MAT_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(MAT_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(MAT_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(MAT_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(MAT_io_pipe_phv_out_is_valid_processor),
    .io_pipe_phv_out_valid(MAT_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(MAT_io_pipe_phv_out_last)
  );
  Executor EXE ( // @[processor.scala 15:21]
    .clock(EXE_clock),
    .io_pipe_phv_in_data_0(EXE_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(EXE_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(EXE_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(EXE_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(EXE_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(EXE_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(EXE_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(EXE_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(EXE_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(EXE_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(EXE_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(EXE_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(EXE_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(EXE_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(EXE_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(EXE_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(EXE_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(EXE_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(EXE_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(EXE_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(EXE_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(EXE_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(EXE_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(EXE_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(EXE_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(EXE_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(EXE_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(EXE_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(EXE_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(EXE_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(EXE_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(EXE_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(EXE_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(EXE_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(EXE_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(EXE_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(EXE_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(EXE_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(EXE_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(EXE_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(EXE_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(EXE_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(EXE_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(EXE_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(EXE_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(EXE_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(EXE_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(EXE_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(EXE_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(EXE_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(EXE_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(EXE_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(EXE_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(EXE_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(EXE_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(EXE_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(EXE_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(EXE_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(EXE_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(EXE_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(EXE_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(EXE_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(EXE_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(EXE_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(EXE_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(EXE_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(EXE_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(EXE_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(EXE_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(EXE_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(EXE_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(EXE_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(EXE_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(EXE_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(EXE_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(EXE_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(EXE_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(EXE_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(EXE_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(EXE_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(EXE_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(EXE_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(EXE_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(EXE_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(EXE_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(EXE_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(EXE_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(EXE_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(EXE_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(EXE_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(EXE_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(EXE_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(EXE_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(EXE_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(EXE_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(EXE_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(EXE_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(EXE_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(EXE_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(EXE_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(EXE_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(EXE_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(EXE_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(EXE_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(EXE_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(EXE_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(EXE_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(EXE_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(EXE_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(EXE_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(EXE_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(EXE_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(EXE_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(EXE_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(EXE_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(EXE_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(EXE_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(EXE_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(EXE_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(EXE_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(EXE_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(EXE_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(EXE_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(EXE_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(EXE_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(EXE_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(EXE_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(EXE_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(EXE_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(EXE_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(EXE_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(EXE_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(EXE_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(EXE_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(EXE_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(EXE_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(EXE_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(EXE_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(EXE_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(EXE_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(EXE_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(EXE_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(EXE_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(EXE_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(EXE_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(EXE_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(EXE_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(EXE_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(EXE_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(EXE_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(EXE_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(EXE_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(EXE_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(EXE_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(EXE_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(EXE_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(EXE_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(EXE_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(EXE_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(EXE_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(EXE_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(EXE_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(EXE_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(EXE_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(EXE_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(EXE_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(EXE_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(EXE_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(EXE_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(EXE_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(EXE_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(EXE_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(EXE_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(EXE_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(EXE_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(EXE_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(EXE_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(EXE_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(EXE_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(EXE_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(EXE_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(EXE_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_in_valid(EXE_io_pipe_phv_in_valid),
    .io_pipe_phv_in_last(EXE_io_pipe_phv_in_last),
    .io_pipe_phv_out_data_0(EXE_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(EXE_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(EXE_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(EXE_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(EXE_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(EXE_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(EXE_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(EXE_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(EXE_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(EXE_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(EXE_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(EXE_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(EXE_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(EXE_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(EXE_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(EXE_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(EXE_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(EXE_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(EXE_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(EXE_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(EXE_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(EXE_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(EXE_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(EXE_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(EXE_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(EXE_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(EXE_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(EXE_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(EXE_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(EXE_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(EXE_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(EXE_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(EXE_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(EXE_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(EXE_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(EXE_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(EXE_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(EXE_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(EXE_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(EXE_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(EXE_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(EXE_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(EXE_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(EXE_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(EXE_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(EXE_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(EXE_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(EXE_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(EXE_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(EXE_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(EXE_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(EXE_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(EXE_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(EXE_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(EXE_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(EXE_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(EXE_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(EXE_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(EXE_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(EXE_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(EXE_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(EXE_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(EXE_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(EXE_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(EXE_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(EXE_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(EXE_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(EXE_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(EXE_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(EXE_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(EXE_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(EXE_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(EXE_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(EXE_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(EXE_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(EXE_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(EXE_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(EXE_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(EXE_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(EXE_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(EXE_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(EXE_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(EXE_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(EXE_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(EXE_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(EXE_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(EXE_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(EXE_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(EXE_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(EXE_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(EXE_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(EXE_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(EXE_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(EXE_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(EXE_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(EXE_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(EXE_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(EXE_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(EXE_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(EXE_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(EXE_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(EXE_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(EXE_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(EXE_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(EXE_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(EXE_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(EXE_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(EXE_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(EXE_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(EXE_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(EXE_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(EXE_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(EXE_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(EXE_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(EXE_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(EXE_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(EXE_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(EXE_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(EXE_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(EXE_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(EXE_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(EXE_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(EXE_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(EXE_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(EXE_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(EXE_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(EXE_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(EXE_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(EXE_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(EXE_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(EXE_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(EXE_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(EXE_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(EXE_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(EXE_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(EXE_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(EXE_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(EXE_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(EXE_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(EXE_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(EXE_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(EXE_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(EXE_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(EXE_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(EXE_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(EXE_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(EXE_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(EXE_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(EXE_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(EXE_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(EXE_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(EXE_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(EXE_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(EXE_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(EXE_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(EXE_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(EXE_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(EXE_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(EXE_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(EXE_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(EXE_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(EXE_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(EXE_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(EXE_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(EXE_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(EXE_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(EXE_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(EXE_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(EXE_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(EXE_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(EXE_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(EXE_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(EXE_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(EXE_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(EXE_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(EXE_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(EXE_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(EXE_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(EXE_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(EXE_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(EXE_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_valid(EXE_io_pipe_phv_out_valid),
    .io_pipe_phv_out_last(EXE_io_pipe_phv_out_last)
  );
  assign io_pipe_phv_out_data_0 = EXE_io_pipe_phv_out_data_0; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_1 = EXE_io_pipe_phv_out_data_1; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_2 = EXE_io_pipe_phv_out_data_2; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_3 = EXE_io_pipe_phv_out_data_3; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_4 = EXE_io_pipe_phv_out_data_4; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_5 = EXE_io_pipe_phv_out_data_5; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_6 = EXE_io_pipe_phv_out_data_6; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_7 = EXE_io_pipe_phv_out_data_7; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_8 = EXE_io_pipe_phv_out_data_8; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_9 = EXE_io_pipe_phv_out_data_9; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_10 = EXE_io_pipe_phv_out_data_10; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_11 = EXE_io_pipe_phv_out_data_11; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_12 = EXE_io_pipe_phv_out_data_12; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_13 = EXE_io_pipe_phv_out_data_13; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_14 = EXE_io_pipe_phv_out_data_14; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_15 = EXE_io_pipe_phv_out_data_15; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_16 = EXE_io_pipe_phv_out_data_16; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_17 = EXE_io_pipe_phv_out_data_17; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_18 = EXE_io_pipe_phv_out_data_18; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_19 = EXE_io_pipe_phv_out_data_19; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_20 = EXE_io_pipe_phv_out_data_20; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_21 = EXE_io_pipe_phv_out_data_21; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_22 = EXE_io_pipe_phv_out_data_22; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_23 = EXE_io_pipe_phv_out_data_23; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_24 = EXE_io_pipe_phv_out_data_24; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_25 = EXE_io_pipe_phv_out_data_25; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_26 = EXE_io_pipe_phv_out_data_26; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_27 = EXE_io_pipe_phv_out_data_27; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_28 = EXE_io_pipe_phv_out_data_28; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_29 = EXE_io_pipe_phv_out_data_29; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_30 = EXE_io_pipe_phv_out_data_30; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_31 = EXE_io_pipe_phv_out_data_31; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_32 = EXE_io_pipe_phv_out_data_32; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_33 = EXE_io_pipe_phv_out_data_33; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_34 = EXE_io_pipe_phv_out_data_34; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_35 = EXE_io_pipe_phv_out_data_35; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_36 = EXE_io_pipe_phv_out_data_36; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_37 = EXE_io_pipe_phv_out_data_37; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_38 = EXE_io_pipe_phv_out_data_38; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_39 = EXE_io_pipe_phv_out_data_39; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_40 = EXE_io_pipe_phv_out_data_40; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_41 = EXE_io_pipe_phv_out_data_41; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_42 = EXE_io_pipe_phv_out_data_42; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_43 = EXE_io_pipe_phv_out_data_43; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_44 = EXE_io_pipe_phv_out_data_44; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_45 = EXE_io_pipe_phv_out_data_45; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_46 = EXE_io_pipe_phv_out_data_46; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_47 = EXE_io_pipe_phv_out_data_47; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_48 = EXE_io_pipe_phv_out_data_48; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_49 = EXE_io_pipe_phv_out_data_49; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_50 = EXE_io_pipe_phv_out_data_50; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_51 = EXE_io_pipe_phv_out_data_51; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_52 = EXE_io_pipe_phv_out_data_52; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_53 = EXE_io_pipe_phv_out_data_53; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_54 = EXE_io_pipe_phv_out_data_54; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_55 = EXE_io_pipe_phv_out_data_55; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_56 = EXE_io_pipe_phv_out_data_56; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_57 = EXE_io_pipe_phv_out_data_57; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_58 = EXE_io_pipe_phv_out_data_58; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_59 = EXE_io_pipe_phv_out_data_59; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_60 = EXE_io_pipe_phv_out_data_60; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_61 = EXE_io_pipe_phv_out_data_61; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_62 = EXE_io_pipe_phv_out_data_62; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_63 = EXE_io_pipe_phv_out_data_63; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_64 = EXE_io_pipe_phv_out_data_64; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_65 = EXE_io_pipe_phv_out_data_65; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_66 = EXE_io_pipe_phv_out_data_66; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_67 = EXE_io_pipe_phv_out_data_67; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_68 = EXE_io_pipe_phv_out_data_68; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_69 = EXE_io_pipe_phv_out_data_69; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_70 = EXE_io_pipe_phv_out_data_70; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_71 = EXE_io_pipe_phv_out_data_71; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_72 = EXE_io_pipe_phv_out_data_72; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_73 = EXE_io_pipe_phv_out_data_73; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_74 = EXE_io_pipe_phv_out_data_74; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_75 = EXE_io_pipe_phv_out_data_75; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_76 = EXE_io_pipe_phv_out_data_76; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_77 = EXE_io_pipe_phv_out_data_77; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_78 = EXE_io_pipe_phv_out_data_78; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_79 = EXE_io_pipe_phv_out_data_79; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_80 = EXE_io_pipe_phv_out_data_80; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_81 = EXE_io_pipe_phv_out_data_81; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_82 = EXE_io_pipe_phv_out_data_82; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_83 = EXE_io_pipe_phv_out_data_83; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_84 = EXE_io_pipe_phv_out_data_84; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_85 = EXE_io_pipe_phv_out_data_85; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_86 = EXE_io_pipe_phv_out_data_86; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_87 = EXE_io_pipe_phv_out_data_87; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_88 = EXE_io_pipe_phv_out_data_88; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_89 = EXE_io_pipe_phv_out_data_89; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_90 = EXE_io_pipe_phv_out_data_90; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_91 = EXE_io_pipe_phv_out_data_91; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_92 = EXE_io_pipe_phv_out_data_92; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_93 = EXE_io_pipe_phv_out_data_93; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_94 = EXE_io_pipe_phv_out_data_94; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_95 = EXE_io_pipe_phv_out_data_95; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_96 = EXE_io_pipe_phv_out_data_96; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_97 = EXE_io_pipe_phv_out_data_97; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_98 = EXE_io_pipe_phv_out_data_98; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_99 = EXE_io_pipe_phv_out_data_99; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_100 = EXE_io_pipe_phv_out_data_100; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_101 = EXE_io_pipe_phv_out_data_101; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_102 = EXE_io_pipe_phv_out_data_102; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_103 = EXE_io_pipe_phv_out_data_103; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_104 = EXE_io_pipe_phv_out_data_104; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_105 = EXE_io_pipe_phv_out_data_105; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_106 = EXE_io_pipe_phv_out_data_106; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_107 = EXE_io_pipe_phv_out_data_107; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_108 = EXE_io_pipe_phv_out_data_108; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_109 = EXE_io_pipe_phv_out_data_109; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_110 = EXE_io_pipe_phv_out_data_110; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_111 = EXE_io_pipe_phv_out_data_111; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_112 = EXE_io_pipe_phv_out_data_112; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_113 = EXE_io_pipe_phv_out_data_113; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_114 = EXE_io_pipe_phv_out_data_114; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_115 = EXE_io_pipe_phv_out_data_115; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_116 = EXE_io_pipe_phv_out_data_116; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_117 = EXE_io_pipe_phv_out_data_117; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_118 = EXE_io_pipe_phv_out_data_118; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_119 = EXE_io_pipe_phv_out_data_119; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_120 = EXE_io_pipe_phv_out_data_120; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_121 = EXE_io_pipe_phv_out_data_121; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_122 = EXE_io_pipe_phv_out_data_122; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_123 = EXE_io_pipe_phv_out_data_123; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_124 = EXE_io_pipe_phv_out_data_124; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_125 = EXE_io_pipe_phv_out_data_125; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_126 = EXE_io_pipe_phv_out_data_126; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_127 = EXE_io_pipe_phv_out_data_127; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_128 = EXE_io_pipe_phv_out_data_128; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_129 = EXE_io_pipe_phv_out_data_129; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_130 = EXE_io_pipe_phv_out_data_130; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_131 = EXE_io_pipe_phv_out_data_131; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_132 = EXE_io_pipe_phv_out_data_132; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_133 = EXE_io_pipe_phv_out_data_133; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_134 = EXE_io_pipe_phv_out_data_134; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_135 = EXE_io_pipe_phv_out_data_135; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_136 = EXE_io_pipe_phv_out_data_136; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_137 = EXE_io_pipe_phv_out_data_137; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_138 = EXE_io_pipe_phv_out_data_138; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_139 = EXE_io_pipe_phv_out_data_139; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_140 = EXE_io_pipe_phv_out_data_140; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_141 = EXE_io_pipe_phv_out_data_141; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_142 = EXE_io_pipe_phv_out_data_142; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_143 = EXE_io_pipe_phv_out_data_143; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_144 = EXE_io_pipe_phv_out_data_144; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_145 = EXE_io_pipe_phv_out_data_145; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_146 = EXE_io_pipe_phv_out_data_146; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_147 = EXE_io_pipe_phv_out_data_147; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_148 = EXE_io_pipe_phv_out_data_148; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_149 = EXE_io_pipe_phv_out_data_149; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_150 = EXE_io_pipe_phv_out_data_150; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_151 = EXE_io_pipe_phv_out_data_151; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_152 = EXE_io_pipe_phv_out_data_152; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_153 = EXE_io_pipe_phv_out_data_153; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_154 = EXE_io_pipe_phv_out_data_154; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_155 = EXE_io_pipe_phv_out_data_155; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_156 = EXE_io_pipe_phv_out_data_156; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_157 = EXE_io_pipe_phv_out_data_157; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_158 = EXE_io_pipe_phv_out_data_158; // @[processor.scala 29:24]
  assign io_pipe_phv_out_data_159 = EXE_io_pipe_phv_out_data_159; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_0 = EXE_io_pipe_phv_out_header_0; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_1 = EXE_io_pipe_phv_out_header_1; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_2 = EXE_io_pipe_phv_out_header_2; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_3 = EXE_io_pipe_phv_out_header_3; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_4 = EXE_io_pipe_phv_out_header_4; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_5 = EXE_io_pipe_phv_out_header_5; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_6 = EXE_io_pipe_phv_out_header_6; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_7 = EXE_io_pipe_phv_out_header_7; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_8 = EXE_io_pipe_phv_out_header_8; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_9 = EXE_io_pipe_phv_out_header_9; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_10 = EXE_io_pipe_phv_out_header_10; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_11 = EXE_io_pipe_phv_out_header_11; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_12 = EXE_io_pipe_phv_out_header_12; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_13 = EXE_io_pipe_phv_out_header_13; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_14 = EXE_io_pipe_phv_out_header_14; // @[processor.scala 29:24]
  assign io_pipe_phv_out_header_15 = EXE_io_pipe_phv_out_header_15; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_current_state = EXE_io_pipe_phv_out_parse_current_state; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_current_offset = EXE_io_pipe_phv_out_parse_current_offset; // @[processor.scala 29:24]
  assign io_pipe_phv_out_parse_transition_field = EXE_io_pipe_phv_out_parse_transition_field; // @[processor.scala 29:24]
  assign io_pipe_phv_out_next_processor_id = EXE_io_pipe_phv_out_next_processor_id; // @[processor.scala 29:24]
  assign io_pipe_phv_out_next_config_id = EXE_io_pipe_phv_out_next_config_id; // @[processor.scala 29:24]
  assign io_pipe_phv_out_valid = EXE_io_pipe_phv_out_valid; // @[processor.scala 29:24]
  assign io_pipe_phv_out_last = EXE_io_pipe_phv_out_last; // @[processor.scala 29:24]
  assign PAR_clock = clock;
  assign PAR_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_valid = io_pipe_phv_in_valid; // @[processor.scala 17:24]
  assign PAR_io_pipe_phv_in_last = io_pipe_phv_in_last; // @[processor.scala 17:24]
  assign MAT_clock = clock;
  assign MAT_io_pipe_phv_in_data_0 = PAR_io_pipe_phv_out_data_0; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_1 = PAR_io_pipe_phv_out_data_1; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_2 = PAR_io_pipe_phv_out_data_2; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_3 = PAR_io_pipe_phv_out_data_3; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_4 = PAR_io_pipe_phv_out_data_4; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_5 = PAR_io_pipe_phv_out_data_5; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_6 = PAR_io_pipe_phv_out_data_6; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_7 = PAR_io_pipe_phv_out_data_7; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_8 = PAR_io_pipe_phv_out_data_8; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_9 = PAR_io_pipe_phv_out_data_9; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_10 = PAR_io_pipe_phv_out_data_10; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_11 = PAR_io_pipe_phv_out_data_11; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_12 = PAR_io_pipe_phv_out_data_12; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_13 = PAR_io_pipe_phv_out_data_13; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_14 = PAR_io_pipe_phv_out_data_14; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_15 = PAR_io_pipe_phv_out_data_15; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_16 = PAR_io_pipe_phv_out_data_16; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_17 = PAR_io_pipe_phv_out_data_17; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_18 = PAR_io_pipe_phv_out_data_18; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_19 = PAR_io_pipe_phv_out_data_19; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_20 = PAR_io_pipe_phv_out_data_20; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_21 = PAR_io_pipe_phv_out_data_21; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_22 = PAR_io_pipe_phv_out_data_22; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_23 = PAR_io_pipe_phv_out_data_23; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_24 = PAR_io_pipe_phv_out_data_24; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_25 = PAR_io_pipe_phv_out_data_25; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_26 = PAR_io_pipe_phv_out_data_26; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_27 = PAR_io_pipe_phv_out_data_27; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_28 = PAR_io_pipe_phv_out_data_28; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_29 = PAR_io_pipe_phv_out_data_29; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_30 = PAR_io_pipe_phv_out_data_30; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_31 = PAR_io_pipe_phv_out_data_31; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_32 = PAR_io_pipe_phv_out_data_32; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_33 = PAR_io_pipe_phv_out_data_33; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_34 = PAR_io_pipe_phv_out_data_34; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_35 = PAR_io_pipe_phv_out_data_35; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_36 = PAR_io_pipe_phv_out_data_36; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_37 = PAR_io_pipe_phv_out_data_37; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_38 = PAR_io_pipe_phv_out_data_38; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_39 = PAR_io_pipe_phv_out_data_39; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_40 = PAR_io_pipe_phv_out_data_40; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_41 = PAR_io_pipe_phv_out_data_41; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_42 = PAR_io_pipe_phv_out_data_42; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_43 = PAR_io_pipe_phv_out_data_43; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_44 = PAR_io_pipe_phv_out_data_44; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_45 = PAR_io_pipe_phv_out_data_45; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_46 = PAR_io_pipe_phv_out_data_46; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_47 = PAR_io_pipe_phv_out_data_47; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_48 = PAR_io_pipe_phv_out_data_48; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_49 = PAR_io_pipe_phv_out_data_49; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_50 = PAR_io_pipe_phv_out_data_50; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_51 = PAR_io_pipe_phv_out_data_51; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_52 = PAR_io_pipe_phv_out_data_52; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_53 = PAR_io_pipe_phv_out_data_53; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_54 = PAR_io_pipe_phv_out_data_54; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_55 = PAR_io_pipe_phv_out_data_55; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_56 = PAR_io_pipe_phv_out_data_56; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_57 = PAR_io_pipe_phv_out_data_57; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_58 = PAR_io_pipe_phv_out_data_58; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_59 = PAR_io_pipe_phv_out_data_59; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_60 = PAR_io_pipe_phv_out_data_60; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_61 = PAR_io_pipe_phv_out_data_61; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_62 = PAR_io_pipe_phv_out_data_62; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_63 = PAR_io_pipe_phv_out_data_63; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_64 = PAR_io_pipe_phv_out_data_64; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_65 = PAR_io_pipe_phv_out_data_65; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_66 = PAR_io_pipe_phv_out_data_66; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_67 = PAR_io_pipe_phv_out_data_67; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_68 = PAR_io_pipe_phv_out_data_68; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_69 = PAR_io_pipe_phv_out_data_69; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_70 = PAR_io_pipe_phv_out_data_70; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_71 = PAR_io_pipe_phv_out_data_71; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_72 = PAR_io_pipe_phv_out_data_72; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_73 = PAR_io_pipe_phv_out_data_73; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_74 = PAR_io_pipe_phv_out_data_74; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_75 = PAR_io_pipe_phv_out_data_75; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_76 = PAR_io_pipe_phv_out_data_76; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_77 = PAR_io_pipe_phv_out_data_77; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_78 = PAR_io_pipe_phv_out_data_78; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_79 = PAR_io_pipe_phv_out_data_79; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_80 = PAR_io_pipe_phv_out_data_80; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_81 = PAR_io_pipe_phv_out_data_81; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_82 = PAR_io_pipe_phv_out_data_82; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_83 = PAR_io_pipe_phv_out_data_83; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_84 = PAR_io_pipe_phv_out_data_84; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_85 = PAR_io_pipe_phv_out_data_85; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_86 = PAR_io_pipe_phv_out_data_86; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_87 = PAR_io_pipe_phv_out_data_87; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_88 = PAR_io_pipe_phv_out_data_88; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_89 = PAR_io_pipe_phv_out_data_89; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_90 = PAR_io_pipe_phv_out_data_90; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_91 = PAR_io_pipe_phv_out_data_91; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_92 = PAR_io_pipe_phv_out_data_92; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_93 = PAR_io_pipe_phv_out_data_93; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_94 = PAR_io_pipe_phv_out_data_94; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_95 = PAR_io_pipe_phv_out_data_95; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_96 = PAR_io_pipe_phv_out_data_96; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_97 = PAR_io_pipe_phv_out_data_97; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_98 = PAR_io_pipe_phv_out_data_98; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_99 = PAR_io_pipe_phv_out_data_99; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_100 = PAR_io_pipe_phv_out_data_100; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_101 = PAR_io_pipe_phv_out_data_101; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_102 = PAR_io_pipe_phv_out_data_102; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_103 = PAR_io_pipe_phv_out_data_103; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_104 = PAR_io_pipe_phv_out_data_104; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_105 = PAR_io_pipe_phv_out_data_105; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_106 = PAR_io_pipe_phv_out_data_106; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_107 = PAR_io_pipe_phv_out_data_107; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_108 = PAR_io_pipe_phv_out_data_108; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_109 = PAR_io_pipe_phv_out_data_109; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_110 = PAR_io_pipe_phv_out_data_110; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_111 = PAR_io_pipe_phv_out_data_111; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_112 = PAR_io_pipe_phv_out_data_112; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_113 = PAR_io_pipe_phv_out_data_113; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_114 = PAR_io_pipe_phv_out_data_114; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_115 = PAR_io_pipe_phv_out_data_115; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_116 = PAR_io_pipe_phv_out_data_116; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_117 = PAR_io_pipe_phv_out_data_117; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_118 = PAR_io_pipe_phv_out_data_118; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_119 = PAR_io_pipe_phv_out_data_119; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_120 = PAR_io_pipe_phv_out_data_120; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_121 = PAR_io_pipe_phv_out_data_121; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_122 = PAR_io_pipe_phv_out_data_122; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_123 = PAR_io_pipe_phv_out_data_123; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_124 = PAR_io_pipe_phv_out_data_124; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_125 = PAR_io_pipe_phv_out_data_125; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_126 = PAR_io_pipe_phv_out_data_126; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_127 = PAR_io_pipe_phv_out_data_127; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_128 = PAR_io_pipe_phv_out_data_128; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_129 = PAR_io_pipe_phv_out_data_129; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_130 = PAR_io_pipe_phv_out_data_130; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_131 = PAR_io_pipe_phv_out_data_131; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_132 = PAR_io_pipe_phv_out_data_132; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_133 = PAR_io_pipe_phv_out_data_133; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_134 = PAR_io_pipe_phv_out_data_134; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_135 = PAR_io_pipe_phv_out_data_135; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_136 = PAR_io_pipe_phv_out_data_136; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_137 = PAR_io_pipe_phv_out_data_137; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_138 = PAR_io_pipe_phv_out_data_138; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_139 = PAR_io_pipe_phv_out_data_139; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_140 = PAR_io_pipe_phv_out_data_140; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_141 = PAR_io_pipe_phv_out_data_141; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_142 = PAR_io_pipe_phv_out_data_142; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_143 = PAR_io_pipe_phv_out_data_143; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_144 = PAR_io_pipe_phv_out_data_144; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_145 = PAR_io_pipe_phv_out_data_145; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_146 = PAR_io_pipe_phv_out_data_146; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_147 = PAR_io_pipe_phv_out_data_147; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_148 = PAR_io_pipe_phv_out_data_148; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_149 = PAR_io_pipe_phv_out_data_149; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_150 = PAR_io_pipe_phv_out_data_150; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_151 = PAR_io_pipe_phv_out_data_151; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_152 = PAR_io_pipe_phv_out_data_152; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_153 = PAR_io_pipe_phv_out_data_153; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_154 = PAR_io_pipe_phv_out_data_154; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_155 = PAR_io_pipe_phv_out_data_155; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_156 = PAR_io_pipe_phv_out_data_156; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_157 = PAR_io_pipe_phv_out_data_157; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_158 = PAR_io_pipe_phv_out_data_158; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_data_159 = PAR_io_pipe_phv_out_data_159; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_0 = PAR_io_pipe_phv_out_header_0; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_1 = PAR_io_pipe_phv_out_header_1; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_2 = PAR_io_pipe_phv_out_header_2; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_3 = PAR_io_pipe_phv_out_header_3; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_4 = PAR_io_pipe_phv_out_header_4; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_5 = PAR_io_pipe_phv_out_header_5; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_6 = PAR_io_pipe_phv_out_header_6; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_7 = PAR_io_pipe_phv_out_header_7; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_8 = PAR_io_pipe_phv_out_header_8; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_9 = PAR_io_pipe_phv_out_header_9; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_10 = PAR_io_pipe_phv_out_header_10; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_11 = PAR_io_pipe_phv_out_header_11; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_12 = PAR_io_pipe_phv_out_header_12; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_13 = PAR_io_pipe_phv_out_header_13; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_14 = PAR_io_pipe_phv_out_header_14; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_header_15 = PAR_io_pipe_phv_out_header_15; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_current_state = PAR_io_pipe_phv_out_parse_current_state; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_current_offset = PAR_io_pipe_phv_out_parse_current_offset; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_parse_transition_field = PAR_io_pipe_phv_out_parse_transition_field; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_next_processor_id = PAR_io_pipe_phv_out_next_processor_id; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_next_config_id = PAR_io_pipe_phv_out_next_config_id; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_is_valid_processor = PAR_io_pipe_phv_out_is_valid_processor; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_valid = PAR_io_pipe_phv_out_valid; // @[processor.scala 20:24]
  assign MAT_io_pipe_phv_in_last = PAR_io_pipe_phv_out_last; // @[processor.scala 20:24]
  assign EXE_clock = clock;
  assign EXE_io_pipe_phv_in_data_0 = MAT_io_pipe_phv_out_data_0; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_1 = MAT_io_pipe_phv_out_data_1; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_2 = MAT_io_pipe_phv_out_data_2; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_3 = MAT_io_pipe_phv_out_data_3; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_4 = MAT_io_pipe_phv_out_data_4; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_5 = MAT_io_pipe_phv_out_data_5; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_6 = MAT_io_pipe_phv_out_data_6; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_7 = MAT_io_pipe_phv_out_data_7; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_8 = MAT_io_pipe_phv_out_data_8; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_9 = MAT_io_pipe_phv_out_data_9; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_10 = MAT_io_pipe_phv_out_data_10; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_11 = MAT_io_pipe_phv_out_data_11; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_12 = MAT_io_pipe_phv_out_data_12; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_13 = MAT_io_pipe_phv_out_data_13; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_14 = MAT_io_pipe_phv_out_data_14; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_15 = MAT_io_pipe_phv_out_data_15; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_16 = MAT_io_pipe_phv_out_data_16; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_17 = MAT_io_pipe_phv_out_data_17; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_18 = MAT_io_pipe_phv_out_data_18; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_19 = MAT_io_pipe_phv_out_data_19; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_20 = MAT_io_pipe_phv_out_data_20; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_21 = MAT_io_pipe_phv_out_data_21; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_22 = MAT_io_pipe_phv_out_data_22; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_23 = MAT_io_pipe_phv_out_data_23; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_24 = MAT_io_pipe_phv_out_data_24; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_25 = MAT_io_pipe_phv_out_data_25; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_26 = MAT_io_pipe_phv_out_data_26; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_27 = MAT_io_pipe_phv_out_data_27; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_28 = MAT_io_pipe_phv_out_data_28; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_29 = MAT_io_pipe_phv_out_data_29; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_30 = MAT_io_pipe_phv_out_data_30; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_31 = MAT_io_pipe_phv_out_data_31; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_32 = MAT_io_pipe_phv_out_data_32; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_33 = MAT_io_pipe_phv_out_data_33; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_34 = MAT_io_pipe_phv_out_data_34; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_35 = MAT_io_pipe_phv_out_data_35; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_36 = MAT_io_pipe_phv_out_data_36; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_37 = MAT_io_pipe_phv_out_data_37; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_38 = MAT_io_pipe_phv_out_data_38; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_39 = MAT_io_pipe_phv_out_data_39; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_40 = MAT_io_pipe_phv_out_data_40; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_41 = MAT_io_pipe_phv_out_data_41; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_42 = MAT_io_pipe_phv_out_data_42; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_43 = MAT_io_pipe_phv_out_data_43; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_44 = MAT_io_pipe_phv_out_data_44; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_45 = MAT_io_pipe_phv_out_data_45; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_46 = MAT_io_pipe_phv_out_data_46; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_47 = MAT_io_pipe_phv_out_data_47; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_48 = MAT_io_pipe_phv_out_data_48; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_49 = MAT_io_pipe_phv_out_data_49; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_50 = MAT_io_pipe_phv_out_data_50; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_51 = MAT_io_pipe_phv_out_data_51; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_52 = MAT_io_pipe_phv_out_data_52; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_53 = MAT_io_pipe_phv_out_data_53; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_54 = MAT_io_pipe_phv_out_data_54; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_55 = MAT_io_pipe_phv_out_data_55; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_56 = MAT_io_pipe_phv_out_data_56; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_57 = MAT_io_pipe_phv_out_data_57; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_58 = MAT_io_pipe_phv_out_data_58; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_59 = MAT_io_pipe_phv_out_data_59; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_60 = MAT_io_pipe_phv_out_data_60; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_61 = MAT_io_pipe_phv_out_data_61; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_62 = MAT_io_pipe_phv_out_data_62; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_63 = MAT_io_pipe_phv_out_data_63; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_64 = MAT_io_pipe_phv_out_data_64; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_65 = MAT_io_pipe_phv_out_data_65; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_66 = MAT_io_pipe_phv_out_data_66; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_67 = MAT_io_pipe_phv_out_data_67; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_68 = MAT_io_pipe_phv_out_data_68; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_69 = MAT_io_pipe_phv_out_data_69; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_70 = MAT_io_pipe_phv_out_data_70; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_71 = MAT_io_pipe_phv_out_data_71; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_72 = MAT_io_pipe_phv_out_data_72; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_73 = MAT_io_pipe_phv_out_data_73; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_74 = MAT_io_pipe_phv_out_data_74; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_75 = MAT_io_pipe_phv_out_data_75; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_76 = MAT_io_pipe_phv_out_data_76; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_77 = MAT_io_pipe_phv_out_data_77; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_78 = MAT_io_pipe_phv_out_data_78; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_79 = MAT_io_pipe_phv_out_data_79; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_80 = MAT_io_pipe_phv_out_data_80; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_81 = MAT_io_pipe_phv_out_data_81; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_82 = MAT_io_pipe_phv_out_data_82; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_83 = MAT_io_pipe_phv_out_data_83; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_84 = MAT_io_pipe_phv_out_data_84; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_85 = MAT_io_pipe_phv_out_data_85; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_86 = MAT_io_pipe_phv_out_data_86; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_87 = MAT_io_pipe_phv_out_data_87; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_88 = MAT_io_pipe_phv_out_data_88; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_89 = MAT_io_pipe_phv_out_data_89; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_90 = MAT_io_pipe_phv_out_data_90; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_91 = MAT_io_pipe_phv_out_data_91; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_92 = MAT_io_pipe_phv_out_data_92; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_93 = MAT_io_pipe_phv_out_data_93; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_94 = MAT_io_pipe_phv_out_data_94; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_95 = MAT_io_pipe_phv_out_data_95; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_96 = MAT_io_pipe_phv_out_data_96; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_97 = MAT_io_pipe_phv_out_data_97; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_98 = MAT_io_pipe_phv_out_data_98; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_99 = MAT_io_pipe_phv_out_data_99; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_100 = MAT_io_pipe_phv_out_data_100; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_101 = MAT_io_pipe_phv_out_data_101; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_102 = MAT_io_pipe_phv_out_data_102; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_103 = MAT_io_pipe_phv_out_data_103; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_104 = MAT_io_pipe_phv_out_data_104; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_105 = MAT_io_pipe_phv_out_data_105; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_106 = MAT_io_pipe_phv_out_data_106; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_107 = MAT_io_pipe_phv_out_data_107; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_108 = MAT_io_pipe_phv_out_data_108; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_109 = MAT_io_pipe_phv_out_data_109; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_110 = MAT_io_pipe_phv_out_data_110; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_111 = MAT_io_pipe_phv_out_data_111; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_112 = MAT_io_pipe_phv_out_data_112; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_113 = MAT_io_pipe_phv_out_data_113; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_114 = MAT_io_pipe_phv_out_data_114; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_115 = MAT_io_pipe_phv_out_data_115; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_116 = MAT_io_pipe_phv_out_data_116; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_117 = MAT_io_pipe_phv_out_data_117; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_118 = MAT_io_pipe_phv_out_data_118; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_119 = MAT_io_pipe_phv_out_data_119; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_120 = MAT_io_pipe_phv_out_data_120; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_121 = MAT_io_pipe_phv_out_data_121; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_122 = MAT_io_pipe_phv_out_data_122; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_123 = MAT_io_pipe_phv_out_data_123; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_124 = MAT_io_pipe_phv_out_data_124; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_125 = MAT_io_pipe_phv_out_data_125; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_126 = MAT_io_pipe_phv_out_data_126; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_127 = MAT_io_pipe_phv_out_data_127; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_128 = MAT_io_pipe_phv_out_data_128; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_129 = MAT_io_pipe_phv_out_data_129; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_130 = MAT_io_pipe_phv_out_data_130; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_131 = MAT_io_pipe_phv_out_data_131; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_132 = MAT_io_pipe_phv_out_data_132; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_133 = MAT_io_pipe_phv_out_data_133; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_134 = MAT_io_pipe_phv_out_data_134; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_135 = MAT_io_pipe_phv_out_data_135; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_136 = MAT_io_pipe_phv_out_data_136; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_137 = MAT_io_pipe_phv_out_data_137; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_138 = MAT_io_pipe_phv_out_data_138; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_139 = MAT_io_pipe_phv_out_data_139; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_140 = MAT_io_pipe_phv_out_data_140; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_141 = MAT_io_pipe_phv_out_data_141; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_142 = MAT_io_pipe_phv_out_data_142; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_143 = MAT_io_pipe_phv_out_data_143; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_144 = MAT_io_pipe_phv_out_data_144; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_145 = MAT_io_pipe_phv_out_data_145; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_146 = MAT_io_pipe_phv_out_data_146; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_147 = MAT_io_pipe_phv_out_data_147; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_148 = MAT_io_pipe_phv_out_data_148; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_149 = MAT_io_pipe_phv_out_data_149; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_150 = MAT_io_pipe_phv_out_data_150; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_151 = MAT_io_pipe_phv_out_data_151; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_152 = MAT_io_pipe_phv_out_data_152; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_153 = MAT_io_pipe_phv_out_data_153; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_154 = MAT_io_pipe_phv_out_data_154; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_155 = MAT_io_pipe_phv_out_data_155; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_156 = MAT_io_pipe_phv_out_data_156; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_157 = MAT_io_pipe_phv_out_data_157; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_158 = MAT_io_pipe_phv_out_data_158; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_data_159 = MAT_io_pipe_phv_out_data_159; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_0 = MAT_io_pipe_phv_out_header_0; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_1 = MAT_io_pipe_phv_out_header_1; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_2 = MAT_io_pipe_phv_out_header_2; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_3 = MAT_io_pipe_phv_out_header_3; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_4 = MAT_io_pipe_phv_out_header_4; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_5 = MAT_io_pipe_phv_out_header_5; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_6 = MAT_io_pipe_phv_out_header_6; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_7 = MAT_io_pipe_phv_out_header_7; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_8 = MAT_io_pipe_phv_out_header_8; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_9 = MAT_io_pipe_phv_out_header_9; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_10 = MAT_io_pipe_phv_out_header_10; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_11 = MAT_io_pipe_phv_out_header_11; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_12 = MAT_io_pipe_phv_out_header_12; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_13 = MAT_io_pipe_phv_out_header_13; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_14 = MAT_io_pipe_phv_out_header_14; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_header_15 = MAT_io_pipe_phv_out_header_15; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_current_state = MAT_io_pipe_phv_out_parse_current_state; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_current_offset = MAT_io_pipe_phv_out_parse_current_offset; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_parse_transition_field = MAT_io_pipe_phv_out_parse_transition_field; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_next_processor_id = MAT_io_pipe_phv_out_next_processor_id; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_next_config_id = MAT_io_pipe_phv_out_next_config_id; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_is_valid_processor = MAT_io_pipe_phv_out_is_valid_processor; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_valid = MAT_io_pipe_phv_out_valid; // @[processor.scala 24:24]
  assign EXE_io_pipe_phv_in_last = MAT_io_pipe_phv_out_last; // @[processor.scala 24:24]
endmodule
