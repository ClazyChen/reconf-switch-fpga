`include "def.svh"

module fixed_parser(
    input wire clk,
    input wire rst,
    input wire start_i,
    input wire [`BYTE_BUS] pkt_hdr_i [0:`HDR_MAX_LEN - 1],
    // output
    output reg ready_o,
    output reg [`DATA_BUS] parsed_hdrs_o [`NUM_HEADERS - 1:0]
);

    // reg
    reg [`DATA_BUS] hdr_id;
    reg [`ADDR_BUS] hdr_addr;
    reg [`HALF_BUS] next_tag;

    // parse graph
    reg [`DATA_BUS] hdr_lens [`NUM_HEADERS - 1:0];
    reg [`DATA_BUS] next_tag_starts[`NUM_HEADERS - 1:0];
    reg [`DATA_BUS] next_tag_lens[`NUM_HEADERS - 1:0];
    reg [`DATA_BUS] next_table[`NUM_HEADERS - 1:0][`NEXT_TABLE_SIZE - 1:0];

    wire [`DATA_BUS] hdr0_len;
    wire [`DATA_BUS] hdr0_tag_start;
    wire [`DATA_BUS] hdr0_tag_len;
    wire [`DATA_BUS] hdr0_next0_tag;
    wire [`DATA_BUS] hdr0_next0_hdr;
    wire [`DATA_BUS] hdr0_next1_tag;
    wire [`DATA_BUS] hdr0_next1_hdr;
    assign hdr0_len = hdr_lens[0];
    assign hdr0_tag_start = next_tag_starts[0];
    assign hdr0_tag_len = next_tag_lens[0];
    assign hdr0_next0_tag = next_table[0][0][31:16];
    assign hdr0_next0_hdr = next_table[0][0][15:0];
    assign hdr0_next1_tag = next_table[0][1][31:16];
    assign hdr0_next1_hdr = next_table[0][1][15:0];

    wire [`DATA_BUS] hdr1_len;
    wire [`DATA_BUS] hdr1_tag_start;
    wire [`DATA_BUS] hdr1_tag_len;
    wire [`DATA_BUS] hdr1_next0_tag;
    wire [`DATA_BUS] hdr1_next0_hdr;
    wire [`DATA_BUS] hdr1_next1_tag;
    wire [`DATA_BUS] hdr1_next1_hdr;
    assign hdr1_len = hdr_lens[1];
    assign hdr1_tag_start = next_tag_starts[1];
    assign hdr1_tag_len = next_tag_lens[1];
    assign hdr1_next0_tag = next_table[1][0][31:16];
    assign hdr1_next0_hdr = next_table[1][0][15:0];
    assign hdr1_next1_tag = next_table[1][1][31:16];
    assign hdr1_next1_hdr = next_table[1][1][15:0];

    wire [`DATA_BUS] hdr2_len;
    wire [`DATA_BUS] hdr2_tag_start;
    wire [`DATA_BUS] hdr2_tag_len;
    wire [`DATA_BUS] hdr2_next0_tag;
    wire [`DATA_BUS] hdr2_next0_hdr;
    wire [`DATA_BUS] hdr2_next1_tag;
    wire [`DATA_BUS] hdr2_next1_hdr;
    assign hdr2_len = hdr_lens[2];
    assign hdr2_tag_start = next_tag_starts[2];
    assign hdr2_tag_len = next_tag_lens[2];
    assign hdr2_next0_tag = next_table[2][0][31:16];
    assign hdr2_next0_hdr = next_table[2][0][15:0];
    assign hdr2_next1_tag = next_table[2][1][31:16];
    assign hdr2_next1_hdr = next_table[2][1][15:0];

    wire [`ADDR_BUS] hdr0_next0_start;
    assign hdr0_next0_start = hdr_addr + hdr0_len + next_tag_starts[hdr0_next0_hdr];
    wire [`ADDR_BUS] hdr0_next1_start;
    assign hdr0_next1_start = hdr_addr + hdr0_len + next_tag_starts[hdr0_next1_hdr];

    wire [`ADDR_BUS] hdr1_next0_start;
    assign hdr1_next0_start = hdr_addr + hdr1_len + next_tag_starts[hdr1_next0_hdr];
    wire [`ADDR_BUS] hdr1_next1_start;
    assign hdr1_next1_start = hdr_addr + hdr1_len + next_tag_starts[hdr1_next1_hdr];

    enum {
        STATE_FREE, STATE_PARSING
    } state;

    always @(posedge clk) begin
        if (rst == `TRUE) begin
            // output
            ready_o <= `FALSE;
            parsed_hdrs_o <= {`NO_HEADER, `NO_HEADER, `NO_HEADER};
            // parser
            for (int i = 2; i < `NUM_HEADERS; i++) begin
                hdr_lens[i] <= i;
                next_tag_starts[i] <= i;
                next_tag_lens[i] <= i;
                for (int j = 0; j < `NEXT_TABLE_SIZE; j++) begin
                    next_table[i][j] <= i;
                end
            end

            // ethernet header
            hdr_lens[0] <= 14;
            next_tag_starts[0] <= 12;
            next_tag_lens[0] <= 2;
            next_table[0] <= {
                {16'h0800, 16'h0001},
                `NO_NEXT_HEADER
            };

            // ip header
            hdr_lens[1] <= 20;
            next_tag_starts[1] <= 9;
            next_tag_lens[1] <= 1;
            next_table[1] <= {
                `NO_NEXT_HEADER,
                `NO_NEXT_HEADER
            };

            // reg
            hdr_id <= `NO_HEADER;
            hdr_addr <= `ZERO_ADDR;
            state <= STATE_FREE;
        end else begin
            case (state)
            STATE_FREE: begin
                if (start_i == `TRUE) begin
                    // output
                    ready_o <= `FALSE;
                    parsed_hdrs_o <= {`NO_HEADER, `NO_HEADER, `NO_HEADER};
                    // reg
                    hdr_id <= 0;
                    hdr_addr <= 0;
                    state <= STATE_PARSING;
                end
            end
            STATE_PARSING: begin
                case (hdr_id)
                0: begin
                    // parse current header offset
                    parsed_hdrs_o[0] <= hdr_addr;
                    hdr_addr <= hdr_addr + hdr0_len;
                    // match next table
                    if (next_tag == hdr0_next0_tag) begin
                        hdr_id <= hdr0_next0_hdr;
                    end else if (next_tag == hdr0_next1_tag) begin
                        hdr_id <= hdr0_next1_hdr;
                    end else begin
                        hdr_id <= `NUM_HEADERS;
                        ready_o <= `TRUE;
                        state <= STATE_FREE;
                    end
                end
                1: begin
                    parsed_hdrs_o[1] <= hdr_addr;
                    hdr_addr <= hdr_addr + hdr1_len;
                    if (next_tag == hdr1_next0_tag) begin
                        hdr_id <= hdr1_next0_hdr;
                    end else if (next_tag == hdr1_next1_tag) begin
                        hdr_id <= hdr1_next1_hdr;
                    end else begin
                        hdr_id <= `NUM_HEADERS;
                        ready_o <= `TRUE;
                        state <= STATE_FREE;
                    end
                end
                2: begin
                    parsed_hdrs_o[2] <= hdr_addr;
                    hdr_addr <= hdr_addr + hdr2_len;
                    if (next_tag == hdr2_next0_tag) begin
                        hdr_id <= hdr2_next0_hdr;
                    end else if (next_tag == hdr2_next1_tag) begin
                        hdr_id <= hdr2_next1_hdr;
                    end else begin
                        hdr_id <= `NUM_HEADERS;
                        ready_o <= `TRUE;
                        state <= STATE_FREE;
                    end
                end
                default: begin
                    hdr_id <= 0;
                end
                endcase
            end
            default: begin
                state <= STATE_FREE;
            end
            endcase
        end
    end

    always @(*) begin
        if (rst == `TRUE) begin
            next_tag = `ZERO_HALF;
        end else begin
            case (hdr_id)
            0: begin
                if (hdr0_tag_len == 1) begin
                    next_tag = {`ZERO_BYTE, pkt_hdr_i[hdr_addr + hdr0_tag_start]};
                end else begin
                    next_tag = {pkt_hdr_i[hdr_addr + hdr0_tag_start],
                                pkt_hdr_i[hdr_addr + hdr0_tag_start + 1]};
                end
            end
            1: begin
                if (hdr1_tag_len == 1) begin
                    next_tag = {`ZERO_BYTE, pkt_hdr_i[hdr_addr + hdr1_tag_start]};
                end else begin
                    next_tag = {pkt_hdr_i[hdr_addr + hdr1_tag_start],
                                pkt_hdr_i[hdr_addr + hdr1_tag_start + 1]};
                end
            end
            2: begin
                if (hdr2_tag_len == 1) begin
                    next_tag = {`ZERO_BYTE, pkt_hdr_i[hdr_addr + hdr2_tag_start]};
                end else begin
                    next_tag = {pkt_hdr_i[hdr_addr + hdr2_tag_start],
                                pkt_hdr_i[hdr_addr + hdr2_tag_start + 1]};
                end
            end
            endcase
        end
    end

endmodule
