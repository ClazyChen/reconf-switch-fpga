module PrimitiveDistributionPISA(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input  [7:0]  io_args_in_0,
  input  [7:0]  io_args_in_1,
  input  [7:0]  io_args_in_2,
  input  [7:0]  io_args_in_3,
  input  [7:0]  io_args_in_4,
  input  [7:0]  io_args_in_5,
  input  [7:0]  io_args_in_6,
  input  [31:0] io_vliw_in_0,
  input  [31:0] io_vliw_in_1,
  input  [31:0] io_vliw_in_2,
  input  [31:0] io_vliw_in_3,
  output [7:0]  io_args_out_0,
  output [7:0]  io_args_out_1,
  output [7:0]  io_args_out_2,
  output [7:0]  io_args_out_3,
  output [7:0]  io_args_out_4,
  output [7:0]  io_args_out_5,
  output [7:0]  io_args_out_6,
  output [17:0] io_vliw_out_0,
  output [17:0] io_vliw_out_1,
  output [17:0] io_vliw_out_2,
  output [17:0] io_vliw_out_3,
  output [17:0] io_vliw_out_4,
  output [17:0] io_vliw_out_5,
  output [17:0] io_vliw_out_6,
  output [17:0] io_vliw_out_7,
  output [17:0] io_vliw_out_8,
  output [17:0] io_vliw_out_9,
  output [17:0] io_vliw_out_10,
  output [17:0] io_vliw_out_11,
  output [17:0] io_vliw_out_12,
  output [17:0] io_vliw_out_13,
  output [17:0] io_vliw_out_14,
  output [17:0] io_vliw_out_15,
  output [17:0] io_vliw_out_16,
  output [17:0] io_vliw_out_17,
  output [17:0] io_vliw_out_18,
  output [17:0] io_vliw_out_19,
  output [17:0] io_vliw_out_20,
  output [17:0] io_vliw_out_21,
  output [17:0] io_vliw_out_22,
  output [17:0] io_vliw_out_23,
  output [17:0] io_vliw_out_24,
  output [17:0] io_vliw_out_25,
  output [17:0] io_vliw_out_26,
  output [17:0] io_vliw_out_27,
  output [17:0] io_vliw_out_28,
  output [17:0] io_vliw_out_29,
  output [17:0] io_vliw_out_30,
  output [17:0] io_vliw_out_31,
  output [17:0] io_vliw_out_32,
  output [17:0] io_vliw_out_33,
  output [17:0] io_vliw_out_34,
  output [17:0] io_vliw_out_35,
  output [17:0] io_vliw_out_36,
  output [17:0] io_vliw_out_37,
  output [17:0] io_vliw_out_38,
  output [17:0] io_vliw_out_39,
  output [17:0] io_vliw_out_40,
  output [17:0] io_vliw_out_41,
  output [17:0] io_vliw_out_42,
  output [17:0] io_vliw_out_43,
  output [17:0] io_vliw_out_44,
  output [17:0] io_vliw_out_45,
  output [17:0] io_vliw_out_46,
  output [17:0] io_vliw_out_47,
  output [17:0] io_vliw_out_48,
  output [17:0] io_vliw_out_49,
  output [17:0] io_vliw_out_50,
  output [17:0] io_vliw_out_51,
  output [17:0] io_vliw_out_52,
  output [17:0] io_vliw_out_53,
  output [17:0] io_vliw_out_54,
  output [17:0] io_vliw_out_55,
  output [17:0] io_vliw_out_56,
  output [17:0] io_vliw_out_57,
  output [17:0] io_vliw_out_58,
  output [17:0] io_vliw_out_59,
  output [17:0] io_vliw_out_60,
  output [17:0] io_vliw_out_61,
  output [17:0] io_vliw_out_62,
  output [17:0] io_vliw_out_63,
  output [17:0] io_vliw_out_64,
  output [17:0] io_vliw_out_65,
  output [17:0] io_vliw_out_66,
  output [17:0] io_vliw_out_67,
  output [17:0] io_vliw_out_68,
  output [17:0] io_vliw_out_69,
  output [14:0] io_nid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_1; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_2; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_3; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_4; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_5; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_6; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_7; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_8; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_9; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_10; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_11; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_12; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_13; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_14; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_15; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_16; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_17; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_18; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_19; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_20; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_21; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_22; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_23; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_24; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_25; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_26; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_27; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_28; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_29; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_30; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_31; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_32; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_33; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_34; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_35; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_36; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_37; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_38; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_39; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_40; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_41; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_42; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_43; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_44; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_45; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_46; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_47; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_48; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_49; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_50; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_51; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_52; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_53; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_54; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_55; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_56; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_57; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_58; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_59; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_60; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_61; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_62; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_63; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_64; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_65; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_66; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_67; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_68; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_69; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_70; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_71; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_72; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_73; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_74; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_75; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_76; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_77; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_78; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_79; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_80; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_81; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_82; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_83; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_84; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_85; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_86; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_87; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_88; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_89; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_90; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_91; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_92; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_93; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_94; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_95; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_96; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_97; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_98; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_99; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_100; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_101; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_102; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_103; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_104; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_105; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_106; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_107; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_108; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_109; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_110; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_111; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_112; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_113; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_114; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_115; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_116; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_117; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_118; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_119; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_120; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_121; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_122; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_123; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_124; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_125; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_126; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_127; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_128; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_129; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_130; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_131; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_132; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_133; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_134; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_135; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_136; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_137; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_138; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_139; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_140; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_141; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_142; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_143; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_144; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_145; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_146; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_147; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_148; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_149; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_150; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_151; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_152; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_153; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_154; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_155; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_156; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_157; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_158; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_159; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_160; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_161; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_162; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_163; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_164; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_165; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_166; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_167; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_168; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_169; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_170; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_171; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_172; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_173; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_174; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_175; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_176; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_177; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_178; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_179; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_180; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_181; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_182; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_183; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_184; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_185; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_186; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_187; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_188; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_189; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_190; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_191; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_192; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_193; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_194; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_195; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_196; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_197; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_198; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_199; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_200; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_201; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_202; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_203; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_204; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_205; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_206; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_207; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_208; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_209; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_210; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_211; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_212; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_213; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_214; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_215; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_216; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_217; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_218; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_219; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_220; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_221; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_222; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_223; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_224; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_225; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_226; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_227; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_228; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_229; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_230; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_231; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_232; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_233; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_234; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_235; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_236; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_237; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_238; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_239; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_240; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_241; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_242; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_243; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_244; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_245; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_246; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_247; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_248; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_249; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_250; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_251; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_252; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_253; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_254; // @[executor_pisa.scala 75:22]
  reg [7:0] phv_data_255; // @[executor_pisa.scala 75:22]
  reg [3:0] phv_next_processor_id; // @[executor_pisa.scala 75:22]
  reg  phv_next_config_id; // @[executor_pisa.scala 75:22]
  reg  phv_is_valid_processor; // @[executor_pisa.scala 75:22]
  reg [7:0] args_0; // @[executor_pisa.scala 79:23]
  reg [7:0] args_1; // @[executor_pisa.scala 79:23]
  reg [7:0] args_2; // @[executor_pisa.scala 79:23]
  reg [7:0] args_3; // @[executor_pisa.scala 79:23]
  reg [7:0] args_4; // @[executor_pisa.scala 79:23]
  reg [7:0] args_5; // @[executor_pisa.scala 79:23]
  reg [7:0] args_6; // @[executor_pisa.scala 79:23]
  reg [31:0] vliw_0; // @[executor_pisa.scala 83:23]
  reg [31:0] vliw_1; // @[executor_pisa.scala 83:23]
  reg [31:0] vliw_2; // @[executor_pisa.scala 83:23]
  reg [31:0] vliw_3; // @[executor_pisa.scala 83:23]
  wire [3:0] vliw_dis_111_hi = vliw_0[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1 = vliw_0[27:14]; // @[primitive.scala 10:44]
  wire [13:0] vliw_dis_111_lo = vliw_0[13:0]; // @[primitive.scala 11:44]
  wire [14:0] _nid_T = {1'h1,vliw_dis_111_lo}; // @[Cat.scala 30:58]
  wire [17:0] _vliw_dis_0_T = {vliw_dis_111_hi,vliw_dis_111_lo}; // @[Cat.scala 30:58]
  wire [17:0] _GEN_0 = 14'h0 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_1 = 14'h1 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_2 = 14'h2 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_3 = 14'h3 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_4 = 14'h4 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_5 = 14'h5 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_6 = 14'h6 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_7 = 14'h7 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_8 = 14'h8 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_9 = 14'h9 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_10 = 14'ha == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_11 = 14'hb == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_12 = 14'hc == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_13 = 14'hd == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_14 = 14'he == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_15 = 14'hf == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_16 = 14'h10 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_17 = 14'h11 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_18 = 14'h12 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_19 = 14'h13 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_20 = 14'h14 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_21 = 14'h15 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_22 = 14'h16 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_23 = 14'h17 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_24 = 14'h18 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_25 = 14'h19 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_26 = 14'h1a == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_27 = 14'h1b == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_28 = 14'h1c == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_29 = 14'h1d == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_30 = 14'h1e == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_31 = 14'h1f == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_32 = 14'h20 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_33 = 14'h21 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_34 = 14'h22 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_35 = 14'h23 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_36 = 14'h24 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_37 = 14'h25 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_38 = 14'h26 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_39 = 14'h27 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_40 = 14'h28 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_41 = 14'h29 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_42 = 14'h2a == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_43 = 14'h2b == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_44 = 14'h2c == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_45 = 14'h2d == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_46 = 14'h2e == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_47 = 14'h2f == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_48 = 14'h30 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_49 = 14'h31 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_50 = 14'h32 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_51 = 14'h33 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_52 = 14'h34 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_53 = 14'h35 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_54 = 14'h36 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_55 = 14'h37 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_56 = 14'h38 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_57 = 14'h39 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_58 = 14'h3a == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_59 = 14'h3b == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_60 = 14'h3c == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_61 = 14'h3d == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_62 = 14'h3e == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_63 = 14'h3f == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_64 = 14'h40 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_65 = 14'h41 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_66 = 14'h42 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_67 = 14'h43 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_68 = 14'h44 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [17:0] _GEN_69 = 14'h45 == parameter_1 ? _vliw_dis_0_T : 18'h0; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41 executor_pisa.scala 88:25]
  wire [14:0] _GEN_112 = vliw_dis_111_hi == 4'hf ? _nid_T : 15'h0; // @[executor_pisa.scala 98:52 executor_pisa.scala 99:25 executor_pisa.scala 91:13]
  wire [17:0] _GEN_113 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_0; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_114 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_1; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_115 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_2; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_116 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_3; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_117 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_4; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_118 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_5; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_119 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_6; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_120 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_7; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_121 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_8; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_122 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_9; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_123 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_10; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_124 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_11; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_125 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_12; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_126 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_13; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_127 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_14; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_128 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_15; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_129 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_16; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_130 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_17; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_131 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_18; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_132 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_19; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_133 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_20; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_134 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_21; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_135 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_22; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_136 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_23; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_137 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_24; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_138 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_25; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_139 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_26; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_140 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_27; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_141 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_28; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_142 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_29; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_143 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_30; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_144 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_31; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_145 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_32; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_146 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_33; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_147 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_34; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_148 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_35; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_149 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_36; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_150 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_37; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_151 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_38; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_152 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_39; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_153 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_40; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_154 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_41; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_155 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_42; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_156 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_43; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_157 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_44; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_158 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_45; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_159 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_46; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_160 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_47; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_161 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_48; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_162 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_49; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_163 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_50; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_164 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_51; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_165 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_52; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_166 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_53; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_167 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_54; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_168 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_55; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_169 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_56; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_170 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_57; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_171 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_58; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_172 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_59; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_173 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_60; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_174 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_61; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_175 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_62; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_176 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_63; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_177 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_64; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_178 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_65; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_179 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_66; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_180 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_67; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_181 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_68; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [17:0] _GEN_182 = vliw_dis_111_hi == 4'hf ? 18'h0 : _GEN_69; // @[executor_pisa.scala 98:52 executor_pisa.scala 88:25]
  wire [3:0] vliw_dis_111_hi_1 = vliw_1[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_1 = vliw_1[27:14]; // @[primitive.scala 10:44]
  wire [13:0] vliw_dis_111_lo_1 = vliw_1[13:0]; // @[primitive.scala 11:44]
  wire [14:0] _nid_T_1 = {1'h1,vliw_dis_111_lo_1}; // @[Cat.scala 30:58]
  wire [17:0] _vliw_dis_0_T_1 = {vliw_dis_111_hi_1,vliw_dis_111_lo_1}; // @[Cat.scala 30:58]
  wire [17:0] _GEN_225 = 14'h0 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_113; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_226 = 14'h1 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_114; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_227 = 14'h2 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_115; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_228 = 14'h3 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_116; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_229 = 14'h4 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_117; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_230 = 14'h5 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_118; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_231 = 14'h6 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_119; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_232 = 14'h7 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_120; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_233 = 14'h8 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_121; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_234 = 14'h9 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_122; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_235 = 14'ha == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_123; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_236 = 14'hb == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_124; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_237 = 14'hc == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_125; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_238 = 14'hd == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_126; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_239 = 14'he == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_127; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_240 = 14'hf == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_128; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_241 = 14'h10 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_129; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_242 = 14'h11 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_130; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_243 = 14'h12 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_131; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_244 = 14'h13 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_132; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_245 = 14'h14 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_133; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_246 = 14'h15 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_134; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_247 = 14'h16 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_135; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_248 = 14'h17 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_136; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_249 = 14'h18 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_137; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_250 = 14'h19 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_138; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_251 = 14'h1a == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_139; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_252 = 14'h1b == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_140; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_253 = 14'h1c == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_141; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_254 = 14'h1d == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_142; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_255 = 14'h1e == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_143; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_256 = 14'h1f == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_144; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_257 = 14'h20 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_145; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_258 = 14'h21 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_146; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_259 = 14'h22 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_147; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_260 = 14'h23 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_148; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_261 = 14'h24 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_149; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_262 = 14'h25 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_150; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_263 = 14'h26 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_151; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_264 = 14'h27 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_152; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_265 = 14'h28 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_153; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_266 = 14'h29 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_154; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_267 = 14'h2a == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_155; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_268 = 14'h2b == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_156; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_269 = 14'h2c == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_157; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_270 = 14'h2d == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_158; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_271 = 14'h2e == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_159; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_272 = 14'h2f == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_160; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_273 = 14'h30 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_161; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_274 = 14'h31 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_162; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_275 = 14'h32 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_163; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_276 = 14'h33 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_164; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_277 = 14'h34 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_165; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_278 = 14'h35 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_166; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_279 = 14'h36 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_167; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_280 = 14'h37 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_168; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_281 = 14'h38 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_169; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_282 = 14'h39 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_170; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_283 = 14'h3a == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_171; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_284 = 14'h3b == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_172; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_285 = 14'h3c == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_173; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_286 = 14'h3d == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_174; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_287 = 14'h3e == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_175; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_288 = 14'h3f == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_176; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_289 = 14'h40 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_177; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_290 = 14'h41 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_178; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_291 = 14'h42 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_179; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_292 = 14'h43 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_180; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_293 = 14'h44 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_181; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_294 = 14'h45 == parameter_1_1 ? _vliw_dis_0_T_1 : _GEN_182; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [14:0] _GEN_337 = vliw_dis_111_hi_1 == 4'hf ? _nid_T_1 : _GEN_112; // @[executor_pisa.scala 98:52 executor_pisa.scala 99:25]
  wire [17:0] _GEN_338 = vliw_dis_111_hi_1 == 4'hf ? _GEN_113 : _GEN_225; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_339 = vliw_dis_111_hi_1 == 4'hf ? _GEN_114 : _GEN_226; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_340 = vliw_dis_111_hi_1 == 4'hf ? _GEN_115 : _GEN_227; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_341 = vliw_dis_111_hi_1 == 4'hf ? _GEN_116 : _GEN_228; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_342 = vliw_dis_111_hi_1 == 4'hf ? _GEN_117 : _GEN_229; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_343 = vliw_dis_111_hi_1 == 4'hf ? _GEN_118 : _GEN_230; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_344 = vliw_dis_111_hi_1 == 4'hf ? _GEN_119 : _GEN_231; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_345 = vliw_dis_111_hi_1 == 4'hf ? _GEN_120 : _GEN_232; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_346 = vliw_dis_111_hi_1 == 4'hf ? _GEN_121 : _GEN_233; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_347 = vliw_dis_111_hi_1 == 4'hf ? _GEN_122 : _GEN_234; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_348 = vliw_dis_111_hi_1 == 4'hf ? _GEN_123 : _GEN_235; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_349 = vliw_dis_111_hi_1 == 4'hf ? _GEN_124 : _GEN_236; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_350 = vliw_dis_111_hi_1 == 4'hf ? _GEN_125 : _GEN_237; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_351 = vliw_dis_111_hi_1 == 4'hf ? _GEN_126 : _GEN_238; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_352 = vliw_dis_111_hi_1 == 4'hf ? _GEN_127 : _GEN_239; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_353 = vliw_dis_111_hi_1 == 4'hf ? _GEN_128 : _GEN_240; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_354 = vliw_dis_111_hi_1 == 4'hf ? _GEN_129 : _GEN_241; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_355 = vliw_dis_111_hi_1 == 4'hf ? _GEN_130 : _GEN_242; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_356 = vliw_dis_111_hi_1 == 4'hf ? _GEN_131 : _GEN_243; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_357 = vliw_dis_111_hi_1 == 4'hf ? _GEN_132 : _GEN_244; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_358 = vliw_dis_111_hi_1 == 4'hf ? _GEN_133 : _GEN_245; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_359 = vliw_dis_111_hi_1 == 4'hf ? _GEN_134 : _GEN_246; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_360 = vliw_dis_111_hi_1 == 4'hf ? _GEN_135 : _GEN_247; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_361 = vliw_dis_111_hi_1 == 4'hf ? _GEN_136 : _GEN_248; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_362 = vliw_dis_111_hi_1 == 4'hf ? _GEN_137 : _GEN_249; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_363 = vliw_dis_111_hi_1 == 4'hf ? _GEN_138 : _GEN_250; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_364 = vliw_dis_111_hi_1 == 4'hf ? _GEN_139 : _GEN_251; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_365 = vliw_dis_111_hi_1 == 4'hf ? _GEN_140 : _GEN_252; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_366 = vliw_dis_111_hi_1 == 4'hf ? _GEN_141 : _GEN_253; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_367 = vliw_dis_111_hi_1 == 4'hf ? _GEN_142 : _GEN_254; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_368 = vliw_dis_111_hi_1 == 4'hf ? _GEN_143 : _GEN_255; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_369 = vliw_dis_111_hi_1 == 4'hf ? _GEN_144 : _GEN_256; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_370 = vliw_dis_111_hi_1 == 4'hf ? _GEN_145 : _GEN_257; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_371 = vliw_dis_111_hi_1 == 4'hf ? _GEN_146 : _GEN_258; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_372 = vliw_dis_111_hi_1 == 4'hf ? _GEN_147 : _GEN_259; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_373 = vliw_dis_111_hi_1 == 4'hf ? _GEN_148 : _GEN_260; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_374 = vliw_dis_111_hi_1 == 4'hf ? _GEN_149 : _GEN_261; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_375 = vliw_dis_111_hi_1 == 4'hf ? _GEN_150 : _GEN_262; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_376 = vliw_dis_111_hi_1 == 4'hf ? _GEN_151 : _GEN_263; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_377 = vliw_dis_111_hi_1 == 4'hf ? _GEN_152 : _GEN_264; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_378 = vliw_dis_111_hi_1 == 4'hf ? _GEN_153 : _GEN_265; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_379 = vliw_dis_111_hi_1 == 4'hf ? _GEN_154 : _GEN_266; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_380 = vliw_dis_111_hi_1 == 4'hf ? _GEN_155 : _GEN_267; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_381 = vliw_dis_111_hi_1 == 4'hf ? _GEN_156 : _GEN_268; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_382 = vliw_dis_111_hi_1 == 4'hf ? _GEN_157 : _GEN_269; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_383 = vliw_dis_111_hi_1 == 4'hf ? _GEN_158 : _GEN_270; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_384 = vliw_dis_111_hi_1 == 4'hf ? _GEN_159 : _GEN_271; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_385 = vliw_dis_111_hi_1 == 4'hf ? _GEN_160 : _GEN_272; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_386 = vliw_dis_111_hi_1 == 4'hf ? _GEN_161 : _GEN_273; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_387 = vliw_dis_111_hi_1 == 4'hf ? _GEN_162 : _GEN_274; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_388 = vliw_dis_111_hi_1 == 4'hf ? _GEN_163 : _GEN_275; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_389 = vliw_dis_111_hi_1 == 4'hf ? _GEN_164 : _GEN_276; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_390 = vliw_dis_111_hi_1 == 4'hf ? _GEN_165 : _GEN_277; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_391 = vliw_dis_111_hi_1 == 4'hf ? _GEN_166 : _GEN_278; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_392 = vliw_dis_111_hi_1 == 4'hf ? _GEN_167 : _GEN_279; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_393 = vliw_dis_111_hi_1 == 4'hf ? _GEN_168 : _GEN_280; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_394 = vliw_dis_111_hi_1 == 4'hf ? _GEN_169 : _GEN_281; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_395 = vliw_dis_111_hi_1 == 4'hf ? _GEN_170 : _GEN_282; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_396 = vliw_dis_111_hi_1 == 4'hf ? _GEN_171 : _GEN_283; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_397 = vliw_dis_111_hi_1 == 4'hf ? _GEN_172 : _GEN_284; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_398 = vliw_dis_111_hi_1 == 4'hf ? _GEN_173 : _GEN_285; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_399 = vliw_dis_111_hi_1 == 4'hf ? _GEN_174 : _GEN_286; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_400 = vliw_dis_111_hi_1 == 4'hf ? _GEN_175 : _GEN_287; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_401 = vliw_dis_111_hi_1 == 4'hf ? _GEN_176 : _GEN_288; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_402 = vliw_dis_111_hi_1 == 4'hf ? _GEN_177 : _GEN_289; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_403 = vliw_dis_111_hi_1 == 4'hf ? _GEN_178 : _GEN_290; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_404 = vliw_dis_111_hi_1 == 4'hf ? _GEN_179 : _GEN_291; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_405 = vliw_dis_111_hi_1 == 4'hf ? _GEN_180 : _GEN_292; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_406 = vliw_dis_111_hi_1 == 4'hf ? _GEN_181 : _GEN_293; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_407 = vliw_dis_111_hi_1 == 4'hf ? _GEN_182 : _GEN_294; // @[executor_pisa.scala 98:52]
  wire [3:0] vliw_dis_111_hi_2 = vliw_2[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_2 = vliw_2[27:14]; // @[primitive.scala 10:44]
  wire [13:0] vliw_dis_111_lo_2 = vliw_2[13:0]; // @[primitive.scala 11:44]
  wire [14:0] _nid_T_2 = {1'h1,vliw_dis_111_lo_2}; // @[Cat.scala 30:58]
  wire [17:0] _vliw_dis_0_T_2 = {vliw_dis_111_hi_2,vliw_dis_111_lo_2}; // @[Cat.scala 30:58]
  wire [17:0] _GEN_450 = 14'h0 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_338; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_451 = 14'h1 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_339; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_452 = 14'h2 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_340; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_453 = 14'h3 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_341; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_454 = 14'h4 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_342; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_455 = 14'h5 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_343; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_456 = 14'h6 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_344; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_457 = 14'h7 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_345; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_458 = 14'h8 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_346; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_459 = 14'h9 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_347; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_460 = 14'ha == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_348; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_461 = 14'hb == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_349; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_462 = 14'hc == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_350; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_463 = 14'hd == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_351; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_464 = 14'he == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_352; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_465 = 14'hf == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_353; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_466 = 14'h10 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_354; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_467 = 14'h11 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_355; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_468 = 14'h12 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_356; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_469 = 14'h13 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_357; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_470 = 14'h14 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_358; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_471 = 14'h15 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_359; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_472 = 14'h16 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_360; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_473 = 14'h17 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_361; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_474 = 14'h18 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_362; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_475 = 14'h19 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_363; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_476 = 14'h1a == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_364; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_477 = 14'h1b == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_365; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_478 = 14'h1c == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_366; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_479 = 14'h1d == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_367; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_480 = 14'h1e == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_368; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_481 = 14'h1f == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_369; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_482 = 14'h20 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_370; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_483 = 14'h21 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_371; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_484 = 14'h22 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_372; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_485 = 14'h23 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_373; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_486 = 14'h24 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_374; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_487 = 14'h25 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_375; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_488 = 14'h26 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_376; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_489 = 14'h27 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_377; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_490 = 14'h28 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_378; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_491 = 14'h29 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_379; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_492 = 14'h2a == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_380; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_493 = 14'h2b == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_381; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_494 = 14'h2c == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_382; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_495 = 14'h2d == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_383; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_496 = 14'h2e == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_384; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_497 = 14'h2f == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_385; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_498 = 14'h30 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_386; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_499 = 14'h31 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_387; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_500 = 14'h32 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_388; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_501 = 14'h33 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_389; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_502 = 14'h34 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_390; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_503 = 14'h35 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_391; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_504 = 14'h36 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_392; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_505 = 14'h37 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_393; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_506 = 14'h38 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_394; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_507 = 14'h39 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_395; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_508 = 14'h3a == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_396; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_509 = 14'h3b == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_397; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_510 = 14'h3c == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_398; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_511 = 14'h3d == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_399; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_512 = 14'h3e == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_400; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_513 = 14'h3f == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_401; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_514 = 14'h40 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_402; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_515 = 14'h41 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_403; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_516 = 14'h42 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_404; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_517 = 14'h43 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_405; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_518 = 14'h44 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_406; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_519 = 14'h45 == parameter_1_2 ? _vliw_dis_0_T_2 : _GEN_407; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [14:0] _GEN_562 = vliw_dis_111_hi_2 == 4'hf ? _nid_T_2 : _GEN_337; // @[executor_pisa.scala 98:52 executor_pisa.scala 99:25]
  wire [17:0] _GEN_563 = vliw_dis_111_hi_2 == 4'hf ? _GEN_338 : _GEN_450; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_564 = vliw_dis_111_hi_2 == 4'hf ? _GEN_339 : _GEN_451; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_565 = vliw_dis_111_hi_2 == 4'hf ? _GEN_340 : _GEN_452; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_566 = vliw_dis_111_hi_2 == 4'hf ? _GEN_341 : _GEN_453; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_567 = vliw_dis_111_hi_2 == 4'hf ? _GEN_342 : _GEN_454; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_568 = vliw_dis_111_hi_2 == 4'hf ? _GEN_343 : _GEN_455; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_569 = vliw_dis_111_hi_2 == 4'hf ? _GEN_344 : _GEN_456; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_570 = vliw_dis_111_hi_2 == 4'hf ? _GEN_345 : _GEN_457; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_571 = vliw_dis_111_hi_2 == 4'hf ? _GEN_346 : _GEN_458; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_572 = vliw_dis_111_hi_2 == 4'hf ? _GEN_347 : _GEN_459; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_573 = vliw_dis_111_hi_2 == 4'hf ? _GEN_348 : _GEN_460; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_574 = vliw_dis_111_hi_2 == 4'hf ? _GEN_349 : _GEN_461; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_575 = vliw_dis_111_hi_2 == 4'hf ? _GEN_350 : _GEN_462; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_576 = vliw_dis_111_hi_2 == 4'hf ? _GEN_351 : _GEN_463; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_577 = vliw_dis_111_hi_2 == 4'hf ? _GEN_352 : _GEN_464; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_578 = vliw_dis_111_hi_2 == 4'hf ? _GEN_353 : _GEN_465; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_579 = vliw_dis_111_hi_2 == 4'hf ? _GEN_354 : _GEN_466; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_580 = vliw_dis_111_hi_2 == 4'hf ? _GEN_355 : _GEN_467; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_581 = vliw_dis_111_hi_2 == 4'hf ? _GEN_356 : _GEN_468; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_582 = vliw_dis_111_hi_2 == 4'hf ? _GEN_357 : _GEN_469; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_583 = vliw_dis_111_hi_2 == 4'hf ? _GEN_358 : _GEN_470; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_584 = vliw_dis_111_hi_2 == 4'hf ? _GEN_359 : _GEN_471; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_585 = vliw_dis_111_hi_2 == 4'hf ? _GEN_360 : _GEN_472; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_586 = vliw_dis_111_hi_2 == 4'hf ? _GEN_361 : _GEN_473; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_587 = vliw_dis_111_hi_2 == 4'hf ? _GEN_362 : _GEN_474; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_588 = vliw_dis_111_hi_2 == 4'hf ? _GEN_363 : _GEN_475; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_589 = vliw_dis_111_hi_2 == 4'hf ? _GEN_364 : _GEN_476; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_590 = vliw_dis_111_hi_2 == 4'hf ? _GEN_365 : _GEN_477; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_591 = vliw_dis_111_hi_2 == 4'hf ? _GEN_366 : _GEN_478; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_592 = vliw_dis_111_hi_2 == 4'hf ? _GEN_367 : _GEN_479; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_593 = vliw_dis_111_hi_2 == 4'hf ? _GEN_368 : _GEN_480; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_594 = vliw_dis_111_hi_2 == 4'hf ? _GEN_369 : _GEN_481; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_595 = vliw_dis_111_hi_2 == 4'hf ? _GEN_370 : _GEN_482; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_596 = vliw_dis_111_hi_2 == 4'hf ? _GEN_371 : _GEN_483; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_597 = vliw_dis_111_hi_2 == 4'hf ? _GEN_372 : _GEN_484; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_598 = vliw_dis_111_hi_2 == 4'hf ? _GEN_373 : _GEN_485; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_599 = vliw_dis_111_hi_2 == 4'hf ? _GEN_374 : _GEN_486; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_600 = vliw_dis_111_hi_2 == 4'hf ? _GEN_375 : _GEN_487; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_601 = vliw_dis_111_hi_2 == 4'hf ? _GEN_376 : _GEN_488; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_602 = vliw_dis_111_hi_2 == 4'hf ? _GEN_377 : _GEN_489; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_603 = vliw_dis_111_hi_2 == 4'hf ? _GEN_378 : _GEN_490; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_604 = vliw_dis_111_hi_2 == 4'hf ? _GEN_379 : _GEN_491; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_605 = vliw_dis_111_hi_2 == 4'hf ? _GEN_380 : _GEN_492; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_606 = vliw_dis_111_hi_2 == 4'hf ? _GEN_381 : _GEN_493; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_607 = vliw_dis_111_hi_2 == 4'hf ? _GEN_382 : _GEN_494; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_608 = vliw_dis_111_hi_2 == 4'hf ? _GEN_383 : _GEN_495; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_609 = vliw_dis_111_hi_2 == 4'hf ? _GEN_384 : _GEN_496; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_610 = vliw_dis_111_hi_2 == 4'hf ? _GEN_385 : _GEN_497; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_611 = vliw_dis_111_hi_2 == 4'hf ? _GEN_386 : _GEN_498; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_612 = vliw_dis_111_hi_2 == 4'hf ? _GEN_387 : _GEN_499; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_613 = vliw_dis_111_hi_2 == 4'hf ? _GEN_388 : _GEN_500; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_614 = vliw_dis_111_hi_2 == 4'hf ? _GEN_389 : _GEN_501; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_615 = vliw_dis_111_hi_2 == 4'hf ? _GEN_390 : _GEN_502; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_616 = vliw_dis_111_hi_2 == 4'hf ? _GEN_391 : _GEN_503; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_617 = vliw_dis_111_hi_2 == 4'hf ? _GEN_392 : _GEN_504; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_618 = vliw_dis_111_hi_2 == 4'hf ? _GEN_393 : _GEN_505; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_619 = vliw_dis_111_hi_2 == 4'hf ? _GEN_394 : _GEN_506; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_620 = vliw_dis_111_hi_2 == 4'hf ? _GEN_395 : _GEN_507; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_621 = vliw_dis_111_hi_2 == 4'hf ? _GEN_396 : _GEN_508; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_622 = vliw_dis_111_hi_2 == 4'hf ? _GEN_397 : _GEN_509; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_623 = vliw_dis_111_hi_2 == 4'hf ? _GEN_398 : _GEN_510; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_624 = vliw_dis_111_hi_2 == 4'hf ? _GEN_399 : _GEN_511; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_625 = vliw_dis_111_hi_2 == 4'hf ? _GEN_400 : _GEN_512; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_626 = vliw_dis_111_hi_2 == 4'hf ? _GEN_401 : _GEN_513; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_627 = vliw_dis_111_hi_2 == 4'hf ? _GEN_402 : _GEN_514; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_628 = vliw_dis_111_hi_2 == 4'hf ? _GEN_403 : _GEN_515; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_629 = vliw_dis_111_hi_2 == 4'hf ? _GEN_404 : _GEN_516; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_630 = vliw_dis_111_hi_2 == 4'hf ? _GEN_405 : _GEN_517; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_631 = vliw_dis_111_hi_2 == 4'hf ? _GEN_406 : _GEN_518; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_632 = vliw_dis_111_hi_2 == 4'hf ? _GEN_407 : _GEN_519; // @[executor_pisa.scala 98:52]
  wire [3:0] vliw_dis_111_hi_3 = vliw_3[31:28]; // @[primitive.scala 9:44]
  wire [13:0] parameter_1_3 = vliw_3[27:14]; // @[primitive.scala 10:44]
  wire [13:0] vliw_dis_111_lo_3 = vliw_3[13:0]; // @[primitive.scala 11:44]
  wire [14:0] _nid_T_3 = {1'h1,vliw_dis_111_lo_3}; // @[Cat.scala 30:58]
  wire [17:0] _vliw_dis_0_T_3 = {vliw_dis_111_hi_3,vliw_dis_111_lo_3}; // @[Cat.scala 30:58]
  wire [17:0] _GEN_675 = 14'h0 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_563; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_676 = 14'h1 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_564; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_677 = 14'h2 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_565; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_678 = 14'h3 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_566; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_679 = 14'h4 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_567; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_680 = 14'h5 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_568; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_681 = 14'h6 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_569; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_682 = 14'h7 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_570; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_683 = 14'h8 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_571; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_684 = 14'h9 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_572; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_685 = 14'ha == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_573; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_686 = 14'hb == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_574; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_687 = 14'hc == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_575; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_688 = 14'hd == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_576; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_689 = 14'he == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_577; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_690 = 14'hf == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_578; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_691 = 14'h10 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_579; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_692 = 14'h11 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_580; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_693 = 14'h12 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_581; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_694 = 14'h13 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_582; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_695 = 14'h14 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_583; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_696 = 14'h15 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_584; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_697 = 14'h16 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_585; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_698 = 14'h17 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_586; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_699 = 14'h18 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_587; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_700 = 14'h19 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_588; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_701 = 14'h1a == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_589; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_702 = 14'h1b == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_590; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_703 = 14'h1c == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_591; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_704 = 14'h1d == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_592; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_705 = 14'h1e == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_593; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_706 = 14'h1f == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_594; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_707 = 14'h20 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_595; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_708 = 14'h21 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_596; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_709 = 14'h22 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_597; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_710 = 14'h23 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_598; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_711 = 14'h24 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_599; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_712 = 14'h25 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_600; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_713 = 14'h26 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_601; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_714 = 14'h27 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_602; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_715 = 14'h28 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_603; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_716 = 14'h29 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_604; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_717 = 14'h2a == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_605; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_718 = 14'h2b == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_606; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_719 = 14'h2c == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_607; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_720 = 14'h2d == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_608; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_721 = 14'h2e == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_609; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_722 = 14'h2f == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_610; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_723 = 14'h30 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_611; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_724 = 14'h31 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_612; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_725 = 14'h32 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_613; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_726 = 14'h33 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_614; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_727 = 14'h34 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_615; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_728 = 14'h35 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_616; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_729 = 14'h36 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_617; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_730 = 14'h37 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_618; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_731 = 14'h38 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_619; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_732 = 14'h39 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_620; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_733 = 14'h3a == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_621; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_734 = 14'h3b == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_622; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_735 = 14'h3c == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_623; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_736 = 14'h3d == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_624; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_737 = 14'h3e == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_625; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_738 = 14'h3f == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_626; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_739 = 14'h40 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_627; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_740 = 14'h41 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_628; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_741 = 14'h42 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_629; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_742 = 14'h43 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_630; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_743 = 14'h44 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_631; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [17:0] _GEN_744 = 14'h45 == parameter_1_3 ? _vliw_dis_0_T_3 : _GEN_632; // @[executor_pisa.scala 102:52 executor_pisa.scala 103:41]
  wire [14:0] _GEN_787 = vliw_dis_111_hi_3 == 4'hf ? _nid_T_3 : _GEN_562; // @[executor_pisa.scala 98:52 executor_pisa.scala 99:25]
  wire [17:0] _GEN_788 = vliw_dis_111_hi_3 == 4'hf ? _GEN_563 : _GEN_675; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_789 = vliw_dis_111_hi_3 == 4'hf ? _GEN_564 : _GEN_676; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_790 = vliw_dis_111_hi_3 == 4'hf ? _GEN_565 : _GEN_677; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_791 = vliw_dis_111_hi_3 == 4'hf ? _GEN_566 : _GEN_678; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_792 = vliw_dis_111_hi_3 == 4'hf ? _GEN_567 : _GEN_679; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_793 = vliw_dis_111_hi_3 == 4'hf ? _GEN_568 : _GEN_680; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_794 = vliw_dis_111_hi_3 == 4'hf ? _GEN_569 : _GEN_681; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_795 = vliw_dis_111_hi_3 == 4'hf ? _GEN_570 : _GEN_682; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_796 = vliw_dis_111_hi_3 == 4'hf ? _GEN_571 : _GEN_683; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_797 = vliw_dis_111_hi_3 == 4'hf ? _GEN_572 : _GEN_684; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_798 = vliw_dis_111_hi_3 == 4'hf ? _GEN_573 : _GEN_685; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_799 = vliw_dis_111_hi_3 == 4'hf ? _GEN_574 : _GEN_686; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_800 = vliw_dis_111_hi_3 == 4'hf ? _GEN_575 : _GEN_687; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_801 = vliw_dis_111_hi_3 == 4'hf ? _GEN_576 : _GEN_688; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_802 = vliw_dis_111_hi_3 == 4'hf ? _GEN_577 : _GEN_689; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_803 = vliw_dis_111_hi_3 == 4'hf ? _GEN_578 : _GEN_690; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_804 = vliw_dis_111_hi_3 == 4'hf ? _GEN_579 : _GEN_691; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_805 = vliw_dis_111_hi_3 == 4'hf ? _GEN_580 : _GEN_692; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_806 = vliw_dis_111_hi_3 == 4'hf ? _GEN_581 : _GEN_693; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_807 = vliw_dis_111_hi_3 == 4'hf ? _GEN_582 : _GEN_694; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_808 = vliw_dis_111_hi_3 == 4'hf ? _GEN_583 : _GEN_695; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_809 = vliw_dis_111_hi_3 == 4'hf ? _GEN_584 : _GEN_696; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_810 = vliw_dis_111_hi_3 == 4'hf ? _GEN_585 : _GEN_697; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_811 = vliw_dis_111_hi_3 == 4'hf ? _GEN_586 : _GEN_698; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_812 = vliw_dis_111_hi_3 == 4'hf ? _GEN_587 : _GEN_699; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_813 = vliw_dis_111_hi_3 == 4'hf ? _GEN_588 : _GEN_700; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_814 = vliw_dis_111_hi_3 == 4'hf ? _GEN_589 : _GEN_701; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_815 = vliw_dis_111_hi_3 == 4'hf ? _GEN_590 : _GEN_702; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_816 = vliw_dis_111_hi_3 == 4'hf ? _GEN_591 : _GEN_703; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_817 = vliw_dis_111_hi_3 == 4'hf ? _GEN_592 : _GEN_704; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_818 = vliw_dis_111_hi_3 == 4'hf ? _GEN_593 : _GEN_705; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_819 = vliw_dis_111_hi_3 == 4'hf ? _GEN_594 : _GEN_706; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_820 = vliw_dis_111_hi_3 == 4'hf ? _GEN_595 : _GEN_707; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_821 = vliw_dis_111_hi_3 == 4'hf ? _GEN_596 : _GEN_708; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_822 = vliw_dis_111_hi_3 == 4'hf ? _GEN_597 : _GEN_709; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_823 = vliw_dis_111_hi_3 == 4'hf ? _GEN_598 : _GEN_710; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_824 = vliw_dis_111_hi_3 == 4'hf ? _GEN_599 : _GEN_711; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_825 = vliw_dis_111_hi_3 == 4'hf ? _GEN_600 : _GEN_712; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_826 = vliw_dis_111_hi_3 == 4'hf ? _GEN_601 : _GEN_713; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_827 = vliw_dis_111_hi_3 == 4'hf ? _GEN_602 : _GEN_714; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_828 = vliw_dis_111_hi_3 == 4'hf ? _GEN_603 : _GEN_715; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_829 = vliw_dis_111_hi_3 == 4'hf ? _GEN_604 : _GEN_716; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_830 = vliw_dis_111_hi_3 == 4'hf ? _GEN_605 : _GEN_717; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_831 = vliw_dis_111_hi_3 == 4'hf ? _GEN_606 : _GEN_718; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_832 = vliw_dis_111_hi_3 == 4'hf ? _GEN_607 : _GEN_719; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_833 = vliw_dis_111_hi_3 == 4'hf ? _GEN_608 : _GEN_720; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_834 = vliw_dis_111_hi_3 == 4'hf ? _GEN_609 : _GEN_721; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_835 = vliw_dis_111_hi_3 == 4'hf ? _GEN_610 : _GEN_722; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_836 = vliw_dis_111_hi_3 == 4'hf ? _GEN_611 : _GEN_723; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_837 = vliw_dis_111_hi_3 == 4'hf ? _GEN_612 : _GEN_724; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_838 = vliw_dis_111_hi_3 == 4'hf ? _GEN_613 : _GEN_725; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_839 = vliw_dis_111_hi_3 == 4'hf ? _GEN_614 : _GEN_726; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_840 = vliw_dis_111_hi_3 == 4'hf ? _GEN_615 : _GEN_727; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_841 = vliw_dis_111_hi_3 == 4'hf ? _GEN_616 : _GEN_728; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_842 = vliw_dis_111_hi_3 == 4'hf ? _GEN_617 : _GEN_729; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_843 = vliw_dis_111_hi_3 == 4'hf ? _GEN_618 : _GEN_730; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_844 = vliw_dis_111_hi_3 == 4'hf ? _GEN_619 : _GEN_731; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_845 = vliw_dis_111_hi_3 == 4'hf ? _GEN_620 : _GEN_732; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_846 = vliw_dis_111_hi_3 == 4'hf ? _GEN_621 : _GEN_733; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_847 = vliw_dis_111_hi_3 == 4'hf ? _GEN_622 : _GEN_734; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_848 = vliw_dis_111_hi_3 == 4'hf ? _GEN_623 : _GEN_735; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_849 = vliw_dis_111_hi_3 == 4'hf ? _GEN_624 : _GEN_736; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_850 = vliw_dis_111_hi_3 == 4'hf ? _GEN_625 : _GEN_737; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_851 = vliw_dis_111_hi_3 == 4'hf ? _GEN_626 : _GEN_738; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_852 = vliw_dis_111_hi_3 == 4'hf ? _GEN_627 : _GEN_739; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_853 = vliw_dis_111_hi_3 == 4'hf ? _GEN_628 : _GEN_740; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_854 = vliw_dis_111_hi_3 == 4'hf ? _GEN_629 : _GEN_741; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_855 = vliw_dis_111_hi_3 == 4'hf ? _GEN_630 : _GEN_742; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_856 = vliw_dis_111_hi_3 == 4'hf ? _GEN_631 : _GEN_743; // @[executor_pisa.scala 98:52]
  wire [17:0] _GEN_857 = vliw_dis_111_hi_3 == 4'hf ? _GEN_632 : _GEN_744; // @[executor_pisa.scala 98:52]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[executor_pisa.scala 77:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[executor_pisa.scala 77:25]
  assign io_args_out_0 = args_0; // @[executor_pisa.scala 81:21]
  assign io_args_out_1 = args_1; // @[executor_pisa.scala 81:21]
  assign io_args_out_2 = args_2; // @[executor_pisa.scala 81:21]
  assign io_args_out_3 = args_3; // @[executor_pisa.scala 81:21]
  assign io_args_out_4 = args_4; // @[executor_pisa.scala 81:21]
  assign io_args_out_5 = args_5; // @[executor_pisa.scala 81:21]
  assign io_args_out_6 = args_6; // @[executor_pisa.scala 81:21]
  assign io_vliw_out_0 = phv_is_valid_processor ? _GEN_788 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_1 = phv_is_valid_processor ? _GEN_789 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_2 = phv_is_valid_processor ? _GEN_790 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_3 = phv_is_valid_processor ? _GEN_791 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_4 = phv_is_valid_processor ? _GEN_792 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_5 = phv_is_valid_processor ? _GEN_793 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_6 = phv_is_valid_processor ? _GEN_794 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_7 = phv_is_valid_processor ? _GEN_795 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_8 = phv_is_valid_processor ? _GEN_796 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_9 = phv_is_valid_processor ? _GEN_797 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_10 = phv_is_valid_processor ? _GEN_798 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_11 = phv_is_valid_processor ? _GEN_799 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_12 = phv_is_valid_processor ? _GEN_800 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_13 = phv_is_valid_processor ? _GEN_801 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_14 = phv_is_valid_processor ? _GEN_802 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_15 = phv_is_valid_processor ? _GEN_803 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_16 = phv_is_valid_processor ? _GEN_804 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_17 = phv_is_valid_processor ? _GEN_805 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_18 = phv_is_valid_processor ? _GEN_806 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_19 = phv_is_valid_processor ? _GEN_807 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_20 = phv_is_valid_processor ? _GEN_808 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_21 = phv_is_valid_processor ? _GEN_809 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_22 = phv_is_valid_processor ? _GEN_810 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_23 = phv_is_valid_processor ? _GEN_811 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_24 = phv_is_valid_processor ? _GEN_812 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_25 = phv_is_valid_processor ? _GEN_813 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_26 = phv_is_valid_processor ? _GEN_814 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_27 = phv_is_valid_processor ? _GEN_815 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_28 = phv_is_valid_processor ? _GEN_816 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_29 = phv_is_valid_processor ? _GEN_817 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_30 = phv_is_valid_processor ? _GEN_818 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_31 = phv_is_valid_processor ? _GEN_819 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_32 = phv_is_valid_processor ? _GEN_820 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_33 = phv_is_valid_processor ? _GEN_821 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_34 = phv_is_valid_processor ? _GEN_822 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_35 = phv_is_valid_processor ? _GEN_823 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_36 = phv_is_valid_processor ? _GEN_824 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_37 = phv_is_valid_processor ? _GEN_825 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_38 = phv_is_valid_processor ? _GEN_826 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_39 = phv_is_valid_processor ? _GEN_827 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_40 = phv_is_valid_processor ? _GEN_828 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_41 = phv_is_valid_processor ? _GEN_829 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_42 = phv_is_valid_processor ? _GEN_830 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_43 = phv_is_valid_processor ? _GEN_831 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_44 = phv_is_valid_processor ? _GEN_832 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_45 = phv_is_valid_processor ? _GEN_833 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_46 = phv_is_valid_processor ? _GEN_834 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_47 = phv_is_valid_processor ? _GEN_835 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_48 = phv_is_valid_processor ? _GEN_836 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_49 = phv_is_valid_processor ? _GEN_837 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_50 = phv_is_valid_processor ? _GEN_838 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_51 = phv_is_valid_processor ? _GEN_839 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_52 = phv_is_valid_processor ? _GEN_840 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_53 = phv_is_valid_processor ? _GEN_841 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_54 = phv_is_valid_processor ? _GEN_842 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_55 = phv_is_valid_processor ? _GEN_843 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_56 = phv_is_valid_processor ? _GEN_844 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_57 = phv_is_valid_processor ? _GEN_845 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_58 = phv_is_valid_processor ? _GEN_846 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_59 = phv_is_valid_processor ? _GEN_847 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_60 = phv_is_valid_processor ? _GEN_848 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_61 = phv_is_valid_processor ? _GEN_849 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_62 = phv_is_valid_processor ? _GEN_850 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_63 = phv_is_valid_processor ? _GEN_851 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_64 = phv_is_valid_processor ? _GEN_852 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_65 = phv_is_valid_processor ? _GEN_853 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_66 = phv_is_valid_processor ? _GEN_854 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_67 = phv_is_valid_processor ? _GEN_855 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_68 = phv_is_valid_processor ? _GEN_856 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_vliw_out_69 = phv_is_valid_processor ? _GEN_857 : 18'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 88:25]
  assign io_nid_out = phv_is_valid_processor ? _GEN_787 : 15'h0; // @[executor_pisa.scala 93:39 executor_pisa.scala 91:13]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[executor_pisa.scala 76:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[executor_pisa.scala 76:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[executor_pisa.scala 76:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[executor_pisa.scala 76:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[executor_pisa.scala 76:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[executor_pisa.scala 76:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[executor_pisa.scala 76:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[executor_pisa.scala 76:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[executor_pisa.scala 76:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[executor_pisa.scala 76:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[executor_pisa.scala 76:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[executor_pisa.scala 76:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[executor_pisa.scala 76:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[executor_pisa.scala 76:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[executor_pisa.scala 76:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[executor_pisa.scala 76:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[executor_pisa.scala 76:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[executor_pisa.scala 76:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[executor_pisa.scala 76:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[executor_pisa.scala 76:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[executor_pisa.scala 76:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[executor_pisa.scala 76:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[executor_pisa.scala 76:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[executor_pisa.scala 76:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[executor_pisa.scala 76:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[executor_pisa.scala 76:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[executor_pisa.scala 76:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[executor_pisa.scala 76:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[executor_pisa.scala 76:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[executor_pisa.scala 76:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[executor_pisa.scala 76:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[executor_pisa.scala 76:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[executor_pisa.scala 76:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[executor_pisa.scala 76:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[executor_pisa.scala 76:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[executor_pisa.scala 76:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[executor_pisa.scala 76:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[executor_pisa.scala 76:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[executor_pisa.scala 76:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[executor_pisa.scala 76:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[executor_pisa.scala 76:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[executor_pisa.scala 76:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[executor_pisa.scala 76:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[executor_pisa.scala 76:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[executor_pisa.scala 76:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[executor_pisa.scala 76:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[executor_pisa.scala 76:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[executor_pisa.scala 76:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[executor_pisa.scala 76:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[executor_pisa.scala 76:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[executor_pisa.scala 76:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[executor_pisa.scala 76:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[executor_pisa.scala 76:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[executor_pisa.scala 76:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[executor_pisa.scala 76:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[executor_pisa.scala 76:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[executor_pisa.scala 76:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[executor_pisa.scala 76:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[executor_pisa.scala 76:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[executor_pisa.scala 76:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[executor_pisa.scala 76:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[executor_pisa.scala 76:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[executor_pisa.scala 76:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[executor_pisa.scala 76:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[executor_pisa.scala 76:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[executor_pisa.scala 76:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[executor_pisa.scala 76:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[executor_pisa.scala 76:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[executor_pisa.scala 76:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[executor_pisa.scala 76:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[executor_pisa.scala 76:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[executor_pisa.scala 76:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[executor_pisa.scala 76:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[executor_pisa.scala 76:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[executor_pisa.scala 76:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[executor_pisa.scala 76:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[executor_pisa.scala 76:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[executor_pisa.scala 76:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[executor_pisa.scala 76:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[executor_pisa.scala 76:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[executor_pisa.scala 76:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[executor_pisa.scala 76:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[executor_pisa.scala 76:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[executor_pisa.scala 76:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[executor_pisa.scala 76:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[executor_pisa.scala 76:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[executor_pisa.scala 76:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[executor_pisa.scala 76:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[executor_pisa.scala 76:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[executor_pisa.scala 76:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[executor_pisa.scala 76:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[executor_pisa.scala 76:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[executor_pisa.scala 76:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[executor_pisa.scala 76:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[executor_pisa.scala 76:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[executor_pisa.scala 76:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[executor_pisa.scala 76:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[executor_pisa.scala 76:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[executor_pisa.scala 76:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[executor_pisa.scala 76:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[executor_pisa.scala 76:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[executor_pisa.scala 76:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[executor_pisa.scala 76:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[executor_pisa.scala 76:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[executor_pisa.scala 76:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[executor_pisa.scala 76:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[executor_pisa.scala 76:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[executor_pisa.scala 76:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[executor_pisa.scala 76:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[executor_pisa.scala 76:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[executor_pisa.scala 76:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[executor_pisa.scala 76:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[executor_pisa.scala 76:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[executor_pisa.scala 76:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[executor_pisa.scala 76:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[executor_pisa.scala 76:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[executor_pisa.scala 76:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[executor_pisa.scala 76:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[executor_pisa.scala 76:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[executor_pisa.scala 76:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[executor_pisa.scala 76:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[executor_pisa.scala 76:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[executor_pisa.scala 76:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[executor_pisa.scala 76:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[executor_pisa.scala 76:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[executor_pisa.scala 76:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[executor_pisa.scala 76:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[executor_pisa.scala 76:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[executor_pisa.scala 76:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[executor_pisa.scala 76:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[executor_pisa.scala 76:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[executor_pisa.scala 76:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[executor_pisa.scala 76:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[executor_pisa.scala 76:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[executor_pisa.scala 76:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[executor_pisa.scala 76:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[executor_pisa.scala 76:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[executor_pisa.scala 76:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[executor_pisa.scala 76:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[executor_pisa.scala 76:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[executor_pisa.scala 76:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[executor_pisa.scala 76:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[executor_pisa.scala 76:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[executor_pisa.scala 76:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[executor_pisa.scala 76:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[executor_pisa.scala 76:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[executor_pisa.scala 76:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[executor_pisa.scala 76:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[executor_pisa.scala 76:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[executor_pisa.scala 76:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[executor_pisa.scala 76:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[executor_pisa.scala 76:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[executor_pisa.scala 76:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[executor_pisa.scala 76:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[executor_pisa.scala 76:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[executor_pisa.scala 76:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[executor_pisa.scala 76:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[executor_pisa.scala 76:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[executor_pisa.scala 76:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[executor_pisa.scala 76:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[executor_pisa.scala 76:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[executor_pisa.scala 76:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[executor_pisa.scala 76:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[executor_pisa.scala 76:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[executor_pisa.scala 76:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[executor_pisa.scala 76:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[executor_pisa.scala 76:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[executor_pisa.scala 76:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[executor_pisa.scala 76:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[executor_pisa.scala 76:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[executor_pisa.scala 76:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[executor_pisa.scala 76:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[executor_pisa.scala 76:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[executor_pisa.scala 76:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[executor_pisa.scala 76:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[executor_pisa.scala 76:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[executor_pisa.scala 76:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[executor_pisa.scala 76:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[executor_pisa.scala 76:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[executor_pisa.scala 76:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[executor_pisa.scala 76:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[executor_pisa.scala 76:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[executor_pisa.scala 76:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[executor_pisa.scala 76:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[executor_pisa.scala 76:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[executor_pisa.scala 76:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[executor_pisa.scala 76:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[executor_pisa.scala 76:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[executor_pisa.scala 76:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[executor_pisa.scala 76:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[executor_pisa.scala 76:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[executor_pisa.scala 76:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[executor_pisa.scala 76:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[executor_pisa.scala 76:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[executor_pisa.scala 76:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[executor_pisa.scala 76:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[executor_pisa.scala 76:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[executor_pisa.scala 76:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[executor_pisa.scala 76:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[executor_pisa.scala 76:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[executor_pisa.scala 76:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[executor_pisa.scala 76:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[executor_pisa.scala 76:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[executor_pisa.scala 76:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[executor_pisa.scala 76:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[executor_pisa.scala 76:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[executor_pisa.scala 76:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[executor_pisa.scala 76:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[executor_pisa.scala 76:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[executor_pisa.scala 76:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[executor_pisa.scala 76:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[executor_pisa.scala 76:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[executor_pisa.scala 76:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[executor_pisa.scala 76:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[executor_pisa.scala 76:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[executor_pisa.scala 76:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[executor_pisa.scala 76:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[executor_pisa.scala 76:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[executor_pisa.scala 76:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[executor_pisa.scala 76:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[executor_pisa.scala 76:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[executor_pisa.scala 76:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[executor_pisa.scala 76:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[executor_pisa.scala 76:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[executor_pisa.scala 76:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[executor_pisa.scala 76:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[executor_pisa.scala 76:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[executor_pisa.scala 76:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[executor_pisa.scala 76:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[executor_pisa.scala 76:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[executor_pisa.scala 76:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[executor_pisa.scala 76:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[executor_pisa.scala 76:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[executor_pisa.scala 76:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[executor_pisa.scala 76:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[executor_pisa.scala 76:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[executor_pisa.scala 76:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[executor_pisa.scala 76:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[executor_pisa.scala 76:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[executor_pisa.scala 76:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[executor_pisa.scala 76:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[executor_pisa.scala 76:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[executor_pisa.scala 76:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[executor_pisa.scala 76:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[executor_pisa.scala 76:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[executor_pisa.scala 76:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[executor_pisa.scala 76:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[executor_pisa.scala 76:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[executor_pisa.scala 76:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[executor_pisa.scala 76:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[executor_pisa.scala 76:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[executor_pisa.scala 76:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[executor_pisa.scala 76:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[executor_pisa.scala 76:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[executor_pisa.scala 76:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[executor_pisa.scala 76:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[executor_pisa.scala 76:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[executor_pisa.scala 76:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[executor_pisa.scala 76:13]
    args_0 <= io_args_in_0; // @[executor_pisa.scala 80:14]
    args_1 <= io_args_in_1; // @[executor_pisa.scala 80:14]
    args_2 <= io_args_in_2; // @[executor_pisa.scala 80:14]
    args_3 <= io_args_in_3; // @[executor_pisa.scala 80:14]
    args_4 <= io_args_in_4; // @[executor_pisa.scala 80:14]
    args_5 <= io_args_in_5; // @[executor_pisa.scala 80:14]
    args_6 <= io_args_in_6; // @[executor_pisa.scala 80:14]
    vliw_0 <= io_vliw_in_0; // @[executor_pisa.scala 84:14]
    vliw_1 <= io_vliw_in_1; // @[executor_pisa.scala 84:14]
    vliw_2 <= io_vliw_in_2; // @[executor_pisa.scala 84:14]
    vliw_3 <= io_vliw_in_3; // @[executor_pisa.scala 84:14]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  phv_next_config_id = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  args_0 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  args_1 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  args_2 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  args_3 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  args_4 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  args_5 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  args_6 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  vliw_0 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  vliw_1 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  vliw_2 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  vliw_3 = _RAND_269[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
