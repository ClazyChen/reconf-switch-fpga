module OutPort(
  input         clock,
  input  [7:0]  io_phv_in_data_0,
  input  [7:0]  io_phv_in_data_1,
  input  [7:0]  io_phv_in_data_2,
  input  [7:0]  io_phv_in_data_3,
  input  [7:0]  io_phv_in_data_4,
  input  [7:0]  io_phv_in_data_5,
  input  [7:0]  io_phv_in_data_6,
  input  [7:0]  io_phv_in_data_7,
  input  [7:0]  io_phv_in_data_8,
  input  [7:0]  io_phv_in_data_9,
  input  [7:0]  io_phv_in_data_10,
  input  [7:0]  io_phv_in_data_11,
  input  [7:0]  io_phv_in_data_12,
  input  [7:0]  io_phv_in_data_13,
  input  [7:0]  io_phv_in_data_14,
  input  [7:0]  io_phv_in_data_15,
  input  [7:0]  io_phv_in_data_16,
  input  [7:0]  io_phv_in_data_17,
  input  [7:0]  io_phv_in_data_18,
  input  [7:0]  io_phv_in_data_19,
  input  [7:0]  io_phv_in_data_20,
  input  [7:0]  io_phv_in_data_21,
  input  [7:0]  io_phv_in_data_22,
  input  [7:0]  io_phv_in_data_23,
  input  [7:0]  io_phv_in_data_24,
  input  [7:0]  io_phv_in_data_25,
  input  [7:0]  io_phv_in_data_26,
  input  [7:0]  io_phv_in_data_27,
  input  [7:0]  io_phv_in_data_28,
  input  [7:0]  io_phv_in_data_29,
  input  [7:0]  io_phv_in_data_30,
  input  [7:0]  io_phv_in_data_31,
  input  [7:0]  io_phv_in_data_32,
  input  [7:0]  io_phv_in_data_33,
  input  [7:0]  io_phv_in_data_34,
  input  [7:0]  io_phv_in_data_35,
  input  [7:0]  io_phv_in_data_36,
  input  [7:0]  io_phv_in_data_37,
  input  [7:0]  io_phv_in_data_38,
  input  [7:0]  io_phv_in_data_39,
  input  [7:0]  io_phv_in_data_40,
  input  [7:0]  io_phv_in_data_41,
  input  [7:0]  io_phv_in_data_42,
  input  [7:0]  io_phv_in_data_43,
  input  [7:0]  io_phv_in_data_44,
  input  [7:0]  io_phv_in_data_45,
  input  [7:0]  io_phv_in_data_46,
  input  [7:0]  io_phv_in_data_47,
  input  [7:0]  io_phv_in_data_48,
  input  [7:0]  io_phv_in_data_49,
  input  [7:0]  io_phv_in_data_50,
  input  [7:0]  io_phv_in_data_51,
  input  [7:0]  io_phv_in_data_52,
  input  [7:0]  io_phv_in_data_53,
  input  [7:0]  io_phv_in_data_54,
  input  [7:0]  io_phv_in_data_55,
  input  [7:0]  io_phv_in_data_56,
  input  [7:0]  io_phv_in_data_57,
  input  [7:0]  io_phv_in_data_58,
  input  [7:0]  io_phv_in_data_59,
  input  [7:0]  io_phv_in_data_60,
  input  [7:0]  io_phv_in_data_61,
  input  [7:0]  io_phv_in_data_62,
  input  [7:0]  io_phv_in_data_63,
  input  [7:0]  io_phv_in_data_64,
  input  [7:0]  io_phv_in_data_65,
  input  [7:0]  io_phv_in_data_66,
  input  [7:0]  io_phv_in_data_67,
  input  [7:0]  io_phv_in_data_68,
  input  [7:0]  io_phv_in_data_69,
  input  [7:0]  io_phv_in_data_70,
  input  [7:0]  io_phv_in_data_71,
  input  [7:0]  io_phv_in_data_72,
  input  [7:0]  io_phv_in_data_73,
  input  [7:0]  io_phv_in_data_74,
  input  [7:0]  io_phv_in_data_75,
  input  [7:0]  io_phv_in_data_76,
  input  [7:0]  io_phv_in_data_77,
  input  [7:0]  io_phv_in_data_78,
  input  [7:0]  io_phv_in_data_79,
  input  [7:0]  io_phv_in_data_80,
  input  [7:0]  io_phv_in_data_81,
  input  [7:0]  io_phv_in_data_82,
  input  [7:0]  io_phv_in_data_83,
  input  [7:0]  io_phv_in_data_84,
  input  [7:0]  io_phv_in_data_85,
  input  [7:0]  io_phv_in_data_86,
  input  [7:0]  io_phv_in_data_87,
  input  [7:0]  io_phv_in_data_88,
  input  [7:0]  io_phv_in_data_89,
  input  [7:0]  io_phv_in_data_90,
  input  [7:0]  io_phv_in_data_91,
  input  [7:0]  io_phv_in_data_92,
  input  [7:0]  io_phv_in_data_93,
  input  [7:0]  io_phv_in_data_94,
  input  [7:0]  io_phv_in_data_95,
  input  [7:0]  io_phv_in_data_96,
  input  [7:0]  io_phv_in_data_97,
  input  [7:0]  io_phv_in_data_98,
  input  [7:0]  io_phv_in_data_99,
  input  [7:0]  io_phv_in_data_100,
  input  [7:0]  io_phv_in_data_101,
  input  [7:0]  io_phv_in_data_102,
  input  [7:0]  io_phv_in_data_103,
  input  [7:0]  io_phv_in_data_104,
  input  [7:0]  io_phv_in_data_105,
  input  [7:0]  io_phv_in_data_106,
  input  [7:0]  io_phv_in_data_107,
  input  [7:0]  io_phv_in_data_108,
  input  [7:0]  io_phv_in_data_109,
  input  [7:0]  io_phv_in_data_110,
  input  [7:0]  io_phv_in_data_111,
  input  [7:0]  io_phv_in_data_112,
  input  [7:0]  io_phv_in_data_113,
  input  [7:0]  io_phv_in_data_114,
  input  [7:0]  io_phv_in_data_115,
  input  [7:0]  io_phv_in_data_116,
  input  [7:0]  io_phv_in_data_117,
  input  [7:0]  io_phv_in_data_118,
  input  [7:0]  io_phv_in_data_119,
  input  [7:0]  io_phv_in_data_120,
  input  [7:0]  io_phv_in_data_121,
  input  [7:0]  io_phv_in_data_122,
  input  [7:0]  io_phv_in_data_123,
  input  [7:0]  io_phv_in_data_124,
  input  [7:0]  io_phv_in_data_125,
  input  [7:0]  io_phv_in_data_126,
  input  [7:0]  io_phv_in_data_127,
  input  [7:0]  io_phv_in_data_128,
  input  [7:0]  io_phv_in_data_129,
  input  [7:0]  io_phv_in_data_130,
  input  [7:0]  io_phv_in_data_131,
  input  [7:0]  io_phv_in_data_132,
  input  [7:0]  io_phv_in_data_133,
  input  [7:0]  io_phv_in_data_134,
  input  [7:0]  io_phv_in_data_135,
  input  [7:0]  io_phv_in_data_136,
  input  [7:0]  io_phv_in_data_137,
  input  [7:0]  io_phv_in_data_138,
  input  [7:0]  io_phv_in_data_139,
  input  [7:0]  io_phv_in_data_140,
  input  [7:0]  io_phv_in_data_141,
  input  [7:0]  io_phv_in_data_142,
  input  [7:0]  io_phv_in_data_143,
  input  [7:0]  io_phv_in_data_144,
  input  [7:0]  io_phv_in_data_145,
  input  [7:0]  io_phv_in_data_146,
  input  [7:0]  io_phv_in_data_147,
  input  [7:0]  io_phv_in_data_148,
  input  [7:0]  io_phv_in_data_149,
  input  [7:0]  io_phv_in_data_150,
  input  [7:0]  io_phv_in_data_151,
  input  [7:0]  io_phv_in_data_152,
  input  [7:0]  io_phv_in_data_153,
  input  [7:0]  io_phv_in_data_154,
  input  [7:0]  io_phv_in_data_155,
  input  [7:0]  io_phv_in_data_156,
  input  [7:0]  io_phv_in_data_157,
  input  [7:0]  io_phv_in_data_158,
  input  [7:0]  io_phv_in_data_159,
  input  [7:0]  io_phv_in_data_160,
  input  [7:0]  io_phv_in_data_161,
  input  [7:0]  io_phv_in_data_162,
  input  [7:0]  io_phv_in_data_163,
  input  [7:0]  io_phv_in_data_164,
  input  [7:0]  io_phv_in_data_165,
  input  [7:0]  io_phv_in_data_166,
  input  [7:0]  io_phv_in_data_167,
  input  [7:0]  io_phv_in_data_168,
  input  [7:0]  io_phv_in_data_169,
  input  [7:0]  io_phv_in_data_170,
  input  [7:0]  io_phv_in_data_171,
  input  [7:0]  io_phv_in_data_172,
  input  [7:0]  io_phv_in_data_173,
  input  [7:0]  io_phv_in_data_174,
  input  [7:0]  io_phv_in_data_175,
  input  [7:0]  io_phv_in_data_176,
  input  [7:0]  io_phv_in_data_177,
  input  [7:0]  io_phv_in_data_178,
  input  [7:0]  io_phv_in_data_179,
  input  [7:0]  io_phv_in_data_180,
  input  [7:0]  io_phv_in_data_181,
  input  [7:0]  io_phv_in_data_182,
  input  [7:0]  io_phv_in_data_183,
  input  [7:0]  io_phv_in_data_184,
  input  [7:0]  io_phv_in_data_185,
  input  [7:0]  io_phv_in_data_186,
  input  [7:0]  io_phv_in_data_187,
  input  [7:0]  io_phv_in_data_188,
  input  [7:0]  io_phv_in_data_189,
  input  [7:0]  io_phv_in_data_190,
  input  [7:0]  io_phv_in_data_191,
  input  [7:0]  io_phv_in_data_192,
  input  [7:0]  io_phv_in_data_193,
  input  [7:0]  io_phv_in_data_194,
  input  [7:0]  io_phv_in_data_195,
  input  [7:0]  io_phv_in_data_196,
  input  [7:0]  io_phv_in_data_197,
  input  [7:0]  io_phv_in_data_198,
  input  [7:0]  io_phv_in_data_199,
  input  [7:0]  io_phv_in_data_200,
  input  [7:0]  io_phv_in_data_201,
  input  [7:0]  io_phv_in_data_202,
  input  [7:0]  io_phv_in_data_203,
  input  [7:0]  io_phv_in_data_204,
  input  [7:0]  io_phv_in_data_205,
  input  [7:0]  io_phv_in_data_206,
  input  [7:0]  io_phv_in_data_207,
  input  [7:0]  io_phv_in_data_208,
  input  [7:0]  io_phv_in_data_209,
  input  [7:0]  io_phv_in_data_210,
  input  [7:0]  io_phv_in_data_211,
  input  [7:0]  io_phv_in_data_212,
  input  [7:0]  io_phv_in_data_213,
  input  [7:0]  io_phv_in_data_214,
  input  [7:0]  io_phv_in_data_215,
  input  [7:0]  io_phv_in_data_216,
  input  [7:0]  io_phv_in_data_217,
  input  [7:0]  io_phv_in_data_218,
  input  [7:0]  io_phv_in_data_219,
  input  [7:0]  io_phv_in_data_220,
  input  [7:0]  io_phv_in_data_221,
  input  [7:0]  io_phv_in_data_222,
  input  [7:0]  io_phv_in_data_223,
  input  [7:0]  io_phv_in_data_224,
  input  [7:0]  io_phv_in_data_225,
  input  [7:0]  io_phv_in_data_226,
  input  [7:0]  io_phv_in_data_227,
  input  [7:0]  io_phv_in_data_228,
  input  [7:0]  io_phv_in_data_229,
  input  [7:0]  io_phv_in_data_230,
  input  [7:0]  io_phv_in_data_231,
  input  [7:0]  io_phv_in_data_232,
  input  [7:0]  io_phv_in_data_233,
  input  [7:0]  io_phv_in_data_234,
  input  [7:0]  io_phv_in_data_235,
  input  [7:0]  io_phv_in_data_236,
  input  [7:0]  io_phv_in_data_237,
  input  [7:0]  io_phv_in_data_238,
  input  [7:0]  io_phv_in_data_239,
  input  [7:0]  io_phv_in_data_240,
  input  [7:0]  io_phv_in_data_241,
  input  [7:0]  io_phv_in_data_242,
  input  [7:0]  io_phv_in_data_243,
  input  [7:0]  io_phv_in_data_244,
  input  [7:0]  io_phv_in_data_245,
  input  [7:0]  io_phv_in_data_246,
  input  [7:0]  io_phv_in_data_247,
  input  [7:0]  io_phv_in_data_248,
  input  [7:0]  io_phv_in_data_249,
  input  [7:0]  io_phv_in_data_250,
  input  [7:0]  io_phv_in_data_251,
  input  [7:0]  io_phv_in_data_252,
  input  [7:0]  io_phv_in_data_253,
  input  [7:0]  io_phv_in_data_254,
  input  [7:0]  io_phv_in_data_255,
  input  [7:0]  io_phv_in_data_256,
  input  [7:0]  io_phv_in_data_257,
  input  [7:0]  io_phv_in_data_258,
  input  [7:0]  io_phv_in_data_259,
  input  [7:0]  io_phv_in_data_260,
  input  [7:0]  io_phv_in_data_261,
  input  [7:0]  io_phv_in_data_262,
  input  [7:0]  io_phv_in_data_263,
  input  [7:0]  io_phv_in_data_264,
  input  [7:0]  io_phv_in_data_265,
  input  [7:0]  io_phv_in_data_266,
  input  [7:0]  io_phv_in_data_267,
  input  [7:0]  io_phv_in_data_268,
  input  [7:0]  io_phv_in_data_269,
  input  [7:0]  io_phv_in_data_270,
  input  [7:0]  io_phv_in_data_271,
  input  [7:0]  io_phv_in_data_272,
  input  [7:0]  io_phv_in_data_273,
  input  [7:0]  io_phv_in_data_274,
  input  [7:0]  io_phv_in_data_275,
  input  [7:0]  io_phv_in_data_276,
  input  [7:0]  io_phv_in_data_277,
  input  [7:0]  io_phv_in_data_278,
  input  [7:0]  io_phv_in_data_279,
  input  [7:0]  io_phv_in_data_280,
  input  [7:0]  io_phv_in_data_281,
  input  [7:0]  io_phv_in_data_282,
  input  [7:0]  io_phv_in_data_283,
  input  [7:0]  io_phv_in_data_284,
  input  [7:0]  io_phv_in_data_285,
  input  [7:0]  io_phv_in_data_286,
  input  [7:0]  io_phv_in_data_287,
  input  [7:0]  io_phv_in_data_288,
  input  [7:0]  io_phv_in_data_289,
  input  [7:0]  io_phv_in_data_290,
  input  [7:0]  io_phv_in_data_291,
  input  [7:0]  io_phv_in_data_292,
  input  [7:0]  io_phv_in_data_293,
  input  [7:0]  io_phv_in_data_294,
  input  [7:0]  io_phv_in_data_295,
  input  [7:0]  io_phv_in_data_296,
  input  [7:0]  io_phv_in_data_297,
  input  [7:0]  io_phv_in_data_298,
  input  [7:0]  io_phv_in_data_299,
  input  [7:0]  io_phv_in_data_300,
  input  [7:0]  io_phv_in_data_301,
  input  [7:0]  io_phv_in_data_302,
  input  [7:0]  io_phv_in_data_303,
  input  [7:0]  io_phv_in_data_304,
  input  [7:0]  io_phv_in_data_305,
  input  [7:0]  io_phv_in_data_306,
  input  [7:0]  io_phv_in_data_307,
  input  [7:0]  io_phv_in_data_308,
  input  [7:0]  io_phv_in_data_309,
  input  [7:0]  io_phv_in_data_310,
  input  [7:0]  io_phv_in_data_311,
  input  [7:0]  io_phv_in_data_312,
  input  [7:0]  io_phv_in_data_313,
  input  [7:0]  io_phv_in_data_314,
  input  [7:0]  io_phv_in_data_315,
  input  [7:0]  io_phv_in_data_316,
  input  [7:0]  io_phv_in_data_317,
  input  [7:0]  io_phv_in_data_318,
  input  [7:0]  io_phv_in_data_319,
  input  [7:0]  io_phv_in_data_320,
  input  [7:0]  io_phv_in_data_321,
  input  [7:0]  io_phv_in_data_322,
  input  [7:0]  io_phv_in_data_323,
  input  [7:0]  io_phv_in_data_324,
  input  [7:0]  io_phv_in_data_325,
  input  [7:0]  io_phv_in_data_326,
  input  [7:0]  io_phv_in_data_327,
  input  [7:0]  io_phv_in_data_328,
  input  [7:0]  io_phv_in_data_329,
  input  [7:0]  io_phv_in_data_330,
  input  [7:0]  io_phv_in_data_331,
  input  [7:0]  io_phv_in_data_332,
  input  [7:0]  io_phv_in_data_333,
  input  [7:0]  io_phv_in_data_334,
  input  [7:0]  io_phv_in_data_335,
  input  [7:0]  io_phv_in_data_336,
  input  [7:0]  io_phv_in_data_337,
  input  [7:0]  io_phv_in_data_338,
  input  [7:0]  io_phv_in_data_339,
  input  [7:0]  io_phv_in_data_340,
  input  [7:0]  io_phv_in_data_341,
  input  [7:0]  io_phv_in_data_342,
  input  [7:0]  io_phv_in_data_343,
  input  [7:0]  io_phv_in_data_344,
  input  [7:0]  io_phv_in_data_345,
  input  [7:0]  io_phv_in_data_346,
  input  [7:0]  io_phv_in_data_347,
  input  [7:0]  io_phv_in_data_348,
  input  [7:0]  io_phv_in_data_349,
  input  [7:0]  io_phv_in_data_350,
  input  [7:0]  io_phv_in_data_351,
  input  [7:0]  io_phv_in_data_352,
  input  [7:0]  io_phv_in_data_353,
  input  [7:0]  io_phv_in_data_354,
  input  [7:0]  io_phv_in_data_355,
  input  [7:0]  io_phv_in_data_356,
  input  [7:0]  io_phv_in_data_357,
  input  [7:0]  io_phv_in_data_358,
  input  [7:0]  io_phv_in_data_359,
  input  [7:0]  io_phv_in_data_360,
  input  [7:0]  io_phv_in_data_361,
  input  [7:0]  io_phv_in_data_362,
  input  [7:0]  io_phv_in_data_363,
  input  [7:0]  io_phv_in_data_364,
  input  [7:0]  io_phv_in_data_365,
  input  [7:0]  io_phv_in_data_366,
  input  [7:0]  io_phv_in_data_367,
  input  [7:0]  io_phv_in_data_368,
  input  [7:0]  io_phv_in_data_369,
  input  [7:0]  io_phv_in_data_370,
  input  [7:0]  io_phv_in_data_371,
  input  [7:0]  io_phv_in_data_372,
  input  [7:0]  io_phv_in_data_373,
  input  [7:0]  io_phv_in_data_374,
  input  [7:0]  io_phv_in_data_375,
  input  [7:0]  io_phv_in_data_376,
  input  [7:0]  io_phv_in_data_377,
  input  [7:0]  io_phv_in_data_378,
  input  [7:0]  io_phv_in_data_379,
  input  [7:0]  io_phv_in_data_380,
  input  [7:0]  io_phv_in_data_381,
  input  [7:0]  io_phv_in_data_382,
  input  [7:0]  io_phv_in_data_383,
  input  [7:0]  io_phv_in_data_384,
  input  [7:0]  io_phv_in_data_385,
  input  [7:0]  io_phv_in_data_386,
  input  [7:0]  io_phv_in_data_387,
  input  [7:0]  io_phv_in_data_388,
  input  [7:0]  io_phv_in_data_389,
  input  [7:0]  io_phv_in_data_390,
  input  [7:0]  io_phv_in_data_391,
  input  [7:0]  io_phv_in_data_392,
  input  [7:0]  io_phv_in_data_393,
  input  [7:0]  io_phv_in_data_394,
  input  [7:0]  io_phv_in_data_395,
  input  [7:0]  io_phv_in_data_396,
  input  [7:0]  io_phv_in_data_397,
  input  [7:0]  io_phv_in_data_398,
  input  [7:0]  io_phv_in_data_399,
  input  [7:0]  io_phv_in_data_400,
  input  [7:0]  io_phv_in_data_401,
  input  [7:0]  io_phv_in_data_402,
  input  [7:0]  io_phv_in_data_403,
  input  [7:0]  io_phv_in_data_404,
  input  [7:0]  io_phv_in_data_405,
  input  [7:0]  io_phv_in_data_406,
  input  [7:0]  io_phv_in_data_407,
  input  [7:0]  io_phv_in_data_408,
  input  [7:0]  io_phv_in_data_409,
  input  [7:0]  io_phv_in_data_410,
  input  [7:0]  io_phv_in_data_411,
  input  [7:0]  io_phv_in_data_412,
  input  [7:0]  io_phv_in_data_413,
  input  [7:0]  io_phv_in_data_414,
  input  [7:0]  io_phv_in_data_415,
  input  [7:0]  io_phv_in_data_416,
  input  [7:0]  io_phv_in_data_417,
  input  [7:0]  io_phv_in_data_418,
  input  [7:0]  io_phv_in_data_419,
  input  [7:0]  io_phv_in_data_420,
  input  [7:0]  io_phv_in_data_421,
  input  [7:0]  io_phv_in_data_422,
  input  [7:0]  io_phv_in_data_423,
  input  [7:0]  io_phv_in_data_424,
  input  [7:0]  io_phv_in_data_425,
  input  [7:0]  io_phv_in_data_426,
  input  [7:0]  io_phv_in_data_427,
  input  [7:0]  io_phv_in_data_428,
  input  [7:0]  io_phv_in_data_429,
  input  [7:0]  io_phv_in_data_430,
  input  [7:0]  io_phv_in_data_431,
  input  [7:0]  io_phv_in_data_432,
  input  [7:0]  io_phv_in_data_433,
  input  [7:0]  io_phv_in_data_434,
  input  [7:0]  io_phv_in_data_435,
  input  [7:0]  io_phv_in_data_436,
  input  [7:0]  io_phv_in_data_437,
  input  [7:0]  io_phv_in_data_438,
  input  [7:0]  io_phv_in_data_439,
  input  [7:0]  io_phv_in_data_440,
  input  [7:0]  io_phv_in_data_441,
  input  [7:0]  io_phv_in_data_442,
  input  [7:0]  io_phv_in_data_443,
  input  [7:0]  io_phv_in_data_444,
  input  [7:0]  io_phv_in_data_445,
  input  [7:0]  io_phv_in_data_446,
  input  [7:0]  io_phv_in_data_447,
  input  [7:0]  io_phv_in_data_448,
  input  [7:0]  io_phv_in_data_449,
  input  [7:0]  io_phv_in_data_450,
  input  [7:0]  io_phv_in_data_451,
  input  [7:0]  io_phv_in_data_452,
  input  [7:0]  io_phv_in_data_453,
  input  [7:0]  io_phv_in_data_454,
  input  [7:0]  io_phv_in_data_455,
  input  [7:0]  io_phv_in_data_456,
  input  [7:0]  io_phv_in_data_457,
  input  [7:0]  io_phv_in_data_458,
  input  [7:0]  io_phv_in_data_459,
  input  [7:0]  io_phv_in_data_460,
  input  [7:0]  io_phv_in_data_461,
  input  [7:0]  io_phv_in_data_462,
  input  [7:0]  io_phv_in_data_463,
  input  [7:0]  io_phv_in_data_464,
  input  [7:0]  io_phv_in_data_465,
  input  [7:0]  io_phv_in_data_466,
  input  [7:0]  io_phv_in_data_467,
  input  [7:0]  io_phv_in_data_468,
  input  [7:0]  io_phv_in_data_469,
  input  [7:0]  io_phv_in_data_470,
  input  [7:0]  io_phv_in_data_471,
  input  [7:0]  io_phv_in_data_472,
  input  [7:0]  io_phv_in_data_473,
  input  [7:0]  io_phv_in_data_474,
  input  [7:0]  io_phv_in_data_475,
  input  [7:0]  io_phv_in_data_476,
  input  [7:0]  io_phv_in_data_477,
  input  [7:0]  io_phv_in_data_478,
  input  [7:0]  io_phv_in_data_479,
  input  [7:0]  io_phv_in_data_480,
  input  [7:0]  io_phv_in_data_481,
  input  [7:0]  io_phv_in_data_482,
  input  [7:0]  io_phv_in_data_483,
  input  [7:0]  io_phv_in_data_484,
  input  [7:0]  io_phv_in_data_485,
  input  [7:0]  io_phv_in_data_486,
  input  [7:0]  io_phv_in_data_487,
  input  [7:0]  io_phv_in_data_488,
  input  [7:0]  io_phv_in_data_489,
  input  [7:0]  io_phv_in_data_490,
  input  [7:0]  io_phv_in_data_491,
  input  [7:0]  io_phv_in_data_492,
  input  [7:0]  io_phv_in_data_493,
  input  [7:0]  io_phv_in_data_494,
  input  [7:0]  io_phv_in_data_495,
  input  [7:0]  io_phv_in_data_496,
  input  [7:0]  io_phv_in_data_497,
  input  [7:0]  io_phv_in_data_498,
  input  [7:0]  io_phv_in_data_499,
  input  [7:0]  io_phv_in_data_500,
  input  [7:0]  io_phv_in_data_501,
  input  [7:0]  io_phv_in_data_502,
  input  [7:0]  io_phv_in_data_503,
  input  [7:0]  io_phv_in_data_504,
  input  [7:0]  io_phv_in_data_505,
  input  [7:0]  io_phv_in_data_506,
  input  [7:0]  io_phv_in_data_507,
  input  [7:0]  io_phv_in_data_508,
  input  [7:0]  io_phv_in_data_509,
  input  [7:0]  io_phv_in_data_510,
  input  [7:0]  io_phv_in_data_511,
  input  [5:0]  io_pcie_o_cs,
  input         io_pcie_o_r_en,
  input  [7:0]  io_pcie_o_r_addr,
  output [63:0] io_pcie_o_r_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  sram_0_clock; // @[outport.scala 23:25]
  wire  sram_0_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_0_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_0_io_w_data; // @[outport.scala 23:25]
  wire  sram_0_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_0_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_0_io_r_data; // @[outport.scala 23:25]
  wire  sram_1_clock; // @[outport.scala 23:25]
  wire  sram_1_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_1_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_1_io_w_data; // @[outport.scala 23:25]
  wire  sram_1_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_1_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_1_io_r_data; // @[outport.scala 23:25]
  wire  sram_2_clock; // @[outport.scala 23:25]
  wire  sram_2_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_2_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_2_io_w_data; // @[outport.scala 23:25]
  wire  sram_2_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_2_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_2_io_r_data; // @[outport.scala 23:25]
  wire  sram_3_clock; // @[outport.scala 23:25]
  wire  sram_3_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_3_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_3_io_w_data; // @[outport.scala 23:25]
  wire  sram_3_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_3_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_3_io_r_data; // @[outport.scala 23:25]
  wire  sram_4_clock; // @[outport.scala 23:25]
  wire  sram_4_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_4_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_4_io_w_data; // @[outport.scala 23:25]
  wire  sram_4_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_4_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_4_io_r_data; // @[outport.scala 23:25]
  wire  sram_5_clock; // @[outport.scala 23:25]
  wire  sram_5_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_5_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_5_io_w_data; // @[outport.scala 23:25]
  wire  sram_5_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_5_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_5_io_r_data; // @[outport.scala 23:25]
  wire  sram_6_clock; // @[outport.scala 23:25]
  wire  sram_6_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_6_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_6_io_w_data; // @[outport.scala 23:25]
  wire  sram_6_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_6_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_6_io_r_data; // @[outport.scala 23:25]
  wire  sram_7_clock; // @[outport.scala 23:25]
  wire  sram_7_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_7_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_7_io_w_data; // @[outport.scala 23:25]
  wire  sram_7_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_7_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_7_io_r_data; // @[outport.scala 23:25]
  wire  sram_8_clock; // @[outport.scala 23:25]
  wire  sram_8_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_8_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_8_io_w_data; // @[outport.scala 23:25]
  wire  sram_8_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_8_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_8_io_r_data; // @[outport.scala 23:25]
  wire  sram_9_clock; // @[outport.scala 23:25]
  wire  sram_9_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_9_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_9_io_w_data; // @[outport.scala 23:25]
  wire  sram_9_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_9_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_9_io_r_data; // @[outport.scala 23:25]
  wire  sram_10_clock; // @[outport.scala 23:25]
  wire  sram_10_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_10_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_10_io_w_data; // @[outport.scala 23:25]
  wire  sram_10_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_10_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_10_io_r_data; // @[outport.scala 23:25]
  wire  sram_11_clock; // @[outport.scala 23:25]
  wire  sram_11_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_11_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_11_io_w_data; // @[outport.scala 23:25]
  wire  sram_11_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_11_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_11_io_r_data; // @[outport.scala 23:25]
  wire  sram_12_clock; // @[outport.scala 23:25]
  wire  sram_12_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_12_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_12_io_w_data; // @[outport.scala 23:25]
  wire  sram_12_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_12_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_12_io_r_data; // @[outport.scala 23:25]
  wire  sram_13_clock; // @[outport.scala 23:25]
  wire  sram_13_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_13_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_13_io_w_data; // @[outport.scala 23:25]
  wire  sram_13_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_13_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_13_io_r_data; // @[outport.scala 23:25]
  wire  sram_14_clock; // @[outport.scala 23:25]
  wire  sram_14_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_14_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_14_io_w_data; // @[outport.scala 23:25]
  wire  sram_14_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_14_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_14_io_r_data; // @[outport.scala 23:25]
  wire  sram_15_clock; // @[outport.scala 23:25]
  wire  sram_15_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_15_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_15_io_w_data; // @[outport.scala 23:25]
  wire  sram_15_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_15_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_15_io_r_data; // @[outport.scala 23:25]
  wire  sram_16_clock; // @[outport.scala 23:25]
  wire  sram_16_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_16_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_16_io_w_data; // @[outport.scala 23:25]
  wire  sram_16_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_16_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_16_io_r_data; // @[outport.scala 23:25]
  wire  sram_17_clock; // @[outport.scala 23:25]
  wire  sram_17_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_17_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_17_io_w_data; // @[outport.scala 23:25]
  wire  sram_17_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_17_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_17_io_r_data; // @[outport.scala 23:25]
  wire  sram_18_clock; // @[outport.scala 23:25]
  wire  sram_18_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_18_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_18_io_w_data; // @[outport.scala 23:25]
  wire  sram_18_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_18_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_18_io_r_data; // @[outport.scala 23:25]
  wire  sram_19_clock; // @[outport.scala 23:25]
  wire  sram_19_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_19_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_19_io_w_data; // @[outport.scala 23:25]
  wire  sram_19_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_19_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_19_io_r_data; // @[outport.scala 23:25]
  wire  sram_20_clock; // @[outport.scala 23:25]
  wire  sram_20_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_20_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_20_io_w_data; // @[outport.scala 23:25]
  wire  sram_20_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_20_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_20_io_r_data; // @[outport.scala 23:25]
  wire  sram_21_clock; // @[outport.scala 23:25]
  wire  sram_21_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_21_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_21_io_w_data; // @[outport.scala 23:25]
  wire  sram_21_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_21_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_21_io_r_data; // @[outport.scala 23:25]
  wire  sram_22_clock; // @[outport.scala 23:25]
  wire  sram_22_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_22_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_22_io_w_data; // @[outport.scala 23:25]
  wire  sram_22_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_22_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_22_io_r_data; // @[outport.scala 23:25]
  wire  sram_23_clock; // @[outport.scala 23:25]
  wire  sram_23_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_23_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_23_io_w_data; // @[outport.scala 23:25]
  wire  sram_23_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_23_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_23_io_r_data; // @[outport.scala 23:25]
  wire  sram_24_clock; // @[outport.scala 23:25]
  wire  sram_24_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_24_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_24_io_w_data; // @[outport.scala 23:25]
  wire  sram_24_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_24_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_24_io_r_data; // @[outport.scala 23:25]
  wire  sram_25_clock; // @[outport.scala 23:25]
  wire  sram_25_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_25_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_25_io_w_data; // @[outport.scala 23:25]
  wire  sram_25_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_25_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_25_io_r_data; // @[outport.scala 23:25]
  wire  sram_26_clock; // @[outport.scala 23:25]
  wire  sram_26_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_26_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_26_io_w_data; // @[outport.scala 23:25]
  wire  sram_26_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_26_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_26_io_r_data; // @[outport.scala 23:25]
  wire  sram_27_clock; // @[outport.scala 23:25]
  wire  sram_27_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_27_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_27_io_w_data; // @[outport.scala 23:25]
  wire  sram_27_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_27_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_27_io_r_data; // @[outport.scala 23:25]
  wire  sram_28_clock; // @[outport.scala 23:25]
  wire  sram_28_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_28_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_28_io_w_data; // @[outport.scala 23:25]
  wire  sram_28_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_28_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_28_io_r_data; // @[outport.scala 23:25]
  wire  sram_29_clock; // @[outport.scala 23:25]
  wire  sram_29_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_29_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_29_io_w_data; // @[outport.scala 23:25]
  wire  sram_29_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_29_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_29_io_r_data; // @[outport.scala 23:25]
  wire  sram_30_clock; // @[outport.scala 23:25]
  wire  sram_30_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_30_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_30_io_w_data; // @[outport.scala 23:25]
  wire  sram_30_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_30_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_30_io_r_data; // @[outport.scala 23:25]
  wire  sram_31_clock; // @[outport.scala 23:25]
  wire  sram_31_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_31_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_31_io_w_data; // @[outport.scala 23:25]
  wire  sram_31_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_31_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_31_io_r_data; // @[outport.scala 23:25]
  wire  sram_32_clock; // @[outport.scala 23:25]
  wire  sram_32_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_32_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_32_io_w_data; // @[outport.scala 23:25]
  wire  sram_32_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_32_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_32_io_r_data; // @[outport.scala 23:25]
  wire  sram_33_clock; // @[outport.scala 23:25]
  wire  sram_33_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_33_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_33_io_w_data; // @[outport.scala 23:25]
  wire  sram_33_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_33_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_33_io_r_data; // @[outport.scala 23:25]
  wire  sram_34_clock; // @[outport.scala 23:25]
  wire  sram_34_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_34_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_34_io_w_data; // @[outport.scala 23:25]
  wire  sram_34_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_34_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_34_io_r_data; // @[outport.scala 23:25]
  wire  sram_35_clock; // @[outport.scala 23:25]
  wire  sram_35_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_35_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_35_io_w_data; // @[outport.scala 23:25]
  wire  sram_35_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_35_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_35_io_r_data; // @[outport.scala 23:25]
  wire  sram_36_clock; // @[outport.scala 23:25]
  wire  sram_36_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_36_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_36_io_w_data; // @[outport.scala 23:25]
  wire  sram_36_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_36_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_36_io_r_data; // @[outport.scala 23:25]
  wire  sram_37_clock; // @[outport.scala 23:25]
  wire  sram_37_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_37_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_37_io_w_data; // @[outport.scala 23:25]
  wire  sram_37_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_37_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_37_io_r_data; // @[outport.scala 23:25]
  wire  sram_38_clock; // @[outport.scala 23:25]
  wire  sram_38_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_38_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_38_io_w_data; // @[outport.scala 23:25]
  wire  sram_38_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_38_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_38_io_r_data; // @[outport.scala 23:25]
  wire  sram_39_clock; // @[outport.scala 23:25]
  wire  sram_39_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_39_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_39_io_w_data; // @[outport.scala 23:25]
  wire  sram_39_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_39_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_39_io_r_data; // @[outport.scala 23:25]
  wire  sram_40_clock; // @[outport.scala 23:25]
  wire  sram_40_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_40_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_40_io_w_data; // @[outport.scala 23:25]
  wire  sram_40_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_40_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_40_io_r_data; // @[outport.scala 23:25]
  wire  sram_41_clock; // @[outport.scala 23:25]
  wire  sram_41_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_41_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_41_io_w_data; // @[outport.scala 23:25]
  wire  sram_41_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_41_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_41_io_r_data; // @[outport.scala 23:25]
  wire  sram_42_clock; // @[outport.scala 23:25]
  wire  sram_42_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_42_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_42_io_w_data; // @[outport.scala 23:25]
  wire  sram_42_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_42_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_42_io_r_data; // @[outport.scala 23:25]
  wire  sram_43_clock; // @[outport.scala 23:25]
  wire  sram_43_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_43_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_43_io_w_data; // @[outport.scala 23:25]
  wire  sram_43_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_43_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_43_io_r_data; // @[outport.scala 23:25]
  wire  sram_44_clock; // @[outport.scala 23:25]
  wire  sram_44_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_44_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_44_io_w_data; // @[outport.scala 23:25]
  wire  sram_44_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_44_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_44_io_r_data; // @[outport.scala 23:25]
  wire  sram_45_clock; // @[outport.scala 23:25]
  wire  sram_45_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_45_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_45_io_w_data; // @[outport.scala 23:25]
  wire  sram_45_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_45_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_45_io_r_data; // @[outport.scala 23:25]
  wire  sram_46_clock; // @[outport.scala 23:25]
  wire  sram_46_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_46_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_46_io_w_data; // @[outport.scala 23:25]
  wire  sram_46_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_46_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_46_io_r_data; // @[outport.scala 23:25]
  wire  sram_47_clock; // @[outport.scala 23:25]
  wire  sram_47_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_47_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_47_io_w_data; // @[outport.scala 23:25]
  wire  sram_47_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_47_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_47_io_r_data; // @[outport.scala 23:25]
  wire  sram_48_clock; // @[outport.scala 23:25]
  wire  sram_48_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_48_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_48_io_w_data; // @[outport.scala 23:25]
  wire  sram_48_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_48_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_48_io_r_data; // @[outport.scala 23:25]
  wire  sram_49_clock; // @[outport.scala 23:25]
  wire  sram_49_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_49_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_49_io_w_data; // @[outport.scala 23:25]
  wire  sram_49_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_49_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_49_io_r_data; // @[outport.scala 23:25]
  wire  sram_50_clock; // @[outport.scala 23:25]
  wire  sram_50_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_50_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_50_io_w_data; // @[outport.scala 23:25]
  wire  sram_50_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_50_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_50_io_r_data; // @[outport.scala 23:25]
  wire  sram_51_clock; // @[outport.scala 23:25]
  wire  sram_51_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_51_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_51_io_w_data; // @[outport.scala 23:25]
  wire  sram_51_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_51_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_51_io_r_data; // @[outport.scala 23:25]
  wire  sram_52_clock; // @[outport.scala 23:25]
  wire  sram_52_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_52_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_52_io_w_data; // @[outport.scala 23:25]
  wire  sram_52_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_52_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_52_io_r_data; // @[outport.scala 23:25]
  wire  sram_53_clock; // @[outport.scala 23:25]
  wire  sram_53_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_53_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_53_io_w_data; // @[outport.scala 23:25]
  wire  sram_53_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_53_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_53_io_r_data; // @[outport.scala 23:25]
  wire  sram_54_clock; // @[outport.scala 23:25]
  wire  sram_54_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_54_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_54_io_w_data; // @[outport.scala 23:25]
  wire  sram_54_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_54_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_54_io_r_data; // @[outport.scala 23:25]
  wire  sram_55_clock; // @[outport.scala 23:25]
  wire  sram_55_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_55_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_55_io_w_data; // @[outport.scala 23:25]
  wire  sram_55_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_55_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_55_io_r_data; // @[outport.scala 23:25]
  wire  sram_56_clock; // @[outport.scala 23:25]
  wire  sram_56_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_56_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_56_io_w_data; // @[outport.scala 23:25]
  wire  sram_56_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_56_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_56_io_r_data; // @[outport.scala 23:25]
  wire  sram_57_clock; // @[outport.scala 23:25]
  wire  sram_57_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_57_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_57_io_w_data; // @[outport.scala 23:25]
  wire  sram_57_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_57_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_57_io_r_data; // @[outport.scala 23:25]
  wire  sram_58_clock; // @[outport.scala 23:25]
  wire  sram_58_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_58_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_58_io_w_data; // @[outport.scala 23:25]
  wire  sram_58_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_58_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_58_io_r_data; // @[outport.scala 23:25]
  wire  sram_59_clock; // @[outport.scala 23:25]
  wire  sram_59_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_59_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_59_io_w_data; // @[outport.scala 23:25]
  wire  sram_59_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_59_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_59_io_r_data; // @[outport.scala 23:25]
  wire  sram_60_clock; // @[outport.scala 23:25]
  wire  sram_60_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_60_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_60_io_w_data; // @[outport.scala 23:25]
  wire  sram_60_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_60_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_60_io_r_data; // @[outport.scala 23:25]
  wire  sram_61_clock; // @[outport.scala 23:25]
  wire  sram_61_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_61_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_61_io_w_data; // @[outport.scala 23:25]
  wire  sram_61_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_61_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_61_io_r_data; // @[outport.scala 23:25]
  wire  sram_62_clock; // @[outport.scala 23:25]
  wire  sram_62_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_62_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_62_io_w_data; // @[outport.scala 23:25]
  wire  sram_62_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_62_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_62_io_r_data; // @[outport.scala 23:25]
  wire  sram_63_clock; // @[outport.scala 23:25]
  wire  sram_63_io_w_en; // @[outport.scala 23:25]
  wire [7:0] sram_63_io_w_addr; // @[outport.scala 23:25]
  wire [63:0] sram_63_io_w_data; // @[outport.scala 23:25]
  wire  sram_63_io_r_en; // @[outport.scala 23:25]
  wire [7:0] sram_63_io_r_addr; // @[outport.scala 23:25]
  wire [63:0] sram_63_io_r_data; // @[outport.scala 23:25]
  reg [7:0] addr; // @[outport.scala 17:19]
  wire [55:0] exe_io_w_data_hi_5 = {io_phv_in_data_0,io_phv_in_data_1,io_phv_in_data_2,io_phv_in_data_3,io_phv_in_data_4
    ,io_phv_in_data_5,io_phv_in_data_6}; // @[Cat.scala 30:58]
  wire  cs_hit = io_pcie_o_cs == 6'h0; // @[outport.scala 31:35]
  wire [63:0] _GEN_0 = cs_hit ? sram_0_io_r_data : 64'h0; // @[outport.scala 34:23 outport.scala 35:31 outport.scala 20:22]
  wire [55:0] exe_io_w_data_hi_11 = {io_phv_in_data_8,io_phv_in_data_9,io_phv_in_data_10,io_phv_in_data_11,
    io_phv_in_data_12,io_phv_in_data_13,io_phv_in_data_14}; // @[Cat.scala 30:58]
  wire  cs_hit_1 = io_pcie_o_cs == 6'h1; // @[outport.scala 31:35]
  wire [63:0] _GEN_1 = cs_hit_1 ? sram_1_io_r_data : _GEN_0; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_17 = {io_phv_in_data_16,io_phv_in_data_17,io_phv_in_data_18,io_phv_in_data_19,
    io_phv_in_data_20,io_phv_in_data_21,io_phv_in_data_22}; // @[Cat.scala 30:58]
  wire  cs_hit_2 = io_pcie_o_cs == 6'h2; // @[outport.scala 31:35]
  wire [63:0] _GEN_2 = cs_hit_2 ? sram_2_io_r_data : _GEN_1; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_23 = {io_phv_in_data_24,io_phv_in_data_25,io_phv_in_data_26,io_phv_in_data_27,
    io_phv_in_data_28,io_phv_in_data_29,io_phv_in_data_30}; // @[Cat.scala 30:58]
  wire  cs_hit_3 = io_pcie_o_cs == 6'h3; // @[outport.scala 31:35]
  wire [63:0] _GEN_3 = cs_hit_3 ? sram_3_io_r_data : _GEN_2; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_29 = {io_phv_in_data_32,io_phv_in_data_33,io_phv_in_data_34,io_phv_in_data_35,
    io_phv_in_data_36,io_phv_in_data_37,io_phv_in_data_38}; // @[Cat.scala 30:58]
  wire  cs_hit_4 = io_pcie_o_cs == 6'h4; // @[outport.scala 31:35]
  wire [63:0] _GEN_4 = cs_hit_4 ? sram_4_io_r_data : _GEN_3; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_35 = {io_phv_in_data_40,io_phv_in_data_41,io_phv_in_data_42,io_phv_in_data_43,
    io_phv_in_data_44,io_phv_in_data_45,io_phv_in_data_46}; // @[Cat.scala 30:58]
  wire  cs_hit_5 = io_pcie_o_cs == 6'h5; // @[outport.scala 31:35]
  wire [63:0] _GEN_5 = cs_hit_5 ? sram_5_io_r_data : _GEN_4; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_41 = {io_phv_in_data_48,io_phv_in_data_49,io_phv_in_data_50,io_phv_in_data_51,
    io_phv_in_data_52,io_phv_in_data_53,io_phv_in_data_54}; // @[Cat.scala 30:58]
  wire  cs_hit_6 = io_pcie_o_cs == 6'h6; // @[outport.scala 31:35]
  wire [63:0] _GEN_6 = cs_hit_6 ? sram_6_io_r_data : _GEN_5; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_47 = {io_phv_in_data_56,io_phv_in_data_57,io_phv_in_data_58,io_phv_in_data_59,
    io_phv_in_data_60,io_phv_in_data_61,io_phv_in_data_62}; // @[Cat.scala 30:58]
  wire  cs_hit_7 = io_pcie_o_cs == 6'h7; // @[outport.scala 31:35]
  wire [63:0] _GEN_7 = cs_hit_7 ? sram_7_io_r_data : _GEN_6; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_53 = {io_phv_in_data_64,io_phv_in_data_65,io_phv_in_data_66,io_phv_in_data_67,
    io_phv_in_data_68,io_phv_in_data_69,io_phv_in_data_70}; // @[Cat.scala 30:58]
  wire  cs_hit_8 = io_pcie_o_cs == 6'h8; // @[outport.scala 31:35]
  wire [63:0] _GEN_8 = cs_hit_8 ? sram_8_io_r_data : _GEN_7; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_59 = {io_phv_in_data_72,io_phv_in_data_73,io_phv_in_data_74,io_phv_in_data_75,
    io_phv_in_data_76,io_phv_in_data_77,io_phv_in_data_78}; // @[Cat.scala 30:58]
  wire  cs_hit_9 = io_pcie_o_cs == 6'h9; // @[outport.scala 31:35]
  wire [63:0] _GEN_9 = cs_hit_9 ? sram_9_io_r_data : _GEN_8; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_65 = {io_phv_in_data_80,io_phv_in_data_81,io_phv_in_data_82,io_phv_in_data_83,
    io_phv_in_data_84,io_phv_in_data_85,io_phv_in_data_86}; // @[Cat.scala 30:58]
  wire  cs_hit_10 = io_pcie_o_cs == 6'ha; // @[outport.scala 31:35]
  wire [63:0] _GEN_10 = cs_hit_10 ? sram_10_io_r_data : _GEN_9; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_71 = {io_phv_in_data_88,io_phv_in_data_89,io_phv_in_data_90,io_phv_in_data_91,
    io_phv_in_data_92,io_phv_in_data_93,io_phv_in_data_94}; // @[Cat.scala 30:58]
  wire  cs_hit_11 = io_pcie_o_cs == 6'hb; // @[outport.scala 31:35]
  wire [63:0] _GEN_11 = cs_hit_11 ? sram_11_io_r_data : _GEN_10; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_77 = {io_phv_in_data_96,io_phv_in_data_97,io_phv_in_data_98,io_phv_in_data_99,
    io_phv_in_data_100,io_phv_in_data_101,io_phv_in_data_102}; // @[Cat.scala 30:58]
  wire  cs_hit_12 = io_pcie_o_cs == 6'hc; // @[outport.scala 31:35]
  wire [63:0] _GEN_12 = cs_hit_12 ? sram_12_io_r_data : _GEN_11; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_83 = {io_phv_in_data_104,io_phv_in_data_105,io_phv_in_data_106,io_phv_in_data_107,
    io_phv_in_data_108,io_phv_in_data_109,io_phv_in_data_110}; // @[Cat.scala 30:58]
  wire  cs_hit_13 = io_pcie_o_cs == 6'hd; // @[outport.scala 31:35]
  wire [63:0] _GEN_13 = cs_hit_13 ? sram_13_io_r_data : _GEN_12; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_89 = {io_phv_in_data_112,io_phv_in_data_113,io_phv_in_data_114,io_phv_in_data_115,
    io_phv_in_data_116,io_phv_in_data_117,io_phv_in_data_118}; // @[Cat.scala 30:58]
  wire  cs_hit_14 = io_pcie_o_cs == 6'he; // @[outport.scala 31:35]
  wire [63:0] _GEN_14 = cs_hit_14 ? sram_14_io_r_data : _GEN_13; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_95 = {io_phv_in_data_120,io_phv_in_data_121,io_phv_in_data_122,io_phv_in_data_123,
    io_phv_in_data_124,io_phv_in_data_125,io_phv_in_data_126}; // @[Cat.scala 30:58]
  wire  cs_hit_15 = io_pcie_o_cs == 6'hf; // @[outport.scala 31:35]
  wire [63:0] _GEN_15 = cs_hit_15 ? sram_15_io_r_data : _GEN_14; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_101 = {io_phv_in_data_128,io_phv_in_data_129,io_phv_in_data_130,io_phv_in_data_131,
    io_phv_in_data_132,io_phv_in_data_133,io_phv_in_data_134}; // @[Cat.scala 30:58]
  wire  cs_hit_16 = io_pcie_o_cs == 6'h10; // @[outport.scala 31:35]
  wire [63:0] _GEN_16 = cs_hit_16 ? sram_16_io_r_data : _GEN_15; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_107 = {io_phv_in_data_136,io_phv_in_data_137,io_phv_in_data_138,io_phv_in_data_139,
    io_phv_in_data_140,io_phv_in_data_141,io_phv_in_data_142}; // @[Cat.scala 30:58]
  wire  cs_hit_17 = io_pcie_o_cs == 6'h11; // @[outport.scala 31:35]
  wire [63:0] _GEN_17 = cs_hit_17 ? sram_17_io_r_data : _GEN_16; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_113 = {io_phv_in_data_144,io_phv_in_data_145,io_phv_in_data_146,io_phv_in_data_147,
    io_phv_in_data_148,io_phv_in_data_149,io_phv_in_data_150}; // @[Cat.scala 30:58]
  wire  cs_hit_18 = io_pcie_o_cs == 6'h12; // @[outport.scala 31:35]
  wire [63:0] _GEN_18 = cs_hit_18 ? sram_18_io_r_data : _GEN_17; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_119 = {io_phv_in_data_152,io_phv_in_data_153,io_phv_in_data_154,io_phv_in_data_155,
    io_phv_in_data_156,io_phv_in_data_157,io_phv_in_data_158}; // @[Cat.scala 30:58]
  wire  cs_hit_19 = io_pcie_o_cs == 6'h13; // @[outport.scala 31:35]
  wire [63:0] _GEN_19 = cs_hit_19 ? sram_19_io_r_data : _GEN_18; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_125 = {io_phv_in_data_160,io_phv_in_data_161,io_phv_in_data_162,io_phv_in_data_163,
    io_phv_in_data_164,io_phv_in_data_165,io_phv_in_data_166}; // @[Cat.scala 30:58]
  wire  cs_hit_20 = io_pcie_o_cs == 6'h14; // @[outport.scala 31:35]
  wire [63:0] _GEN_20 = cs_hit_20 ? sram_20_io_r_data : _GEN_19; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_131 = {io_phv_in_data_168,io_phv_in_data_169,io_phv_in_data_170,io_phv_in_data_171,
    io_phv_in_data_172,io_phv_in_data_173,io_phv_in_data_174}; // @[Cat.scala 30:58]
  wire  cs_hit_21 = io_pcie_o_cs == 6'h15; // @[outport.scala 31:35]
  wire [63:0] _GEN_21 = cs_hit_21 ? sram_21_io_r_data : _GEN_20; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_137 = {io_phv_in_data_176,io_phv_in_data_177,io_phv_in_data_178,io_phv_in_data_179,
    io_phv_in_data_180,io_phv_in_data_181,io_phv_in_data_182}; // @[Cat.scala 30:58]
  wire  cs_hit_22 = io_pcie_o_cs == 6'h16; // @[outport.scala 31:35]
  wire [63:0] _GEN_22 = cs_hit_22 ? sram_22_io_r_data : _GEN_21; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_143 = {io_phv_in_data_184,io_phv_in_data_185,io_phv_in_data_186,io_phv_in_data_187,
    io_phv_in_data_188,io_phv_in_data_189,io_phv_in_data_190}; // @[Cat.scala 30:58]
  wire  cs_hit_23 = io_pcie_o_cs == 6'h17; // @[outport.scala 31:35]
  wire [63:0] _GEN_23 = cs_hit_23 ? sram_23_io_r_data : _GEN_22; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_149 = {io_phv_in_data_192,io_phv_in_data_193,io_phv_in_data_194,io_phv_in_data_195,
    io_phv_in_data_196,io_phv_in_data_197,io_phv_in_data_198}; // @[Cat.scala 30:58]
  wire  cs_hit_24 = io_pcie_o_cs == 6'h18; // @[outport.scala 31:35]
  wire [63:0] _GEN_24 = cs_hit_24 ? sram_24_io_r_data : _GEN_23; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_155 = {io_phv_in_data_200,io_phv_in_data_201,io_phv_in_data_202,io_phv_in_data_203,
    io_phv_in_data_204,io_phv_in_data_205,io_phv_in_data_206}; // @[Cat.scala 30:58]
  wire  cs_hit_25 = io_pcie_o_cs == 6'h19; // @[outport.scala 31:35]
  wire [63:0] _GEN_25 = cs_hit_25 ? sram_25_io_r_data : _GEN_24; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_161 = {io_phv_in_data_208,io_phv_in_data_209,io_phv_in_data_210,io_phv_in_data_211,
    io_phv_in_data_212,io_phv_in_data_213,io_phv_in_data_214}; // @[Cat.scala 30:58]
  wire  cs_hit_26 = io_pcie_o_cs == 6'h1a; // @[outport.scala 31:35]
  wire [63:0] _GEN_26 = cs_hit_26 ? sram_26_io_r_data : _GEN_25; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_167 = {io_phv_in_data_216,io_phv_in_data_217,io_phv_in_data_218,io_phv_in_data_219,
    io_phv_in_data_220,io_phv_in_data_221,io_phv_in_data_222}; // @[Cat.scala 30:58]
  wire  cs_hit_27 = io_pcie_o_cs == 6'h1b; // @[outport.scala 31:35]
  wire [63:0] _GEN_27 = cs_hit_27 ? sram_27_io_r_data : _GEN_26; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_173 = {io_phv_in_data_224,io_phv_in_data_225,io_phv_in_data_226,io_phv_in_data_227,
    io_phv_in_data_228,io_phv_in_data_229,io_phv_in_data_230}; // @[Cat.scala 30:58]
  wire  cs_hit_28 = io_pcie_o_cs == 6'h1c; // @[outport.scala 31:35]
  wire [63:0] _GEN_28 = cs_hit_28 ? sram_28_io_r_data : _GEN_27; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_179 = {io_phv_in_data_232,io_phv_in_data_233,io_phv_in_data_234,io_phv_in_data_235,
    io_phv_in_data_236,io_phv_in_data_237,io_phv_in_data_238}; // @[Cat.scala 30:58]
  wire  cs_hit_29 = io_pcie_o_cs == 6'h1d; // @[outport.scala 31:35]
  wire [63:0] _GEN_29 = cs_hit_29 ? sram_29_io_r_data : _GEN_28; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_185 = {io_phv_in_data_240,io_phv_in_data_241,io_phv_in_data_242,io_phv_in_data_243,
    io_phv_in_data_244,io_phv_in_data_245,io_phv_in_data_246}; // @[Cat.scala 30:58]
  wire  cs_hit_30 = io_pcie_o_cs == 6'h1e; // @[outport.scala 31:35]
  wire [63:0] _GEN_30 = cs_hit_30 ? sram_30_io_r_data : _GEN_29; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_191 = {io_phv_in_data_248,io_phv_in_data_249,io_phv_in_data_250,io_phv_in_data_251,
    io_phv_in_data_252,io_phv_in_data_253,io_phv_in_data_254}; // @[Cat.scala 30:58]
  wire  cs_hit_31 = io_pcie_o_cs == 6'h1f; // @[outport.scala 31:35]
  wire [63:0] _GEN_31 = cs_hit_31 ? sram_31_io_r_data : _GEN_30; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_197 = {io_phv_in_data_256,io_phv_in_data_257,io_phv_in_data_258,io_phv_in_data_259,
    io_phv_in_data_260,io_phv_in_data_261,io_phv_in_data_262}; // @[Cat.scala 30:58]
  wire  cs_hit_32 = io_pcie_o_cs == 6'h20; // @[outport.scala 31:35]
  wire [63:0] _GEN_32 = cs_hit_32 ? sram_32_io_r_data : _GEN_31; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_203 = {io_phv_in_data_264,io_phv_in_data_265,io_phv_in_data_266,io_phv_in_data_267,
    io_phv_in_data_268,io_phv_in_data_269,io_phv_in_data_270}; // @[Cat.scala 30:58]
  wire  cs_hit_33 = io_pcie_o_cs == 6'h21; // @[outport.scala 31:35]
  wire [63:0] _GEN_33 = cs_hit_33 ? sram_33_io_r_data : _GEN_32; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_209 = {io_phv_in_data_272,io_phv_in_data_273,io_phv_in_data_274,io_phv_in_data_275,
    io_phv_in_data_276,io_phv_in_data_277,io_phv_in_data_278}; // @[Cat.scala 30:58]
  wire  cs_hit_34 = io_pcie_o_cs == 6'h22; // @[outport.scala 31:35]
  wire [63:0] _GEN_34 = cs_hit_34 ? sram_34_io_r_data : _GEN_33; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_215 = {io_phv_in_data_280,io_phv_in_data_281,io_phv_in_data_282,io_phv_in_data_283,
    io_phv_in_data_284,io_phv_in_data_285,io_phv_in_data_286}; // @[Cat.scala 30:58]
  wire  cs_hit_35 = io_pcie_o_cs == 6'h23; // @[outport.scala 31:35]
  wire [63:0] _GEN_35 = cs_hit_35 ? sram_35_io_r_data : _GEN_34; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_221 = {io_phv_in_data_288,io_phv_in_data_289,io_phv_in_data_290,io_phv_in_data_291,
    io_phv_in_data_292,io_phv_in_data_293,io_phv_in_data_294}; // @[Cat.scala 30:58]
  wire  cs_hit_36 = io_pcie_o_cs == 6'h24; // @[outport.scala 31:35]
  wire [63:0] _GEN_36 = cs_hit_36 ? sram_36_io_r_data : _GEN_35; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_227 = {io_phv_in_data_296,io_phv_in_data_297,io_phv_in_data_298,io_phv_in_data_299,
    io_phv_in_data_300,io_phv_in_data_301,io_phv_in_data_302}; // @[Cat.scala 30:58]
  wire  cs_hit_37 = io_pcie_o_cs == 6'h25; // @[outport.scala 31:35]
  wire [63:0] _GEN_37 = cs_hit_37 ? sram_37_io_r_data : _GEN_36; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_233 = {io_phv_in_data_304,io_phv_in_data_305,io_phv_in_data_306,io_phv_in_data_307,
    io_phv_in_data_308,io_phv_in_data_309,io_phv_in_data_310}; // @[Cat.scala 30:58]
  wire  cs_hit_38 = io_pcie_o_cs == 6'h26; // @[outport.scala 31:35]
  wire [63:0] _GEN_38 = cs_hit_38 ? sram_38_io_r_data : _GEN_37; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_239 = {io_phv_in_data_312,io_phv_in_data_313,io_phv_in_data_314,io_phv_in_data_315,
    io_phv_in_data_316,io_phv_in_data_317,io_phv_in_data_318}; // @[Cat.scala 30:58]
  wire  cs_hit_39 = io_pcie_o_cs == 6'h27; // @[outport.scala 31:35]
  wire [63:0] _GEN_39 = cs_hit_39 ? sram_39_io_r_data : _GEN_38; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_245 = {io_phv_in_data_320,io_phv_in_data_321,io_phv_in_data_322,io_phv_in_data_323,
    io_phv_in_data_324,io_phv_in_data_325,io_phv_in_data_326}; // @[Cat.scala 30:58]
  wire  cs_hit_40 = io_pcie_o_cs == 6'h28; // @[outport.scala 31:35]
  wire [63:0] _GEN_40 = cs_hit_40 ? sram_40_io_r_data : _GEN_39; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_251 = {io_phv_in_data_328,io_phv_in_data_329,io_phv_in_data_330,io_phv_in_data_331,
    io_phv_in_data_332,io_phv_in_data_333,io_phv_in_data_334}; // @[Cat.scala 30:58]
  wire  cs_hit_41 = io_pcie_o_cs == 6'h29; // @[outport.scala 31:35]
  wire [63:0] _GEN_41 = cs_hit_41 ? sram_41_io_r_data : _GEN_40; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_257 = {io_phv_in_data_336,io_phv_in_data_337,io_phv_in_data_338,io_phv_in_data_339,
    io_phv_in_data_340,io_phv_in_data_341,io_phv_in_data_342}; // @[Cat.scala 30:58]
  wire  cs_hit_42 = io_pcie_o_cs == 6'h2a; // @[outport.scala 31:35]
  wire [63:0] _GEN_42 = cs_hit_42 ? sram_42_io_r_data : _GEN_41; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_263 = {io_phv_in_data_344,io_phv_in_data_345,io_phv_in_data_346,io_phv_in_data_347,
    io_phv_in_data_348,io_phv_in_data_349,io_phv_in_data_350}; // @[Cat.scala 30:58]
  wire  cs_hit_43 = io_pcie_o_cs == 6'h2b; // @[outport.scala 31:35]
  wire [63:0] _GEN_43 = cs_hit_43 ? sram_43_io_r_data : _GEN_42; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_269 = {io_phv_in_data_352,io_phv_in_data_353,io_phv_in_data_354,io_phv_in_data_355,
    io_phv_in_data_356,io_phv_in_data_357,io_phv_in_data_358}; // @[Cat.scala 30:58]
  wire  cs_hit_44 = io_pcie_o_cs == 6'h2c; // @[outport.scala 31:35]
  wire [63:0] _GEN_44 = cs_hit_44 ? sram_44_io_r_data : _GEN_43; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_275 = {io_phv_in_data_360,io_phv_in_data_361,io_phv_in_data_362,io_phv_in_data_363,
    io_phv_in_data_364,io_phv_in_data_365,io_phv_in_data_366}; // @[Cat.scala 30:58]
  wire  cs_hit_45 = io_pcie_o_cs == 6'h2d; // @[outport.scala 31:35]
  wire [63:0] _GEN_45 = cs_hit_45 ? sram_45_io_r_data : _GEN_44; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_281 = {io_phv_in_data_368,io_phv_in_data_369,io_phv_in_data_370,io_phv_in_data_371,
    io_phv_in_data_372,io_phv_in_data_373,io_phv_in_data_374}; // @[Cat.scala 30:58]
  wire  cs_hit_46 = io_pcie_o_cs == 6'h2e; // @[outport.scala 31:35]
  wire [63:0] _GEN_46 = cs_hit_46 ? sram_46_io_r_data : _GEN_45; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_287 = {io_phv_in_data_376,io_phv_in_data_377,io_phv_in_data_378,io_phv_in_data_379,
    io_phv_in_data_380,io_phv_in_data_381,io_phv_in_data_382}; // @[Cat.scala 30:58]
  wire  cs_hit_47 = io_pcie_o_cs == 6'h2f; // @[outport.scala 31:35]
  wire [63:0] _GEN_47 = cs_hit_47 ? sram_47_io_r_data : _GEN_46; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_293 = {io_phv_in_data_384,io_phv_in_data_385,io_phv_in_data_386,io_phv_in_data_387,
    io_phv_in_data_388,io_phv_in_data_389,io_phv_in_data_390}; // @[Cat.scala 30:58]
  wire  cs_hit_48 = io_pcie_o_cs == 6'h30; // @[outport.scala 31:35]
  wire [63:0] _GEN_48 = cs_hit_48 ? sram_48_io_r_data : _GEN_47; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_299 = {io_phv_in_data_392,io_phv_in_data_393,io_phv_in_data_394,io_phv_in_data_395,
    io_phv_in_data_396,io_phv_in_data_397,io_phv_in_data_398}; // @[Cat.scala 30:58]
  wire  cs_hit_49 = io_pcie_o_cs == 6'h31; // @[outport.scala 31:35]
  wire [63:0] _GEN_49 = cs_hit_49 ? sram_49_io_r_data : _GEN_48; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_305 = {io_phv_in_data_400,io_phv_in_data_401,io_phv_in_data_402,io_phv_in_data_403,
    io_phv_in_data_404,io_phv_in_data_405,io_phv_in_data_406}; // @[Cat.scala 30:58]
  wire  cs_hit_50 = io_pcie_o_cs == 6'h32; // @[outport.scala 31:35]
  wire [63:0] _GEN_50 = cs_hit_50 ? sram_50_io_r_data : _GEN_49; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_311 = {io_phv_in_data_408,io_phv_in_data_409,io_phv_in_data_410,io_phv_in_data_411,
    io_phv_in_data_412,io_phv_in_data_413,io_phv_in_data_414}; // @[Cat.scala 30:58]
  wire  cs_hit_51 = io_pcie_o_cs == 6'h33; // @[outport.scala 31:35]
  wire [63:0] _GEN_51 = cs_hit_51 ? sram_51_io_r_data : _GEN_50; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_317 = {io_phv_in_data_416,io_phv_in_data_417,io_phv_in_data_418,io_phv_in_data_419,
    io_phv_in_data_420,io_phv_in_data_421,io_phv_in_data_422}; // @[Cat.scala 30:58]
  wire  cs_hit_52 = io_pcie_o_cs == 6'h34; // @[outport.scala 31:35]
  wire [63:0] _GEN_52 = cs_hit_52 ? sram_52_io_r_data : _GEN_51; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_323 = {io_phv_in_data_424,io_phv_in_data_425,io_phv_in_data_426,io_phv_in_data_427,
    io_phv_in_data_428,io_phv_in_data_429,io_phv_in_data_430}; // @[Cat.scala 30:58]
  wire  cs_hit_53 = io_pcie_o_cs == 6'h35; // @[outport.scala 31:35]
  wire [63:0] _GEN_53 = cs_hit_53 ? sram_53_io_r_data : _GEN_52; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_329 = {io_phv_in_data_432,io_phv_in_data_433,io_phv_in_data_434,io_phv_in_data_435,
    io_phv_in_data_436,io_phv_in_data_437,io_phv_in_data_438}; // @[Cat.scala 30:58]
  wire  cs_hit_54 = io_pcie_o_cs == 6'h36; // @[outport.scala 31:35]
  wire [63:0] _GEN_54 = cs_hit_54 ? sram_54_io_r_data : _GEN_53; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_335 = {io_phv_in_data_440,io_phv_in_data_441,io_phv_in_data_442,io_phv_in_data_443,
    io_phv_in_data_444,io_phv_in_data_445,io_phv_in_data_446}; // @[Cat.scala 30:58]
  wire  cs_hit_55 = io_pcie_o_cs == 6'h37; // @[outport.scala 31:35]
  wire [63:0] _GEN_55 = cs_hit_55 ? sram_55_io_r_data : _GEN_54; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_341 = {io_phv_in_data_448,io_phv_in_data_449,io_phv_in_data_450,io_phv_in_data_451,
    io_phv_in_data_452,io_phv_in_data_453,io_phv_in_data_454}; // @[Cat.scala 30:58]
  wire  cs_hit_56 = io_pcie_o_cs == 6'h38; // @[outport.scala 31:35]
  wire [63:0] _GEN_56 = cs_hit_56 ? sram_56_io_r_data : _GEN_55; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_347 = {io_phv_in_data_456,io_phv_in_data_457,io_phv_in_data_458,io_phv_in_data_459,
    io_phv_in_data_460,io_phv_in_data_461,io_phv_in_data_462}; // @[Cat.scala 30:58]
  wire  cs_hit_57 = io_pcie_o_cs == 6'h39; // @[outport.scala 31:35]
  wire [63:0] _GEN_57 = cs_hit_57 ? sram_57_io_r_data : _GEN_56; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_353 = {io_phv_in_data_464,io_phv_in_data_465,io_phv_in_data_466,io_phv_in_data_467,
    io_phv_in_data_468,io_phv_in_data_469,io_phv_in_data_470}; // @[Cat.scala 30:58]
  wire  cs_hit_58 = io_pcie_o_cs == 6'h3a; // @[outport.scala 31:35]
  wire [63:0] _GEN_58 = cs_hit_58 ? sram_58_io_r_data : _GEN_57; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_359 = {io_phv_in_data_472,io_phv_in_data_473,io_phv_in_data_474,io_phv_in_data_475,
    io_phv_in_data_476,io_phv_in_data_477,io_phv_in_data_478}; // @[Cat.scala 30:58]
  wire  cs_hit_59 = io_pcie_o_cs == 6'h3b; // @[outport.scala 31:35]
  wire [63:0] _GEN_59 = cs_hit_59 ? sram_59_io_r_data : _GEN_58; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_365 = {io_phv_in_data_480,io_phv_in_data_481,io_phv_in_data_482,io_phv_in_data_483,
    io_phv_in_data_484,io_phv_in_data_485,io_phv_in_data_486}; // @[Cat.scala 30:58]
  wire  cs_hit_60 = io_pcie_o_cs == 6'h3c; // @[outport.scala 31:35]
  wire [63:0] _GEN_60 = cs_hit_60 ? sram_60_io_r_data : _GEN_59; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_371 = {io_phv_in_data_488,io_phv_in_data_489,io_phv_in_data_490,io_phv_in_data_491,
    io_phv_in_data_492,io_phv_in_data_493,io_phv_in_data_494}; // @[Cat.scala 30:58]
  wire  cs_hit_61 = io_pcie_o_cs == 6'h3d; // @[outport.scala 31:35]
  wire [63:0] _GEN_61 = cs_hit_61 ? sram_61_io_r_data : _GEN_60; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_377 = {io_phv_in_data_496,io_phv_in_data_497,io_phv_in_data_498,io_phv_in_data_499,
    io_phv_in_data_500,io_phv_in_data_501,io_phv_in_data_502}; // @[Cat.scala 30:58]
  wire  cs_hit_62 = io_pcie_o_cs == 6'h3e; // @[outport.scala 31:35]
  wire [63:0] _GEN_62 = cs_hit_62 ? sram_62_io_r_data : _GEN_61; // @[outport.scala 34:23 outport.scala 35:31]
  wire [55:0] exe_io_w_data_hi_383 = {io_phv_in_data_504,io_phv_in_data_505,io_phv_in_data_506,io_phv_in_data_507,
    io_phv_in_data_508,io_phv_in_data_509,io_phv_in_data_510}; // @[Cat.scala 30:58]
  wire  cs_hit_63 = io_pcie_o_cs == 6'h3f; // @[outport.scala 31:35]
  SRAM sram_0 ( // @[outport.scala 23:25]
    .clock(sram_0_clock),
    .io_w_en(sram_0_io_w_en),
    .io_w_addr(sram_0_io_w_addr),
    .io_w_data(sram_0_io_w_data),
    .io_r_en(sram_0_io_r_en),
    .io_r_addr(sram_0_io_r_addr),
    .io_r_data(sram_0_io_r_data)
  );
  SRAM sram_1 ( // @[outport.scala 23:25]
    .clock(sram_1_clock),
    .io_w_en(sram_1_io_w_en),
    .io_w_addr(sram_1_io_w_addr),
    .io_w_data(sram_1_io_w_data),
    .io_r_en(sram_1_io_r_en),
    .io_r_addr(sram_1_io_r_addr),
    .io_r_data(sram_1_io_r_data)
  );
  SRAM sram_2 ( // @[outport.scala 23:25]
    .clock(sram_2_clock),
    .io_w_en(sram_2_io_w_en),
    .io_w_addr(sram_2_io_w_addr),
    .io_w_data(sram_2_io_w_data),
    .io_r_en(sram_2_io_r_en),
    .io_r_addr(sram_2_io_r_addr),
    .io_r_data(sram_2_io_r_data)
  );
  SRAM sram_3 ( // @[outport.scala 23:25]
    .clock(sram_3_clock),
    .io_w_en(sram_3_io_w_en),
    .io_w_addr(sram_3_io_w_addr),
    .io_w_data(sram_3_io_w_data),
    .io_r_en(sram_3_io_r_en),
    .io_r_addr(sram_3_io_r_addr),
    .io_r_data(sram_3_io_r_data)
  );
  SRAM sram_4 ( // @[outport.scala 23:25]
    .clock(sram_4_clock),
    .io_w_en(sram_4_io_w_en),
    .io_w_addr(sram_4_io_w_addr),
    .io_w_data(sram_4_io_w_data),
    .io_r_en(sram_4_io_r_en),
    .io_r_addr(sram_4_io_r_addr),
    .io_r_data(sram_4_io_r_data)
  );
  SRAM sram_5 ( // @[outport.scala 23:25]
    .clock(sram_5_clock),
    .io_w_en(sram_5_io_w_en),
    .io_w_addr(sram_5_io_w_addr),
    .io_w_data(sram_5_io_w_data),
    .io_r_en(sram_5_io_r_en),
    .io_r_addr(sram_5_io_r_addr),
    .io_r_data(sram_5_io_r_data)
  );
  SRAM sram_6 ( // @[outport.scala 23:25]
    .clock(sram_6_clock),
    .io_w_en(sram_6_io_w_en),
    .io_w_addr(sram_6_io_w_addr),
    .io_w_data(sram_6_io_w_data),
    .io_r_en(sram_6_io_r_en),
    .io_r_addr(sram_6_io_r_addr),
    .io_r_data(sram_6_io_r_data)
  );
  SRAM sram_7 ( // @[outport.scala 23:25]
    .clock(sram_7_clock),
    .io_w_en(sram_7_io_w_en),
    .io_w_addr(sram_7_io_w_addr),
    .io_w_data(sram_7_io_w_data),
    .io_r_en(sram_7_io_r_en),
    .io_r_addr(sram_7_io_r_addr),
    .io_r_data(sram_7_io_r_data)
  );
  SRAM sram_8 ( // @[outport.scala 23:25]
    .clock(sram_8_clock),
    .io_w_en(sram_8_io_w_en),
    .io_w_addr(sram_8_io_w_addr),
    .io_w_data(sram_8_io_w_data),
    .io_r_en(sram_8_io_r_en),
    .io_r_addr(sram_8_io_r_addr),
    .io_r_data(sram_8_io_r_data)
  );
  SRAM sram_9 ( // @[outport.scala 23:25]
    .clock(sram_9_clock),
    .io_w_en(sram_9_io_w_en),
    .io_w_addr(sram_9_io_w_addr),
    .io_w_data(sram_9_io_w_data),
    .io_r_en(sram_9_io_r_en),
    .io_r_addr(sram_9_io_r_addr),
    .io_r_data(sram_9_io_r_data)
  );
  SRAM sram_10 ( // @[outport.scala 23:25]
    .clock(sram_10_clock),
    .io_w_en(sram_10_io_w_en),
    .io_w_addr(sram_10_io_w_addr),
    .io_w_data(sram_10_io_w_data),
    .io_r_en(sram_10_io_r_en),
    .io_r_addr(sram_10_io_r_addr),
    .io_r_data(sram_10_io_r_data)
  );
  SRAM sram_11 ( // @[outport.scala 23:25]
    .clock(sram_11_clock),
    .io_w_en(sram_11_io_w_en),
    .io_w_addr(sram_11_io_w_addr),
    .io_w_data(sram_11_io_w_data),
    .io_r_en(sram_11_io_r_en),
    .io_r_addr(sram_11_io_r_addr),
    .io_r_data(sram_11_io_r_data)
  );
  SRAM sram_12 ( // @[outport.scala 23:25]
    .clock(sram_12_clock),
    .io_w_en(sram_12_io_w_en),
    .io_w_addr(sram_12_io_w_addr),
    .io_w_data(sram_12_io_w_data),
    .io_r_en(sram_12_io_r_en),
    .io_r_addr(sram_12_io_r_addr),
    .io_r_data(sram_12_io_r_data)
  );
  SRAM sram_13 ( // @[outport.scala 23:25]
    .clock(sram_13_clock),
    .io_w_en(sram_13_io_w_en),
    .io_w_addr(sram_13_io_w_addr),
    .io_w_data(sram_13_io_w_data),
    .io_r_en(sram_13_io_r_en),
    .io_r_addr(sram_13_io_r_addr),
    .io_r_data(sram_13_io_r_data)
  );
  SRAM sram_14 ( // @[outport.scala 23:25]
    .clock(sram_14_clock),
    .io_w_en(sram_14_io_w_en),
    .io_w_addr(sram_14_io_w_addr),
    .io_w_data(sram_14_io_w_data),
    .io_r_en(sram_14_io_r_en),
    .io_r_addr(sram_14_io_r_addr),
    .io_r_data(sram_14_io_r_data)
  );
  SRAM sram_15 ( // @[outport.scala 23:25]
    .clock(sram_15_clock),
    .io_w_en(sram_15_io_w_en),
    .io_w_addr(sram_15_io_w_addr),
    .io_w_data(sram_15_io_w_data),
    .io_r_en(sram_15_io_r_en),
    .io_r_addr(sram_15_io_r_addr),
    .io_r_data(sram_15_io_r_data)
  );
  SRAM sram_16 ( // @[outport.scala 23:25]
    .clock(sram_16_clock),
    .io_w_en(sram_16_io_w_en),
    .io_w_addr(sram_16_io_w_addr),
    .io_w_data(sram_16_io_w_data),
    .io_r_en(sram_16_io_r_en),
    .io_r_addr(sram_16_io_r_addr),
    .io_r_data(sram_16_io_r_data)
  );
  SRAM sram_17 ( // @[outport.scala 23:25]
    .clock(sram_17_clock),
    .io_w_en(sram_17_io_w_en),
    .io_w_addr(sram_17_io_w_addr),
    .io_w_data(sram_17_io_w_data),
    .io_r_en(sram_17_io_r_en),
    .io_r_addr(sram_17_io_r_addr),
    .io_r_data(sram_17_io_r_data)
  );
  SRAM sram_18 ( // @[outport.scala 23:25]
    .clock(sram_18_clock),
    .io_w_en(sram_18_io_w_en),
    .io_w_addr(sram_18_io_w_addr),
    .io_w_data(sram_18_io_w_data),
    .io_r_en(sram_18_io_r_en),
    .io_r_addr(sram_18_io_r_addr),
    .io_r_data(sram_18_io_r_data)
  );
  SRAM sram_19 ( // @[outport.scala 23:25]
    .clock(sram_19_clock),
    .io_w_en(sram_19_io_w_en),
    .io_w_addr(sram_19_io_w_addr),
    .io_w_data(sram_19_io_w_data),
    .io_r_en(sram_19_io_r_en),
    .io_r_addr(sram_19_io_r_addr),
    .io_r_data(sram_19_io_r_data)
  );
  SRAM sram_20 ( // @[outport.scala 23:25]
    .clock(sram_20_clock),
    .io_w_en(sram_20_io_w_en),
    .io_w_addr(sram_20_io_w_addr),
    .io_w_data(sram_20_io_w_data),
    .io_r_en(sram_20_io_r_en),
    .io_r_addr(sram_20_io_r_addr),
    .io_r_data(sram_20_io_r_data)
  );
  SRAM sram_21 ( // @[outport.scala 23:25]
    .clock(sram_21_clock),
    .io_w_en(sram_21_io_w_en),
    .io_w_addr(sram_21_io_w_addr),
    .io_w_data(sram_21_io_w_data),
    .io_r_en(sram_21_io_r_en),
    .io_r_addr(sram_21_io_r_addr),
    .io_r_data(sram_21_io_r_data)
  );
  SRAM sram_22 ( // @[outport.scala 23:25]
    .clock(sram_22_clock),
    .io_w_en(sram_22_io_w_en),
    .io_w_addr(sram_22_io_w_addr),
    .io_w_data(sram_22_io_w_data),
    .io_r_en(sram_22_io_r_en),
    .io_r_addr(sram_22_io_r_addr),
    .io_r_data(sram_22_io_r_data)
  );
  SRAM sram_23 ( // @[outport.scala 23:25]
    .clock(sram_23_clock),
    .io_w_en(sram_23_io_w_en),
    .io_w_addr(sram_23_io_w_addr),
    .io_w_data(sram_23_io_w_data),
    .io_r_en(sram_23_io_r_en),
    .io_r_addr(sram_23_io_r_addr),
    .io_r_data(sram_23_io_r_data)
  );
  SRAM sram_24 ( // @[outport.scala 23:25]
    .clock(sram_24_clock),
    .io_w_en(sram_24_io_w_en),
    .io_w_addr(sram_24_io_w_addr),
    .io_w_data(sram_24_io_w_data),
    .io_r_en(sram_24_io_r_en),
    .io_r_addr(sram_24_io_r_addr),
    .io_r_data(sram_24_io_r_data)
  );
  SRAM sram_25 ( // @[outport.scala 23:25]
    .clock(sram_25_clock),
    .io_w_en(sram_25_io_w_en),
    .io_w_addr(sram_25_io_w_addr),
    .io_w_data(sram_25_io_w_data),
    .io_r_en(sram_25_io_r_en),
    .io_r_addr(sram_25_io_r_addr),
    .io_r_data(sram_25_io_r_data)
  );
  SRAM sram_26 ( // @[outport.scala 23:25]
    .clock(sram_26_clock),
    .io_w_en(sram_26_io_w_en),
    .io_w_addr(sram_26_io_w_addr),
    .io_w_data(sram_26_io_w_data),
    .io_r_en(sram_26_io_r_en),
    .io_r_addr(sram_26_io_r_addr),
    .io_r_data(sram_26_io_r_data)
  );
  SRAM sram_27 ( // @[outport.scala 23:25]
    .clock(sram_27_clock),
    .io_w_en(sram_27_io_w_en),
    .io_w_addr(sram_27_io_w_addr),
    .io_w_data(sram_27_io_w_data),
    .io_r_en(sram_27_io_r_en),
    .io_r_addr(sram_27_io_r_addr),
    .io_r_data(sram_27_io_r_data)
  );
  SRAM sram_28 ( // @[outport.scala 23:25]
    .clock(sram_28_clock),
    .io_w_en(sram_28_io_w_en),
    .io_w_addr(sram_28_io_w_addr),
    .io_w_data(sram_28_io_w_data),
    .io_r_en(sram_28_io_r_en),
    .io_r_addr(sram_28_io_r_addr),
    .io_r_data(sram_28_io_r_data)
  );
  SRAM sram_29 ( // @[outport.scala 23:25]
    .clock(sram_29_clock),
    .io_w_en(sram_29_io_w_en),
    .io_w_addr(sram_29_io_w_addr),
    .io_w_data(sram_29_io_w_data),
    .io_r_en(sram_29_io_r_en),
    .io_r_addr(sram_29_io_r_addr),
    .io_r_data(sram_29_io_r_data)
  );
  SRAM sram_30 ( // @[outport.scala 23:25]
    .clock(sram_30_clock),
    .io_w_en(sram_30_io_w_en),
    .io_w_addr(sram_30_io_w_addr),
    .io_w_data(sram_30_io_w_data),
    .io_r_en(sram_30_io_r_en),
    .io_r_addr(sram_30_io_r_addr),
    .io_r_data(sram_30_io_r_data)
  );
  SRAM sram_31 ( // @[outport.scala 23:25]
    .clock(sram_31_clock),
    .io_w_en(sram_31_io_w_en),
    .io_w_addr(sram_31_io_w_addr),
    .io_w_data(sram_31_io_w_data),
    .io_r_en(sram_31_io_r_en),
    .io_r_addr(sram_31_io_r_addr),
    .io_r_data(sram_31_io_r_data)
  );
  SRAM sram_32 ( // @[outport.scala 23:25]
    .clock(sram_32_clock),
    .io_w_en(sram_32_io_w_en),
    .io_w_addr(sram_32_io_w_addr),
    .io_w_data(sram_32_io_w_data),
    .io_r_en(sram_32_io_r_en),
    .io_r_addr(sram_32_io_r_addr),
    .io_r_data(sram_32_io_r_data)
  );
  SRAM sram_33 ( // @[outport.scala 23:25]
    .clock(sram_33_clock),
    .io_w_en(sram_33_io_w_en),
    .io_w_addr(sram_33_io_w_addr),
    .io_w_data(sram_33_io_w_data),
    .io_r_en(sram_33_io_r_en),
    .io_r_addr(sram_33_io_r_addr),
    .io_r_data(sram_33_io_r_data)
  );
  SRAM sram_34 ( // @[outport.scala 23:25]
    .clock(sram_34_clock),
    .io_w_en(sram_34_io_w_en),
    .io_w_addr(sram_34_io_w_addr),
    .io_w_data(sram_34_io_w_data),
    .io_r_en(sram_34_io_r_en),
    .io_r_addr(sram_34_io_r_addr),
    .io_r_data(sram_34_io_r_data)
  );
  SRAM sram_35 ( // @[outport.scala 23:25]
    .clock(sram_35_clock),
    .io_w_en(sram_35_io_w_en),
    .io_w_addr(sram_35_io_w_addr),
    .io_w_data(sram_35_io_w_data),
    .io_r_en(sram_35_io_r_en),
    .io_r_addr(sram_35_io_r_addr),
    .io_r_data(sram_35_io_r_data)
  );
  SRAM sram_36 ( // @[outport.scala 23:25]
    .clock(sram_36_clock),
    .io_w_en(sram_36_io_w_en),
    .io_w_addr(sram_36_io_w_addr),
    .io_w_data(sram_36_io_w_data),
    .io_r_en(sram_36_io_r_en),
    .io_r_addr(sram_36_io_r_addr),
    .io_r_data(sram_36_io_r_data)
  );
  SRAM sram_37 ( // @[outport.scala 23:25]
    .clock(sram_37_clock),
    .io_w_en(sram_37_io_w_en),
    .io_w_addr(sram_37_io_w_addr),
    .io_w_data(sram_37_io_w_data),
    .io_r_en(sram_37_io_r_en),
    .io_r_addr(sram_37_io_r_addr),
    .io_r_data(sram_37_io_r_data)
  );
  SRAM sram_38 ( // @[outport.scala 23:25]
    .clock(sram_38_clock),
    .io_w_en(sram_38_io_w_en),
    .io_w_addr(sram_38_io_w_addr),
    .io_w_data(sram_38_io_w_data),
    .io_r_en(sram_38_io_r_en),
    .io_r_addr(sram_38_io_r_addr),
    .io_r_data(sram_38_io_r_data)
  );
  SRAM sram_39 ( // @[outport.scala 23:25]
    .clock(sram_39_clock),
    .io_w_en(sram_39_io_w_en),
    .io_w_addr(sram_39_io_w_addr),
    .io_w_data(sram_39_io_w_data),
    .io_r_en(sram_39_io_r_en),
    .io_r_addr(sram_39_io_r_addr),
    .io_r_data(sram_39_io_r_data)
  );
  SRAM sram_40 ( // @[outport.scala 23:25]
    .clock(sram_40_clock),
    .io_w_en(sram_40_io_w_en),
    .io_w_addr(sram_40_io_w_addr),
    .io_w_data(sram_40_io_w_data),
    .io_r_en(sram_40_io_r_en),
    .io_r_addr(sram_40_io_r_addr),
    .io_r_data(sram_40_io_r_data)
  );
  SRAM sram_41 ( // @[outport.scala 23:25]
    .clock(sram_41_clock),
    .io_w_en(sram_41_io_w_en),
    .io_w_addr(sram_41_io_w_addr),
    .io_w_data(sram_41_io_w_data),
    .io_r_en(sram_41_io_r_en),
    .io_r_addr(sram_41_io_r_addr),
    .io_r_data(sram_41_io_r_data)
  );
  SRAM sram_42 ( // @[outport.scala 23:25]
    .clock(sram_42_clock),
    .io_w_en(sram_42_io_w_en),
    .io_w_addr(sram_42_io_w_addr),
    .io_w_data(sram_42_io_w_data),
    .io_r_en(sram_42_io_r_en),
    .io_r_addr(sram_42_io_r_addr),
    .io_r_data(sram_42_io_r_data)
  );
  SRAM sram_43 ( // @[outport.scala 23:25]
    .clock(sram_43_clock),
    .io_w_en(sram_43_io_w_en),
    .io_w_addr(sram_43_io_w_addr),
    .io_w_data(sram_43_io_w_data),
    .io_r_en(sram_43_io_r_en),
    .io_r_addr(sram_43_io_r_addr),
    .io_r_data(sram_43_io_r_data)
  );
  SRAM sram_44 ( // @[outport.scala 23:25]
    .clock(sram_44_clock),
    .io_w_en(sram_44_io_w_en),
    .io_w_addr(sram_44_io_w_addr),
    .io_w_data(sram_44_io_w_data),
    .io_r_en(sram_44_io_r_en),
    .io_r_addr(sram_44_io_r_addr),
    .io_r_data(sram_44_io_r_data)
  );
  SRAM sram_45 ( // @[outport.scala 23:25]
    .clock(sram_45_clock),
    .io_w_en(sram_45_io_w_en),
    .io_w_addr(sram_45_io_w_addr),
    .io_w_data(sram_45_io_w_data),
    .io_r_en(sram_45_io_r_en),
    .io_r_addr(sram_45_io_r_addr),
    .io_r_data(sram_45_io_r_data)
  );
  SRAM sram_46 ( // @[outport.scala 23:25]
    .clock(sram_46_clock),
    .io_w_en(sram_46_io_w_en),
    .io_w_addr(sram_46_io_w_addr),
    .io_w_data(sram_46_io_w_data),
    .io_r_en(sram_46_io_r_en),
    .io_r_addr(sram_46_io_r_addr),
    .io_r_data(sram_46_io_r_data)
  );
  SRAM sram_47 ( // @[outport.scala 23:25]
    .clock(sram_47_clock),
    .io_w_en(sram_47_io_w_en),
    .io_w_addr(sram_47_io_w_addr),
    .io_w_data(sram_47_io_w_data),
    .io_r_en(sram_47_io_r_en),
    .io_r_addr(sram_47_io_r_addr),
    .io_r_data(sram_47_io_r_data)
  );
  SRAM sram_48 ( // @[outport.scala 23:25]
    .clock(sram_48_clock),
    .io_w_en(sram_48_io_w_en),
    .io_w_addr(sram_48_io_w_addr),
    .io_w_data(sram_48_io_w_data),
    .io_r_en(sram_48_io_r_en),
    .io_r_addr(sram_48_io_r_addr),
    .io_r_data(sram_48_io_r_data)
  );
  SRAM sram_49 ( // @[outport.scala 23:25]
    .clock(sram_49_clock),
    .io_w_en(sram_49_io_w_en),
    .io_w_addr(sram_49_io_w_addr),
    .io_w_data(sram_49_io_w_data),
    .io_r_en(sram_49_io_r_en),
    .io_r_addr(sram_49_io_r_addr),
    .io_r_data(sram_49_io_r_data)
  );
  SRAM sram_50 ( // @[outport.scala 23:25]
    .clock(sram_50_clock),
    .io_w_en(sram_50_io_w_en),
    .io_w_addr(sram_50_io_w_addr),
    .io_w_data(sram_50_io_w_data),
    .io_r_en(sram_50_io_r_en),
    .io_r_addr(sram_50_io_r_addr),
    .io_r_data(sram_50_io_r_data)
  );
  SRAM sram_51 ( // @[outport.scala 23:25]
    .clock(sram_51_clock),
    .io_w_en(sram_51_io_w_en),
    .io_w_addr(sram_51_io_w_addr),
    .io_w_data(sram_51_io_w_data),
    .io_r_en(sram_51_io_r_en),
    .io_r_addr(sram_51_io_r_addr),
    .io_r_data(sram_51_io_r_data)
  );
  SRAM sram_52 ( // @[outport.scala 23:25]
    .clock(sram_52_clock),
    .io_w_en(sram_52_io_w_en),
    .io_w_addr(sram_52_io_w_addr),
    .io_w_data(sram_52_io_w_data),
    .io_r_en(sram_52_io_r_en),
    .io_r_addr(sram_52_io_r_addr),
    .io_r_data(sram_52_io_r_data)
  );
  SRAM sram_53 ( // @[outport.scala 23:25]
    .clock(sram_53_clock),
    .io_w_en(sram_53_io_w_en),
    .io_w_addr(sram_53_io_w_addr),
    .io_w_data(sram_53_io_w_data),
    .io_r_en(sram_53_io_r_en),
    .io_r_addr(sram_53_io_r_addr),
    .io_r_data(sram_53_io_r_data)
  );
  SRAM sram_54 ( // @[outport.scala 23:25]
    .clock(sram_54_clock),
    .io_w_en(sram_54_io_w_en),
    .io_w_addr(sram_54_io_w_addr),
    .io_w_data(sram_54_io_w_data),
    .io_r_en(sram_54_io_r_en),
    .io_r_addr(sram_54_io_r_addr),
    .io_r_data(sram_54_io_r_data)
  );
  SRAM sram_55 ( // @[outport.scala 23:25]
    .clock(sram_55_clock),
    .io_w_en(sram_55_io_w_en),
    .io_w_addr(sram_55_io_w_addr),
    .io_w_data(sram_55_io_w_data),
    .io_r_en(sram_55_io_r_en),
    .io_r_addr(sram_55_io_r_addr),
    .io_r_data(sram_55_io_r_data)
  );
  SRAM sram_56 ( // @[outport.scala 23:25]
    .clock(sram_56_clock),
    .io_w_en(sram_56_io_w_en),
    .io_w_addr(sram_56_io_w_addr),
    .io_w_data(sram_56_io_w_data),
    .io_r_en(sram_56_io_r_en),
    .io_r_addr(sram_56_io_r_addr),
    .io_r_data(sram_56_io_r_data)
  );
  SRAM sram_57 ( // @[outport.scala 23:25]
    .clock(sram_57_clock),
    .io_w_en(sram_57_io_w_en),
    .io_w_addr(sram_57_io_w_addr),
    .io_w_data(sram_57_io_w_data),
    .io_r_en(sram_57_io_r_en),
    .io_r_addr(sram_57_io_r_addr),
    .io_r_data(sram_57_io_r_data)
  );
  SRAM sram_58 ( // @[outport.scala 23:25]
    .clock(sram_58_clock),
    .io_w_en(sram_58_io_w_en),
    .io_w_addr(sram_58_io_w_addr),
    .io_w_data(sram_58_io_w_data),
    .io_r_en(sram_58_io_r_en),
    .io_r_addr(sram_58_io_r_addr),
    .io_r_data(sram_58_io_r_data)
  );
  SRAM sram_59 ( // @[outport.scala 23:25]
    .clock(sram_59_clock),
    .io_w_en(sram_59_io_w_en),
    .io_w_addr(sram_59_io_w_addr),
    .io_w_data(sram_59_io_w_data),
    .io_r_en(sram_59_io_r_en),
    .io_r_addr(sram_59_io_r_addr),
    .io_r_data(sram_59_io_r_data)
  );
  SRAM sram_60 ( // @[outport.scala 23:25]
    .clock(sram_60_clock),
    .io_w_en(sram_60_io_w_en),
    .io_w_addr(sram_60_io_w_addr),
    .io_w_data(sram_60_io_w_data),
    .io_r_en(sram_60_io_r_en),
    .io_r_addr(sram_60_io_r_addr),
    .io_r_data(sram_60_io_r_data)
  );
  SRAM sram_61 ( // @[outport.scala 23:25]
    .clock(sram_61_clock),
    .io_w_en(sram_61_io_w_en),
    .io_w_addr(sram_61_io_w_addr),
    .io_w_data(sram_61_io_w_data),
    .io_r_en(sram_61_io_r_en),
    .io_r_addr(sram_61_io_r_addr),
    .io_r_data(sram_61_io_r_data)
  );
  SRAM sram_62 ( // @[outport.scala 23:25]
    .clock(sram_62_clock),
    .io_w_en(sram_62_io_w_en),
    .io_w_addr(sram_62_io_w_addr),
    .io_w_data(sram_62_io_w_data),
    .io_r_en(sram_62_io_r_en),
    .io_r_addr(sram_62_io_r_addr),
    .io_r_data(sram_62_io_r_data)
  );
  SRAM sram_63 ( // @[outport.scala 23:25]
    .clock(sram_63_clock),
    .io_w_en(sram_63_io_w_en),
    .io_w_addr(sram_63_io_w_addr),
    .io_w_data(sram_63_io_w_data),
    .io_r_en(sram_63_io_r_en),
    .io_r_addr(sram_63_io_r_addr),
    .io_r_data(sram_63_io_r_data)
  );
  assign io_pcie_o_r_data = cs_hit_63 ? sram_63_io_r_data : _GEN_62; // @[outport.scala 34:23 outport.scala 35:31]
  assign sram_0_clock = clock;
  assign sram_0_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_0_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_0_io_w_data = {exe_io_w_data_hi_5,io_phv_in_data_7}; // @[Cat.scala 30:58]
  assign sram_0_io_r_en = io_pcie_o_r_en & cs_hit; // @[outport.scala 32:42]
  assign sram_0_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_1_clock = clock;
  assign sram_1_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_1_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_1_io_w_data = {exe_io_w_data_hi_11,io_phv_in_data_15}; // @[Cat.scala 30:58]
  assign sram_1_io_r_en = io_pcie_o_r_en & cs_hit_1; // @[outport.scala 32:42]
  assign sram_1_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_2_clock = clock;
  assign sram_2_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_2_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_2_io_w_data = {exe_io_w_data_hi_17,io_phv_in_data_23}; // @[Cat.scala 30:58]
  assign sram_2_io_r_en = io_pcie_o_r_en & cs_hit_2; // @[outport.scala 32:42]
  assign sram_2_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_3_clock = clock;
  assign sram_3_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_3_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_3_io_w_data = {exe_io_w_data_hi_23,io_phv_in_data_31}; // @[Cat.scala 30:58]
  assign sram_3_io_r_en = io_pcie_o_r_en & cs_hit_3; // @[outport.scala 32:42]
  assign sram_3_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_4_clock = clock;
  assign sram_4_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_4_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_4_io_w_data = {exe_io_w_data_hi_29,io_phv_in_data_39}; // @[Cat.scala 30:58]
  assign sram_4_io_r_en = io_pcie_o_r_en & cs_hit_4; // @[outport.scala 32:42]
  assign sram_4_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_5_clock = clock;
  assign sram_5_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_5_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_5_io_w_data = {exe_io_w_data_hi_35,io_phv_in_data_47}; // @[Cat.scala 30:58]
  assign sram_5_io_r_en = io_pcie_o_r_en & cs_hit_5; // @[outport.scala 32:42]
  assign sram_5_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_6_clock = clock;
  assign sram_6_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_6_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_6_io_w_data = {exe_io_w_data_hi_41,io_phv_in_data_55}; // @[Cat.scala 30:58]
  assign sram_6_io_r_en = io_pcie_o_r_en & cs_hit_6; // @[outport.scala 32:42]
  assign sram_6_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_7_clock = clock;
  assign sram_7_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_7_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_7_io_w_data = {exe_io_w_data_hi_47,io_phv_in_data_63}; // @[Cat.scala 30:58]
  assign sram_7_io_r_en = io_pcie_o_r_en & cs_hit_7; // @[outport.scala 32:42]
  assign sram_7_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_8_clock = clock;
  assign sram_8_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_8_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_8_io_w_data = {exe_io_w_data_hi_53,io_phv_in_data_71}; // @[Cat.scala 30:58]
  assign sram_8_io_r_en = io_pcie_o_r_en & cs_hit_8; // @[outport.scala 32:42]
  assign sram_8_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_9_clock = clock;
  assign sram_9_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_9_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_9_io_w_data = {exe_io_w_data_hi_59,io_phv_in_data_79}; // @[Cat.scala 30:58]
  assign sram_9_io_r_en = io_pcie_o_r_en & cs_hit_9; // @[outport.scala 32:42]
  assign sram_9_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_10_clock = clock;
  assign sram_10_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_10_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_10_io_w_data = {exe_io_w_data_hi_65,io_phv_in_data_87}; // @[Cat.scala 30:58]
  assign sram_10_io_r_en = io_pcie_o_r_en & cs_hit_10; // @[outport.scala 32:42]
  assign sram_10_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_11_clock = clock;
  assign sram_11_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_11_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_11_io_w_data = {exe_io_w_data_hi_71,io_phv_in_data_95}; // @[Cat.scala 30:58]
  assign sram_11_io_r_en = io_pcie_o_r_en & cs_hit_11; // @[outport.scala 32:42]
  assign sram_11_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_12_clock = clock;
  assign sram_12_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_12_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_12_io_w_data = {exe_io_w_data_hi_77,io_phv_in_data_103}; // @[Cat.scala 30:58]
  assign sram_12_io_r_en = io_pcie_o_r_en & cs_hit_12; // @[outport.scala 32:42]
  assign sram_12_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_13_clock = clock;
  assign sram_13_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_13_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_13_io_w_data = {exe_io_w_data_hi_83,io_phv_in_data_111}; // @[Cat.scala 30:58]
  assign sram_13_io_r_en = io_pcie_o_r_en & cs_hit_13; // @[outport.scala 32:42]
  assign sram_13_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_14_clock = clock;
  assign sram_14_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_14_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_14_io_w_data = {exe_io_w_data_hi_89,io_phv_in_data_119}; // @[Cat.scala 30:58]
  assign sram_14_io_r_en = io_pcie_o_r_en & cs_hit_14; // @[outport.scala 32:42]
  assign sram_14_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_15_clock = clock;
  assign sram_15_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_15_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_15_io_w_data = {exe_io_w_data_hi_95,io_phv_in_data_127}; // @[Cat.scala 30:58]
  assign sram_15_io_r_en = io_pcie_o_r_en & cs_hit_15; // @[outport.scala 32:42]
  assign sram_15_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_16_clock = clock;
  assign sram_16_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_16_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_16_io_w_data = {exe_io_w_data_hi_101,io_phv_in_data_135}; // @[Cat.scala 30:58]
  assign sram_16_io_r_en = io_pcie_o_r_en & cs_hit_16; // @[outport.scala 32:42]
  assign sram_16_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_17_clock = clock;
  assign sram_17_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_17_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_17_io_w_data = {exe_io_w_data_hi_107,io_phv_in_data_143}; // @[Cat.scala 30:58]
  assign sram_17_io_r_en = io_pcie_o_r_en & cs_hit_17; // @[outport.scala 32:42]
  assign sram_17_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_18_clock = clock;
  assign sram_18_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_18_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_18_io_w_data = {exe_io_w_data_hi_113,io_phv_in_data_151}; // @[Cat.scala 30:58]
  assign sram_18_io_r_en = io_pcie_o_r_en & cs_hit_18; // @[outport.scala 32:42]
  assign sram_18_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_19_clock = clock;
  assign sram_19_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_19_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_19_io_w_data = {exe_io_w_data_hi_119,io_phv_in_data_159}; // @[Cat.scala 30:58]
  assign sram_19_io_r_en = io_pcie_o_r_en & cs_hit_19; // @[outport.scala 32:42]
  assign sram_19_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_20_clock = clock;
  assign sram_20_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_20_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_20_io_w_data = {exe_io_w_data_hi_125,io_phv_in_data_167}; // @[Cat.scala 30:58]
  assign sram_20_io_r_en = io_pcie_o_r_en & cs_hit_20; // @[outport.scala 32:42]
  assign sram_20_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_21_clock = clock;
  assign sram_21_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_21_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_21_io_w_data = {exe_io_w_data_hi_131,io_phv_in_data_175}; // @[Cat.scala 30:58]
  assign sram_21_io_r_en = io_pcie_o_r_en & cs_hit_21; // @[outport.scala 32:42]
  assign sram_21_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_22_clock = clock;
  assign sram_22_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_22_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_22_io_w_data = {exe_io_w_data_hi_137,io_phv_in_data_183}; // @[Cat.scala 30:58]
  assign sram_22_io_r_en = io_pcie_o_r_en & cs_hit_22; // @[outport.scala 32:42]
  assign sram_22_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_23_clock = clock;
  assign sram_23_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_23_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_23_io_w_data = {exe_io_w_data_hi_143,io_phv_in_data_191}; // @[Cat.scala 30:58]
  assign sram_23_io_r_en = io_pcie_o_r_en & cs_hit_23; // @[outport.scala 32:42]
  assign sram_23_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_24_clock = clock;
  assign sram_24_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_24_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_24_io_w_data = {exe_io_w_data_hi_149,io_phv_in_data_199}; // @[Cat.scala 30:58]
  assign sram_24_io_r_en = io_pcie_o_r_en & cs_hit_24; // @[outport.scala 32:42]
  assign sram_24_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_25_clock = clock;
  assign sram_25_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_25_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_25_io_w_data = {exe_io_w_data_hi_155,io_phv_in_data_207}; // @[Cat.scala 30:58]
  assign sram_25_io_r_en = io_pcie_o_r_en & cs_hit_25; // @[outport.scala 32:42]
  assign sram_25_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_26_clock = clock;
  assign sram_26_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_26_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_26_io_w_data = {exe_io_w_data_hi_161,io_phv_in_data_215}; // @[Cat.scala 30:58]
  assign sram_26_io_r_en = io_pcie_o_r_en & cs_hit_26; // @[outport.scala 32:42]
  assign sram_26_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_27_clock = clock;
  assign sram_27_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_27_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_27_io_w_data = {exe_io_w_data_hi_167,io_phv_in_data_223}; // @[Cat.scala 30:58]
  assign sram_27_io_r_en = io_pcie_o_r_en & cs_hit_27; // @[outport.scala 32:42]
  assign sram_27_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_28_clock = clock;
  assign sram_28_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_28_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_28_io_w_data = {exe_io_w_data_hi_173,io_phv_in_data_231}; // @[Cat.scala 30:58]
  assign sram_28_io_r_en = io_pcie_o_r_en & cs_hit_28; // @[outport.scala 32:42]
  assign sram_28_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_29_clock = clock;
  assign sram_29_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_29_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_29_io_w_data = {exe_io_w_data_hi_179,io_phv_in_data_239}; // @[Cat.scala 30:58]
  assign sram_29_io_r_en = io_pcie_o_r_en & cs_hit_29; // @[outport.scala 32:42]
  assign sram_29_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_30_clock = clock;
  assign sram_30_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_30_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_30_io_w_data = {exe_io_w_data_hi_185,io_phv_in_data_247}; // @[Cat.scala 30:58]
  assign sram_30_io_r_en = io_pcie_o_r_en & cs_hit_30; // @[outport.scala 32:42]
  assign sram_30_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_31_clock = clock;
  assign sram_31_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_31_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_31_io_w_data = {exe_io_w_data_hi_191,io_phv_in_data_255}; // @[Cat.scala 30:58]
  assign sram_31_io_r_en = io_pcie_o_r_en & cs_hit_31; // @[outport.scala 32:42]
  assign sram_31_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_32_clock = clock;
  assign sram_32_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_32_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_32_io_w_data = {exe_io_w_data_hi_197,io_phv_in_data_263}; // @[Cat.scala 30:58]
  assign sram_32_io_r_en = io_pcie_o_r_en & cs_hit_32; // @[outport.scala 32:42]
  assign sram_32_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_33_clock = clock;
  assign sram_33_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_33_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_33_io_w_data = {exe_io_w_data_hi_203,io_phv_in_data_271}; // @[Cat.scala 30:58]
  assign sram_33_io_r_en = io_pcie_o_r_en & cs_hit_33; // @[outport.scala 32:42]
  assign sram_33_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_34_clock = clock;
  assign sram_34_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_34_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_34_io_w_data = {exe_io_w_data_hi_209,io_phv_in_data_279}; // @[Cat.scala 30:58]
  assign sram_34_io_r_en = io_pcie_o_r_en & cs_hit_34; // @[outport.scala 32:42]
  assign sram_34_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_35_clock = clock;
  assign sram_35_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_35_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_35_io_w_data = {exe_io_w_data_hi_215,io_phv_in_data_287}; // @[Cat.scala 30:58]
  assign sram_35_io_r_en = io_pcie_o_r_en & cs_hit_35; // @[outport.scala 32:42]
  assign sram_35_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_36_clock = clock;
  assign sram_36_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_36_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_36_io_w_data = {exe_io_w_data_hi_221,io_phv_in_data_295}; // @[Cat.scala 30:58]
  assign sram_36_io_r_en = io_pcie_o_r_en & cs_hit_36; // @[outport.scala 32:42]
  assign sram_36_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_37_clock = clock;
  assign sram_37_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_37_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_37_io_w_data = {exe_io_w_data_hi_227,io_phv_in_data_303}; // @[Cat.scala 30:58]
  assign sram_37_io_r_en = io_pcie_o_r_en & cs_hit_37; // @[outport.scala 32:42]
  assign sram_37_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_38_clock = clock;
  assign sram_38_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_38_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_38_io_w_data = {exe_io_w_data_hi_233,io_phv_in_data_311}; // @[Cat.scala 30:58]
  assign sram_38_io_r_en = io_pcie_o_r_en & cs_hit_38; // @[outport.scala 32:42]
  assign sram_38_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_39_clock = clock;
  assign sram_39_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_39_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_39_io_w_data = {exe_io_w_data_hi_239,io_phv_in_data_319}; // @[Cat.scala 30:58]
  assign sram_39_io_r_en = io_pcie_o_r_en & cs_hit_39; // @[outport.scala 32:42]
  assign sram_39_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_40_clock = clock;
  assign sram_40_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_40_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_40_io_w_data = {exe_io_w_data_hi_245,io_phv_in_data_327}; // @[Cat.scala 30:58]
  assign sram_40_io_r_en = io_pcie_o_r_en & cs_hit_40; // @[outport.scala 32:42]
  assign sram_40_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_41_clock = clock;
  assign sram_41_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_41_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_41_io_w_data = {exe_io_w_data_hi_251,io_phv_in_data_335}; // @[Cat.scala 30:58]
  assign sram_41_io_r_en = io_pcie_o_r_en & cs_hit_41; // @[outport.scala 32:42]
  assign sram_41_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_42_clock = clock;
  assign sram_42_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_42_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_42_io_w_data = {exe_io_w_data_hi_257,io_phv_in_data_343}; // @[Cat.scala 30:58]
  assign sram_42_io_r_en = io_pcie_o_r_en & cs_hit_42; // @[outport.scala 32:42]
  assign sram_42_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_43_clock = clock;
  assign sram_43_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_43_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_43_io_w_data = {exe_io_w_data_hi_263,io_phv_in_data_351}; // @[Cat.scala 30:58]
  assign sram_43_io_r_en = io_pcie_o_r_en & cs_hit_43; // @[outport.scala 32:42]
  assign sram_43_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_44_clock = clock;
  assign sram_44_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_44_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_44_io_w_data = {exe_io_w_data_hi_269,io_phv_in_data_359}; // @[Cat.scala 30:58]
  assign sram_44_io_r_en = io_pcie_o_r_en & cs_hit_44; // @[outport.scala 32:42]
  assign sram_44_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_45_clock = clock;
  assign sram_45_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_45_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_45_io_w_data = {exe_io_w_data_hi_275,io_phv_in_data_367}; // @[Cat.scala 30:58]
  assign sram_45_io_r_en = io_pcie_o_r_en & cs_hit_45; // @[outport.scala 32:42]
  assign sram_45_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_46_clock = clock;
  assign sram_46_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_46_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_46_io_w_data = {exe_io_w_data_hi_281,io_phv_in_data_375}; // @[Cat.scala 30:58]
  assign sram_46_io_r_en = io_pcie_o_r_en & cs_hit_46; // @[outport.scala 32:42]
  assign sram_46_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_47_clock = clock;
  assign sram_47_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_47_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_47_io_w_data = {exe_io_w_data_hi_287,io_phv_in_data_383}; // @[Cat.scala 30:58]
  assign sram_47_io_r_en = io_pcie_o_r_en & cs_hit_47; // @[outport.scala 32:42]
  assign sram_47_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_48_clock = clock;
  assign sram_48_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_48_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_48_io_w_data = {exe_io_w_data_hi_293,io_phv_in_data_391}; // @[Cat.scala 30:58]
  assign sram_48_io_r_en = io_pcie_o_r_en & cs_hit_48; // @[outport.scala 32:42]
  assign sram_48_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_49_clock = clock;
  assign sram_49_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_49_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_49_io_w_data = {exe_io_w_data_hi_299,io_phv_in_data_399}; // @[Cat.scala 30:58]
  assign sram_49_io_r_en = io_pcie_o_r_en & cs_hit_49; // @[outport.scala 32:42]
  assign sram_49_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_50_clock = clock;
  assign sram_50_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_50_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_50_io_w_data = {exe_io_w_data_hi_305,io_phv_in_data_407}; // @[Cat.scala 30:58]
  assign sram_50_io_r_en = io_pcie_o_r_en & cs_hit_50; // @[outport.scala 32:42]
  assign sram_50_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_51_clock = clock;
  assign sram_51_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_51_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_51_io_w_data = {exe_io_w_data_hi_311,io_phv_in_data_415}; // @[Cat.scala 30:58]
  assign sram_51_io_r_en = io_pcie_o_r_en & cs_hit_51; // @[outport.scala 32:42]
  assign sram_51_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_52_clock = clock;
  assign sram_52_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_52_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_52_io_w_data = {exe_io_w_data_hi_317,io_phv_in_data_423}; // @[Cat.scala 30:58]
  assign sram_52_io_r_en = io_pcie_o_r_en & cs_hit_52; // @[outport.scala 32:42]
  assign sram_52_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_53_clock = clock;
  assign sram_53_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_53_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_53_io_w_data = {exe_io_w_data_hi_323,io_phv_in_data_431}; // @[Cat.scala 30:58]
  assign sram_53_io_r_en = io_pcie_o_r_en & cs_hit_53; // @[outport.scala 32:42]
  assign sram_53_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_54_clock = clock;
  assign sram_54_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_54_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_54_io_w_data = {exe_io_w_data_hi_329,io_phv_in_data_439}; // @[Cat.scala 30:58]
  assign sram_54_io_r_en = io_pcie_o_r_en & cs_hit_54; // @[outport.scala 32:42]
  assign sram_54_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_55_clock = clock;
  assign sram_55_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_55_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_55_io_w_data = {exe_io_w_data_hi_335,io_phv_in_data_447}; // @[Cat.scala 30:58]
  assign sram_55_io_r_en = io_pcie_o_r_en & cs_hit_55; // @[outport.scala 32:42]
  assign sram_55_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_56_clock = clock;
  assign sram_56_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_56_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_56_io_w_data = {exe_io_w_data_hi_341,io_phv_in_data_455}; // @[Cat.scala 30:58]
  assign sram_56_io_r_en = io_pcie_o_r_en & cs_hit_56; // @[outport.scala 32:42]
  assign sram_56_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_57_clock = clock;
  assign sram_57_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_57_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_57_io_w_data = {exe_io_w_data_hi_347,io_phv_in_data_463}; // @[Cat.scala 30:58]
  assign sram_57_io_r_en = io_pcie_o_r_en & cs_hit_57; // @[outport.scala 32:42]
  assign sram_57_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_58_clock = clock;
  assign sram_58_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_58_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_58_io_w_data = {exe_io_w_data_hi_353,io_phv_in_data_471}; // @[Cat.scala 30:58]
  assign sram_58_io_r_en = io_pcie_o_r_en & cs_hit_58; // @[outport.scala 32:42]
  assign sram_58_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_59_clock = clock;
  assign sram_59_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_59_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_59_io_w_data = {exe_io_w_data_hi_359,io_phv_in_data_479}; // @[Cat.scala 30:58]
  assign sram_59_io_r_en = io_pcie_o_r_en & cs_hit_59; // @[outport.scala 32:42]
  assign sram_59_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_60_clock = clock;
  assign sram_60_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_60_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_60_io_w_data = {exe_io_w_data_hi_365,io_phv_in_data_487}; // @[Cat.scala 30:58]
  assign sram_60_io_r_en = io_pcie_o_r_en & cs_hit_60; // @[outport.scala 32:42]
  assign sram_60_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_61_clock = clock;
  assign sram_61_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_61_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_61_io_w_data = {exe_io_w_data_hi_371,io_phv_in_data_495}; // @[Cat.scala 30:58]
  assign sram_61_io_r_en = io_pcie_o_r_en & cs_hit_61; // @[outport.scala 32:42]
  assign sram_61_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_62_clock = clock;
  assign sram_62_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_62_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_62_io_w_data = {exe_io_w_data_hi_377,io_phv_in_data_503}; // @[Cat.scala 30:58]
  assign sram_62_io_r_en = io_pcie_o_r_en & cs_hit_62; // @[outport.scala 32:42]
  assign sram_62_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  assign sram_63_clock = clock;
  assign sram_63_io_w_en = 1'h1; // @[outport.scala 24:24]
  assign sram_63_io_w_addr = addr; // @[outport.scala 25:24]
  assign sram_63_io_w_data = {exe_io_w_data_hi_383,io_phv_in_data_511}; // @[Cat.scala 30:58]
  assign sram_63_io_r_en = io_pcie_o_r_en & cs_hit_63; // @[outport.scala 32:42]
  assign sram_63_io_r_addr = io_pcie_o_r_addr; // @[outport.scala 33:24]
  always @(posedge clock) begin
    addr <= addr + 8'h1; // @[outport.scala 18:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
