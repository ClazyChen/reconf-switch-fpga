module HashSumLevel(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [7:0]   io_pipe_phv_in_data_160,
  input  [7:0]   io_pipe_phv_in_data_161,
  input  [7:0]   io_pipe_phv_in_data_162,
  input  [7:0]   io_pipe_phv_in_data_163,
  input  [7:0]   io_pipe_phv_in_data_164,
  input  [7:0]   io_pipe_phv_in_data_165,
  input  [7:0]   io_pipe_phv_in_data_166,
  input  [7:0]   io_pipe_phv_in_data_167,
  input  [7:0]   io_pipe_phv_in_data_168,
  input  [7:0]   io_pipe_phv_in_data_169,
  input  [7:0]   io_pipe_phv_in_data_170,
  input  [7:0]   io_pipe_phv_in_data_171,
  input  [7:0]   io_pipe_phv_in_data_172,
  input  [7:0]   io_pipe_phv_in_data_173,
  input  [7:0]   io_pipe_phv_in_data_174,
  input  [7:0]   io_pipe_phv_in_data_175,
  input  [7:0]   io_pipe_phv_in_data_176,
  input  [7:0]   io_pipe_phv_in_data_177,
  input  [7:0]   io_pipe_phv_in_data_178,
  input  [7:0]   io_pipe_phv_in_data_179,
  input  [7:0]   io_pipe_phv_in_data_180,
  input  [7:0]   io_pipe_phv_in_data_181,
  input  [7:0]   io_pipe_phv_in_data_182,
  input  [7:0]   io_pipe_phv_in_data_183,
  input  [7:0]   io_pipe_phv_in_data_184,
  input  [7:0]   io_pipe_phv_in_data_185,
  input  [7:0]   io_pipe_phv_in_data_186,
  input  [7:0]   io_pipe_phv_in_data_187,
  input  [7:0]   io_pipe_phv_in_data_188,
  input  [7:0]   io_pipe_phv_in_data_189,
  input  [7:0]   io_pipe_phv_in_data_190,
  input  [7:0]   io_pipe_phv_in_data_191,
  input  [7:0]   io_pipe_phv_in_data_192,
  input  [7:0]   io_pipe_phv_in_data_193,
  input  [7:0]   io_pipe_phv_in_data_194,
  input  [7:0]   io_pipe_phv_in_data_195,
  input  [7:0]   io_pipe_phv_in_data_196,
  input  [7:0]   io_pipe_phv_in_data_197,
  input  [7:0]   io_pipe_phv_in_data_198,
  input  [7:0]   io_pipe_phv_in_data_199,
  input  [7:0]   io_pipe_phv_in_data_200,
  input  [7:0]   io_pipe_phv_in_data_201,
  input  [7:0]   io_pipe_phv_in_data_202,
  input  [7:0]   io_pipe_phv_in_data_203,
  input  [7:0]   io_pipe_phv_in_data_204,
  input  [7:0]   io_pipe_phv_in_data_205,
  input  [7:0]   io_pipe_phv_in_data_206,
  input  [7:0]   io_pipe_phv_in_data_207,
  input  [7:0]   io_pipe_phv_in_data_208,
  input  [7:0]   io_pipe_phv_in_data_209,
  input  [7:0]   io_pipe_phv_in_data_210,
  input  [7:0]   io_pipe_phv_in_data_211,
  input  [7:0]   io_pipe_phv_in_data_212,
  input  [7:0]   io_pipe_phv_in_data_213,
  input  [7:0]   io_pipe_phv_in_data_214,
  input  [7:0]   io_pipe_phv_in_data_215,
  input  [7:0]   io_pipe_phv_in_data_216,
  input  [7:0]   io_pipe_phv_in_data_217,
  input  [7:0]   io_pipe_phv_in_data_218,
  input  [7:0]   io_pipe_phv_in_data_219,
  input  [7:0]   io_pipe_phv_in_data_220,
  input  [7:0]   io_pipe_phv_in_data_221,
  input  [7:0]   io_pipe_phv_in_data_222,
  input  [7:0]   io_pipe_phv_in_data_223,
  input  [7:0]   io_pipe_phv_in_data_224,
  input  [7:0]   io_pipe_phv_in_data_225,
  input  [7:0]   io_pipe_phv_in_data_226,
  input  [7:0]   io_pipe_phv_in_data_227,
  input  [7:0]   io_pipe_phv_in_data_228,
  input  [7:0]   io_pipe_phv_in_data_229,
  input  [7:0]   io_pipe_phv_in_data_230,
  input  [7:0]   io_pipe_phv_in_data_231,
  input  [7:0]   io_pipe_phv_in_data_232,
  input  [7:0]   io_pipe_phv_in_data_233,
  input  [7:0]   io_pipe_phv_in_data_234,
  input  [7:0]   io_pipe_phv_in_data_235,
  input  [7:0]   io_pipe_phv_in_data_236,
  input  [7:0]   io_pipe_phv_in_data_237,
  input  [7:0]   io_pipe_phv_in_data_238,
  input  [7:0]   io_pipe_phv_in_data_239,
  input  [7:0]   io_pipe_phv_in_data_240,
  input  [7:0]   io_pipe_phv_in_data_241,
  input  [7:0]   io_pipe_phv_in_data_242,
  input  [7:0]   io_pipe_phv_in_data_243,
  input  [7:0]   io_pipe_phv_in_data_244,
  input  [7:0]   io_pipe_phv_in_data_245,
  input  [7:0]   io_pipe_phv_in_data_246,
  input  [7:0]   io_pipe_phv_in_data_247,
  input  [7:0]   io_pipe_phv_in_data_248,
  input  [7:0]   io_pipe_phv_in_data_249,
  input  [7:0]   io_pipe_phv_in_data_250,
  input  [7:0]   io_pipe_phv_in_data_251,
  input  [7:0]   io_pipe_phv_in_data_252,
  input  [7:0]   io_pipe_phv_in_data_253,
  input  [7:0]   io_pipe_phv_in_data_254,
  input  [7:0]   io_pipe_phv_in_data_255,
  input  [7:0]   io_pipe_phv_in_data_256,
  input  [7:0]   io_pipe_phv_in_data_257,
  input  [7:0]   io_pipe_phv_in_data_258,
  input  [7:0]   io_pipe_phv_in_data_259,
  input  [7:0]   io_pipe_phv_in_data_260,
  input  [7:0]   io_pipe_phv_in_data_261,
  input  [7:0]   io_pipe_phv_in_data_262,
  input  [7:0]   io_pipe_phv_in_data_263,
  input  [7:0]   io_pipe_phv_in_data_264,
  input  [7:0]   io_pipe_phv_in_data_265,
  input  [7:0]   io_pipe_phv_in_data_266,
  input  [7:0]   io_pipe_phv_in_data_267,
  input  [7:0]   io_pipe_phv_in_data_268,
  input  [7:0]   io_pipe_phv_in_data_269,
  input  [7:0]   io_pipe_phv_in_data_270,
  input  [7:0]   io_pipe_phv_in_data_271,
  input  [7:0]   io_pipe_phv_in_data_272,
  input  [7:0]   io_pipe_phv_in_data_273,
  input  [7:0]   io_pipe_phv_in_data_274,
  input  [7:0]   io_pipe_phv_in_data_275,
  input  [7:0]   io_pipe_phv_in_data_276,
  input  [7:0]   io_pipe_phv_in_data_277,
  input  [7:0]   io_pipe_phv_in_data_278,
  input  [7:0]   io_pipe_phv_in_data_279,
  input  [7:0]   io_pipe_phv_in_data_280,
  input  [7:0]   io_pipe_phv_in_data_281,
  input  [7:0]   io_pipe_phv_in_data_282,
  input  [7:0]   io_pipe_phv_in_data_283,
  input  [7:0]   io_pipe_phv_in_data_284,
  input  [7:0]   io_pipe_phv_in_data_285,
  input  [7:0]   io_pipe_phv_in_data_286,
  input  [7:0]   io_pipe_phv_in_data_287,
  input  [7:0]   io_pipe_phv_in_data_288,
  input  [7:0]   io_pipe_phv_in_data_289,
  input  [7:0]   io_pipe_phv_in_data_290,
  input  [7:0]   io_pipe_phv_in_data_291,
  input  [7:0]   io_pipe_phv_in_data_292,
  input  [7:0]   io_pipe_phv_in_data_293,
  input  [7:0]   io_pipe_phv_in_data_294,
  input  [7:0]   io_pipe_phv_in_data_295,
  input  [7:0]   io_pipe_phv_in_data_296,
  input  [7:0]   io_pipe_phv_in_data_297,
  input  [7:0]   io_pipe_phv_in_data_298,
  input  [7:0]   io_pipe_phv_in_data_299,
  input  [7:0]   io_pipe_phv_in_data_300,
  input  [7:0]   io_pipe_phv_in_data_301,
  input  [7:0]   io_pipe_phv_in_data_302,
  input  [7:0]   io_pipe_phv_in_data_303,
  input  [7:0]   io_pipe_phv_in_data_304,
  input  [7:0]   io_pipe_phv_in_data_305,
  input  [7:0]   io_pipe_phv_in_data_306,
  input  [7:0]   io_pipe_phv_in_data_307,
  input  [7:0]   io_pipe_phv_in_data_308,
  input  [7:0]   io_pipe_phv_in_data_309,
  input  [7:0]   io_pipe_phv_in_data_310,
  input  [7:0]   io_pipe_phv_in_data_311,
  input  [7:0]   io_pipe_phv_in_data_312,
  input  [7:0]   io_pipe_phv_in_data_313,
  input  [7:0]   io_pipe_phv_in_data_314,
  input  [7:0]   io_pipe_phv_in_data_315,
  input  [7:0]   io_pipe_phv_in_data_316,
  input  [7:0]   io_pipe_phv_in_data_317,
  input  [7:0]   io_pipe_phv_in_data_318,
  input  [7:0]   io_pipe_phv_in_data_319,
  input  [7:0]   io_pipe_phv_in_data_320,
  input  [7:0]   io_pipe_phv_in_data_321,
  input  [7:0]   io_pipe_phv_in_data_322,
  input  [7:0]   io_pipe_phv_in_data_323,
  input  [7:0]   io_pipe_phv_in_data_324,
  input  [7:0]   io_pipe_phv_in_data_325,
  input  [7:0]   io_pipe_phv_in_data_326,
  input  [7:0]   io_pipe_phv_in_data_327,
  input  [7:0]   io_pipe_phv_in_data_328,
  input  [7:0]   io_pipe_phv_in_data_329,
  input  [7:0]   io_pipe_phv_in_data_330,
  input  [7:0]   io_pipe_phv_in_data_331,
  input  [7:0]   io_pipe_phv_in_data_332,
  input  [7:0]   io_pipe_phv_in_data_333,
  input  [7:0]   io_pipe_phv_in_data_334,
  input  [7:0]   io_pipe_phv_in_data_335,
  input  [7:0]   io_pipe_phv_in_data_336,
  input  [7:0]   io_pipe_phv_in_data_337,
  input  [7:0]   io_pipe_phv_in_data_338,
  input  [7:0]   io_pipe_phv_in_data_339,
  input  [7:0]   io_pipe_phv_in_data_340,
  input  [7:0]   io_pipe_phv_in_data_341,
  input  [7:0]   io_pipe_phv_in_data_342,
  input  [7:0]   io_pipe_phv_in_data_343,
  input  [7:0]   io_pipe_phv_in_data_344,
  input  [7:0]   io_pipe_phv_in_data_345,
  input  [7:0]   io_pipe_phv_in_data_346,
  input  [7:0]   io_pipe_phv_in_data_347,
  input  [7:0]   io_pipe_phv_in_data_348,
  input  [7:0]   io_pipe_phv_in_data_349,
  input  [7:0]   io_pipe_phv_in_data_350,
  input  [7:0]   io_pipe_phv_in_data_351,
  input  [7:0]   io_pipe_phv_in_data_352,
  input  [7:0]   io_pipe_phv_in_data_353,
  input  [7:0]   io_pipe_phv_in_data_354,
  input  [7:0]   io_pipe_phv_in_data_355,
  input  [7:0]   io_pipe_phv_in_data_356,
  input  [7:0]   io_pipe_phv_in_data_357,
  input  [7:0]   io_pipe_phv_in_data_358,
  input  [7:0]   io_pipe_phv_in_data_359,
  input  [7:0]   io_pipe_phv_in_data_360,
  input  [7:0]   io_pipe_phv_in_data_361,
  input  [7:0]   io_pipe_phv_in_data_362,
  input  [7:0]   io_pipe_phv_in_data_363,
  input  [7:0]   io_pipe_phv_in_data_364,
  input  [7:0]   io_pipe_phv_in_data_365,
  input  [7:0]   io_pipe_phv_in_data_366,
  input  [7:0]   io_pipe_phv_in_data_367,
  input  [7:0]   io_pipe_phv_in_data_368,
  input  [7:0]   io_pipe_phv_in_data_369,
  input  [7:0]   io_pipe_phv_in_data_370,
  input  [7:0]   io_pipe_phv_in_data_371,
  input  [7:0]   io_pipe_phv_in_data_372,
  input  [7:0]   io_pipe_phv_in_data_373,
  input  [7:0]   io_pipe_phv_in_data_374,
  input  [7:0]   io_pipe_phv_in_data_375,
  input  [7:0]   io_pipe_phv_in_data_376,
  input  [7:0]   io_pipe_phv_in_data_377,
  input  [7:0]   io_pipe_phv_in_data_378,
  input  [7:0]   io_pipe_phv_in_data_379,
  input  [7:0]   io_pipe_phv_in_data_380,
  input  [7:0]   io_pipe_phv_in_data_381,
  input  [7:0]   io_pipe_phv_in_data_382,
  input  [7:0]   io_pipe_phv_in_data_383,
  input  [7:0]   io_pipe_phv_in_data_384,
  input  [7:0]   io_pipe_phv_in_data_385,
  input  [7:0]   io_pipe_phv_in_data_386,
  input  [7:0]   io_pipe_phv_in_data_387,
  input  [7:0]   io_pipe_phv_in_data_388,
  input  [7:0]   io_pipe_phv_in_data_389,
  input  [7:0]   io_pipe_phv_in_data_390,
  input  [7:0]   io_pipe_phv_in_data_391,
  input  [7:0]   io_pipe_phv_in_data_392,
  input  [7:0]   io_pipe_phv_in_data_393,
  input  [7:0]   io_pipe_phv_in_data_394,
  input  [7:0]   io_pipe_phv_in_data_395,
  input  [7:0]   io_pipe_phv_in_data_396,
  input  [7:0]   io_pipe_phv_in_data_397,
  input  [7:0]   io_pipe_phv_in_data_398,
  input  [7:0]   io_pipe_phv_in_data_399,
  input  [7:0]   io_pipe_phv_in_data_400,
  input  [7:0]   io_pipe_phv_in_data_401,
  input  [7:0]   io_pipe_phv_in_data_402,
  input  [7:0]   io_pipe_phv_in_data_403,
  input  [7:0]   io_pipe_phv_in_data_404,
  input  [7:0]   io_pipe_phv_in_data_405,
  input  [7:0]   io_pipe_phv_in_data_406,
  input  [7:0]   io_pipe_phv_in_data_407,
  input  [7:0]   io_pipe_phv_in_data_408,
  input  [7:0]   io_pipe_phv_in_data_409,
  input  [7:0]   io_pipe_phv_in_data_410,
  input  [7:0]   io_pipe_phv_in_data_411,
  input  [7:0]   io_pipe_phv_in_data_412,
  input  [7:0]   io_pipe_phv_in_data_413,
  input  [7:0]   io_pipe_phv_in_data_414,
  input  [7:0]   io_pipe_phv_in_data_415,
  input  [7:0]   io_pipe_phv_in_data_416,
  input  [7:0]   io_pipe_phv_in_data_417,
  input  [7:0]   io_pipe_phv_in_data_418,
  input  [7:0]   io_pipe_phv_in_data_419,
  input  [7:0]   io_pipe_phv_in_data_420,
  input  [7:0]   io_pipe_phv_in_data_421,
  input  [7:0]   io_pipe_phv_in_data_422,
  input  [7:0]   io_pipe_phv_in_data_423,
  input  [7:0]   io_pipe_phv_in_data_424,
  input  [7:0]   io_pipe_phv_in_data_425,
  input  [7:0]   io_pipe_phv_in_data_426,
  input  [7:0]   io_pipe_phv_in_data_427,
  input  [7:0]   io_pipe_phv_in_data_428,
  input  [7:0]   io_pipe_phv_in_data_429,
  input  [7:0]   io_pipe_phv_in_data_430,
  input  [7:0]   io_pipe_phv_in_data_431,
  input  [7:0]   io_pipe_phv_in_data_432,
  input  [7:0]   io_pipe_phv_in_data_433,
  input  [7:0]   io_pipe_phv_in_data_434,
  input  [7:0]   io_pipe_phv_in_data_435,
  input  [7:0]   io_pipe_phv_in_data_436,
  input  [7:0]   io_pipe_phv_in_data_437,
  input  [7:0]   io_pipe_phv_in_data_438,
  input  [7:0]   io_pipe_phv_in_data_439,
  input  [7:0]   io_pipe_phv_in_data_440,
  input  [7:0]   io_pipe_phv_in_data_441,
  input  [7:0]   io_pipe_phv_in_data_442,
  input  [7:0]   io_pipe_phv_in_data_443,
  input  [7:0]   io_pipe_phv_in_data_444,
  input  [7:0]   io_pipe_phv_in_data_445,
  input  [7:0]   io_pipe_phv_in_data_446,
  input  [7:0]   io_pipe_phv_in_data_447,
  input  [7:0]   io_pipe_phv_in_data_448,
  input  [7:0]   io_pipe_phv_in_data_449,
  input  [7:0]   io_pipe_phv_in_data_450,
  input  [7:0]   io_pipe_phv_in_data_451,
  input  [7:0]   io_pipe_phv_in_data_452,
  input  [7:0]   io_pipe_phv_in_data_453,
  input  [7:0]   io_pipe_phv_in_data_454,
  input  [7:0]   io_pipe_phv_in_data_455,
  input  [7:0]   io_pipe_phv_in_data_456,
  input  [7:0]   io_pipe_phv_in_data_457,
  input  [7:0]   io_pipe_phv_in_data_458,
  input  [7:0]   io_pipe_phv_in_data_459,
  input  [7:0]   io_pipe_phv_in_data_460,
  input  [7:0]   io_pipe_phv_in_data_461,
  input  [7:0]   io_pipe_phv_in_data_462,
  input  [7:0]   io_pipe_phv_in_data_463,
  input  [7:0]   io_pipe_phv_in_data_464,
  input  [7:0]   io_pipe_phv_in_data_465,
  input  [7:0]   io_pipe_phv_in_data_466,
  input  [7:0]   io_pipe_phv_in_data_467,
  input  [7:0]   io_pipe_phv_in_data_468,
  input  [7:0]   io_pipe_phv_in_data_469,
  input  [7:0]   io_pipe_phv_in_data_470,
  input  [7:0]   io_pipe_phv_in_data_471,
  input  [7:0]   io_pipe_phv_in_data_472,
  input  [7:0]   io_pipe_phv_in_data_473,
  input  [7:0]   io_pipe_phv_in_data_474,
  input  [7:0]   io_pipe_phv_in_data_475,
  input  [7:0]   io_pipe_phv_in_data_476,
  input  [7:0]   io_pipe_phv_in_data_477,
  input  [7:0]   io_pipe_phv_in_data_478,
  input  [7:0]   io_pipe_phv_in_data_479,
  input  [7:0]   io_pipe_phv_in_data_480,
  input  [7:0]   io_pipe_phv_in_data_481,
  input  [7:0]   io_pipe_phv_in_data_482,
  input  [7:0]   io_pipe_phv_in_data_483,
  input  [7:0]   io_pipe_phv_in_data_484,
  input  [7:0]   io_pipe_phv_in_data_485,
  input  [7:0]   io_pipe_phv_in_data_486,
  input  [7:0]   io_pipe_phv_in_data_487,
  input  [7:0]   io_pipe_phv_in_data_488,
  input  [7:0]   io_pipe_phv_in_data_489,
  input  [7:0]   io_pipe_phv_in_data_490,
  input  [7:0]   io_pipe_phv_in_data_491,
  input  [7:0]   io_pipe_phv_in_data_492,
  input  [7:0]   io_pipe_phv_in_data_493,
  input  [7:0]   io_pipe_phv_in_data_494,
  input  [7:0]   io_pipe_phv_in_data_495,
  input  [7:0]   io_pipe_phv_in_data_496,
  input  [7:0]   io_pipe_phv_in_data_497,
  input  [7:0]   io_pipe_phv_in_data_498,
  input  [7:0]   io_pipe_phv_in_data_499,
  input  [7:0]   io_pipe_phv_in_data_500,
  input  [7:0]   io_pipe_phv_in_data_501,
  input  [7:0]   io_pipe_phv_in_data_502,
  input  [7:0]   io_pipe_phv_in_data_503,
  input  [7:0]   io_pipe_phv_in_data_504,
  input  [7:0]   io_pipe_phv_in_data_505,
  input  [7:0]   io_pipe_phv_in_data_506,
  input  [7:0]   io_pipe_phv_in_data_507,
  input  [7:0]   io_pipe_phv_in_data_508,
  input  [7:0]   io_pipe_phv_in_data_509,
  input  [7:0]   io_pipe_phv_in_data_510,
  input  [7:0]   io_pipe_phv_in_data_511,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [7:0]   io_pipe_phv_out_data_160,
  output [7:0]   io_pipe_phv_out_data_161,
  output [7:0]   io_pipe_phv_out_data_162,
  output [7:0]   io_pipe_phv_out_data_163,
  output [7:0]   io_pipe_phv_out_data_164,
  output [7:0]   io_pipe_phv_out_data_165,
  output [7:0]   io_pipe_phv_out_data_166,
  output [7:0]   io_pipe_phv_out_data_167,
  output [7:0]   io_pipe_phv_out_data_168,
  output [7:0]   io_pipe_phv_out_data_169,
  output [7:0]   io_pipe_phv_out_data_170,
  output [7:0]   io_pipe_phv_out_data_171,
  output [7:0]   io_pipe_phv_out_data_172,
  output [7:0]   io_pipe_phv_out_data_173,
  output [7:0]   io_pipe_phv_out_data_174,
  output [7:0]   io_pipe_phv_out_data_175,
  output [7:0]   io_pipe_phv_out_data_176,
  output [7:0]   io_pipe_phv_out_data_177,
  output [7:0]   io_pipe_phv_out_data_178,
  output [7:0]   io_pipe_phv_out_data_179,
  output [7:0]   io_pipe_phv_out_data_180,
  output [7:0]   io_pipe_phv_out_data_181,
  output [7:0]   io_pipe_phv_out_data_182,
  output [7:0]   io_pipe_phv_out_data_183,
  output [7:0]   io_pipe_phv_out_data_184,
  output [7:0]   io_pipe_phv_out_data_185,
  output [7:0]   io_pipe_phv_out_data_186,
  output [7:0]   io_pipe_phv_out_data_187,
  output [7:0]   io_pipe_phv_out_data_188,
  output [7:0]   io_pipe_phv_out_data_189,
  output [7:0]   io_pipe_phv_out_data_190,
  output [7:0]   io_pipe_phv_out_data_191,
  output [7:0]   io_pipe_phv_out_data_192,
  output [7:0]   io_pipe_phv_out_data_193,
  output [7:0]   io_pipe_phv_out_data_194,
  output [7:0]   io_pipe_phv_out_data_195,
  output [7:0]   io_pipe_phv_out_data_196,
  output [7:0]   io_pipe_phv_out_data_197,
  output [7:0]   io_pipe_phv_out_data_198,
  output [7:0]   io_pipe_phv_out_data_199,
  output [7:0]   io_pipe_phv_out_data_200,
  output [7:0]   io_pipe_phv_out_data_201,
  output [7:0]   io_pipe_phv_out_data_202,
  output [7:0]   io_pipe_phv_out_data_203,
  output [7:0]   io_pipe_phv_out_data_204,
  output [7:0]   io_pipe_phv_out_data_205,
  output [7:0]   io_pipe_phv_out_data_206,
  output [7:0]   io_pipe_phv_out_data_207,
  output [7:0]   io_pipe_phv_out_data_208,
  output [7:0]   io_pipe_phv_out_data_209,
  output [7:0]   io_pipe_phv_out_data_210,
  output [7:0]   io_pipe_phv_out_data_211,
  output [7:0]   io_pipe_phv_out_data_212,
  output [7:0]   io_pipe_phv_out_data_213,
  output [7:0]   io_pipe_phv_out_data_214,
  output [7:0]   io_pipe_phv_out_data_215,
  output [7:0]   io_pipe_phv_out_data_216,
  output [7:0]   io_pipe_phv_out_data_217,
  output [7:0]   io_pipe_phv_out_data_218,
  output [7:0]   io_pipe_phv_out_data_219,
  output [7:0]   io_pipe_phv_out_data_220,
  output [7:0]   io_pipe_phv_out_data_221,
  output [7:0]   io_pipe_phv_out_data_222,
  output [7:0]   io_pipe_phv_out_data_223,
  output [7:0]   io_pipe_phv_out_data_224,
  output [7:0]   io_pipe_phv_out_data_225,
  output [7:0]   io_pipe_phv_out_data_226,
  output [7:0]   io_pipe_phv_out_data_227,
  output [7:0]   io_pipe_phv_out_data_228,
  output [7:0]   io_pipe_phv_out_data_229,
  output [7:0]   io_pipe_phv_out_data_230,
  output [7:0]   io_pipe_phv_out_data_231,
  output [7:0]   io_pipe_phv_out_data_232,
  output [7:0]   io_pipe_phv_out_data_233,
  output [7:0]   io_pipe_phv_out_data_234,
  output [7:0]   io_pipe_phv_out_data_235,
  output [7:0]   io_pipe_phv_out_data_236,
  output [7:0]   io_pipe_phv_out_data_237,
  output [7:0]   io_pipe_phv_out_data_238,
  output [7:0]   io_pipe_phv_out_data_239,
  output [7:0]   io_pipe_phv_out_data_240,
  output [7:0]   io_pipe_phv_out_data_241,
  output [7:0]   io_pipe_phv_out_data_242,
  output [7:0]   io_pipe_phv_out_data_243,
  output [7:0]   io_pipe_phv_out_data_244,
  output [7:0]   io_pipe_phv_out_data_245,
  output [7:0]   io_pipe_phv_out_data_246,
  output [7:0]   io_pipe_phv_out_data_247,
  output [7:0]   io_pipe_phv_out_data_248,
  output [7:0]   io_pipe_phv_out_data_249,
  output [7:0]   io_pipe_phv_out_data_250,
  output [7:0]   io_pipe_phv_out_data_251,
  output [7:0]   io_pipe_phv_out_data_252,
  output [7:0]   io_pipe_phv_out_data_253,
  output [7:0]   io_pipe_phv_out_data_254,
  output [7:0]   io_pipe_phv_out_data_255,
  output [7:0]   io_pipe_phv_out_data_256,
  output [7:0]   io_pipe_phv_out_data_257,
  output [7:0]   io_pipe_phv_out_data_258,
  output [7:0]   io_pipe_phv_out_data_259,
  output [7:0]   io_pipe_phv_out_data_260,
  output [7:0]   io_pipe_phv_out_data_261,
  output [7:0]   io_pipe_phv_out_data_262,
  output [7:0]   io_pipe_phv_out_data_263,
  output [7:0]   io_pipe_phv_out_data_264,
  output [7:0]   io_pipe_phv_out_data_265,
  output [7:0]   io_pipe_phv_out_data_266,
  output [7:0]   io_pipe_phv_out_data_267,
  output [7:0]   io_pipe_phv_out_data_268,
  output [7:0]   io_pipe_phv_out_data_269,
  output [7:0]   io_pipe_phv_out_data_270,
  output [7:0]   io_pipe_phv_out_data_271,
  output [7:0]   io_pipe_phv_out_data_272,
  output [7:0]   io_pipe_phv_out_data_273,
  output [7:0]   io_pipe_phv_out_data_274,
  output [7:0]   io_pipe_phv_out_data_275,
  output [7:0]   io_pipe_phv_out_data_276,
  output [7:0]   io_pipe_phv_out_data_277,
  output [7:0]   io_pipe_phv_out_data_278,
  output [7:0]   io_pipe_phv_out_data_279,
  output [7:0]   io_pipe_phv_out_data_280,
  output [7:0]   io_pipe_phv_out_data_281,
  output [7:0]   io_pipe_phv_out_data_282,
  output [7:0]   io_pipe_phv_out_data_283,
  output [7:0]   io_pipe_phv_out_data_284,
  output [7:0]   io_pipe_phv_out_data_285,
  output [7:0]   io_pipe_phv_out_data_286,
  output [7:0]   io_pipe_phv_out_data_287,
  output [7:0]   io_pipe_phv_out_data_288,
  output [7:0]   io_pipe_phv_out_data_289,
  output [7:0]   io_pipe_phv_out_data_290,
  output [7:0]   io_pipe_phv_out_data_291,
  output [7:0]   io_pipe_phv_out_data_292,
  output [7:0]   io_pipe_phv_out_data_293,
  output [7:0]   io_pipe_phv_out_data_294,
  output [7:0]   io_pipe_phv_out_data_295,
  output [7:0]   io_pipe_phv_out_data_296,
  output [7:0]   io_pipe_phv_out_data_297,
  output [7:0]   io_pipe_phv_out_data_298,
  output [7:0]   io_pipe_phv_out_data_299,
  output [7:0]   io_pipe_phv_out_data_300,
  output [7:0]   io_pipe_phv_out_data_301,
  output [7:0]   io_pipe_phv_out_data_302,
  output [7:0]   io_pipe_phv_out_data_303,
  output [7:0]   io_pipe_phv_out_data_304,
  output [7:0]   io_pipe_phv_out_data_305,
  output [7:0]   io_pipe_phv_out_data_306,
  output [7:0]   io_pipe_phv_out_data_307,
  output [7:0]   io_pipe_phv_out_data_308,
  output [7:0]   io_pipe_phv_out_data_309,
  output [7:0]   io_pipe_phv_out_data_310,
  output [7:0]   io_pipe_phv_out_data_311,
  output [7:0]   io_pipe_phv_out_data_312,
  output [7:0]   io_pipe_phv_out_data_313,
  output [7:0]   io_pipe_phv_out_data_314,
  output [7:0]   io_pipe_phv_out_data_315,
  output [7:0]   io_pipe_phv_out_data_316,
  output [7:0]   io_pipe_phv_out_data_317,
  output [7:0]   io_pipe_phv_out_data_318,
  output [7:0]   io_pipe_phv_out_data_319,
  output [7:0]   io_pipe_phv_out_data_320,
  output [7:0]   io_pipe_phv_out_data_321,
  output [7:0]   io_pipe_phv_out_data_322,
  output [7:0]   io_pipe_phv_out_data_323,
  output [7:0]   io_pipe_phv_out_data_324,
  output [7:0]   io_pipe_phv_out_data_325,
  output [7:0]   io_pipe_phv_out_data_326,
  output [7:0]   io_pipe_phv_out_data_327,
  output [7:0]   io_pipe_phv_out_data_328,
  output [7:0]   io_pipe_phv_out_data_329,
  output [7:0]   io_pipe_phv_out_data_330,
  output [7:0]   io_pipe_phv_out_data_331,
  output [7:0]   io_pipe_phv_out_data_332,
  output [7:0]   io_pipe_phv_out_data_333,
  output [7:0]   io_pipe_phv_out_data_334,
  output [7:0]   io_pipe_phv_out_data_335,
  output [7:0]   io_pipe_phv_out_data_336,
  output [7:0]   io_pipe_phv_out_data_337,
  output [7:0]   io_pipe_phv_out_data_338,
  output [7:0]   io_pipe_phv_out_data_339,
  output [7:0]   io_pipe_phv_out_data_340,
  output [7:0]   io_pipe_phv_out_data_341,
  output [7:0]   io_pipe_phv_out_data_342,
  output [7:0]   io_pipe_phv_out_data_343,
  output [7:0]   io_pipe_phv_out_data_344,
  output [7:0]   io_pipe_phv_out_data_345,
  output [7:0]   io_pipe_phv_out_data_346,
  output [7:0]   io_pipe_phv_out_data_347,
  output [7:0]   io_pipe_phv_out_data_348,
  output [7:0]   io_pipe_phv_out_data_349,
  output [7:0]   io_pipe_phv_out_data_350,
  output [7:0]   io_pipe_phv_out_data_351,
  output [7:0]   io_pipe_phv_out_data_352,
  output [7:0]   io_pipe_phv_out_data_353,
  output [7:0]   io_pipe_phv_out_data_354,
  output [7:0]   io_pipe_phv_out_data_355,
  output [7:0]   io_pipe_phv_out_data_356,
  output [7:0]   io_pipe_phv_out_data_357,
  output [7:0]   io_pipe_phv_out_data_358,
  output [7:0]   io_pipe_phv_out_data_359,
  output [7:0]   io_pipe_phv_out_data_360,
  output [7:0]   io_pipe_phv_out_data_361,
  output [7:0]   io_pipe_phv_out_data_362,
  output [7:0]   io_pipe_phv_out_data_363,
  output [7:0]   io_pipe_phv_out_data_364,
  output [7:0]   io_pipe_phv_out_data_365,
  output [7:0]   io_pipe_phv_out_data_366,
  output [7:0]   io_pipe_phv_out_data_367,
  output [7:0]   io_pipe_phv_out_data_368,
  output [7:0]   io_pipe_phv_out_data_369,
  output [7:0]   io_pipe_phv_out_data_370,
  output [7:0]   io_pipe_phv_out_data_371,
  output [7:0]   io_pipe_phv_out_data_372,
  output [7:0]   io_pipe_phv_out_data_373,
  output [7:0]   io_pipe_phv_out_data_374,
  output [7:0]   io_pipe_phv_out_data_375,
  output [7:0]   io_pipe_phv_out_data_376,
  output [7:0]   io_pipe_phv_out_data_377,
  output [7:0]   io_pipe_phv_out_data_378,
  output [7:0]   io_pipe_phv_out_data_379,
  output [7:0]   io_pipe_phv_out_data_380,
  output [7:0]   io_pipe_phv_out_data_381,
  output [7:0]   io_pipe_phv_out_data_382,
  output [7:0]   io_pipe_phv_out_data_383,
  output [7:0]   io_pipe_phv_out_data_384,
  output [7:0]   io_pipe_phv_out_data_385,
  output [7:0]   io_pipe_phv_out_data_386,
  output [7:0]   io_pipe_phv_out_data_387,
  output [7:0]   io_pipe_phv_out_data_388,
  output [7:0]   io_pipe_phv_out_data_389,
  output [7:0]   io_pipe_phv_out_data_390,
  output [7:0]   io_pipe_phv_out_data_391,
  output [7:0]   io_pipe_phv_out_data_392,
  output [7:0]   io_pipe_phv_out_data_393,
  output [7:0]   io_pipe_phv_out_data_394,
  output [7:0]   io_pipe_phv_out_data_395,
  output [7:0]   io_pipe_phv_out_data_396,
  output [7:0]   io_pipe_phv_out_data_397,
  output [7:0]   io_pipe_phv_out_data_398,
  output [7:0]   io_pipe_phv_out_data_399,
  output [7:0]   io_pipe_phv_out_data_400,
  output [7:0]   io_pipe_phv_out_data_401,
  output [7:0]   io_pipe_phv_out_data_402,
  output [7:0]   io_pipe_phv_out_data_403,
  output [7:0]   io_pipe_phv_out_data_404,
  output [7:0]   io_pipe_phv_out_data_405,
  output [7:0]   io_pipe_phv_out_data_406,
  output [7:0]   io_pipe_phv_out_data_407,
  output [7:0]   io_pipe_phv_out_data_408,
  output [7:0]   io_pipe_phv_out_data_409,
  output [7:0]   io_pipe_phv_out_data_410,
  output [7:0]   io_pipe_phv_out_data_411,
  output [7:0]   io_pipe_phv_out_data_412,
  output [7:0]   io_pipe_phv_out_data_413,
  output [7:0]   io_pipe_phv_out_data_414,
  output [7:0]   io_pipe_phv_out_data_415,
  output [7:0]   io_pipe_phv_out_data_416,
  output [7:0]   io_pipe_phv_out_data_417,
  output [7:0]   io_pipe_phv_out_data_418,
  output [7:0]   io_pipe_phv_out_data_419,
  output [7:0]   io_pipe_phv_out_data_420,
  output [7:0]   io_pipe_phv_out_data_421,
  output [7:0]   io_pipe_phv_out_data_422,
  output [7:0]   io_pipe_phv_out_data_423,
  output [7:0]   io_pipe_phv_out_data_424,
  output [7:0]   io_pipe_phv_out_data_425,
  output [7:0]   io_pipe_phv_out_data_426,
  output [7:0]   io_pipe_phv_out_data_427,
  output [7:0]   io_pipe_phv_out_data_428,
  output [7:0]   io_pipe_phv_out_data_429,
  output [7:0]   io_pipe_phv_out_data_430,
  output [7:0]   io_pipe_phv_out_data_431,
  output [7:0]   io_pipe_phv_out_data_432,
  output [7:0]   io_pipe_phv_out_data_433,
  output [7:0]   io_pipe_phv_out_data_434,
  output [7:0]   io_pipe_phv_out_data_435,
  output [7:0]   io_pipe_phv_out_data_436,
  output [7:0]   io_pipe_phv_out_data_437,
  output [7:0]   io_pipe_phv_out_data_438,
  output [7:0]   io_pipe_phv_out_data_439,
  output [7:0]   io_pipe_phv_out_data_440,
  output [7:0]   io_pipe_phv_out_data_441,
  output [7:0]   io_pipe_phv_out_data_442,
  output [7:0]   io_pipe_phv_out_data_443,
  output [7:0]   io_pipe_phv_out_data_444,
  output [7:0]   io_pipe_phv_out_data_445,
  output [7:0]   io_pipe_phv_out_data_446,
  output [7:0]   io_pipe_phv_out_data_447,
  output [7:0]   io_pipe_phv_out_data_448,
  output [7:0]   io_pipe_phv_out_data_449,
  output [7:0]   io_pipe_phv_out_data_450,
  output [7:0]   io_pipe_phv_out_data_451,
  output [7:0]   io_pipe_phv_out_data_452,
  output [7:0]   io_pipe_phv_out_data_453,
  output [7:0]   io_pipe_phv_out_data_454,
  output [7:0]   io_pipe_phv_out_data_455,
  output [7:0]   io_pipe_phv_out_data_456,
  output [7:0]   io_pipe_phv_out_data_457,
  output [7:0]   io_pipe_phv_out_data_458,
  output [7:0]   io_pipe_phv_out_data_459,
  output [7:0]   io_pipe_phv_out_data_460,
  output [7:0]   io_pipe_phv_out_data_461,
  output [7:0]   io_pipe_phv_out_data_462,
  output [7:0]   io_pipe_phv_out_data_463,
  output [7:0]   io_pipe_phv_out_data_464,
  output [7:0]   io_pipe_phv_out_data_465,
  output [7:0]   io_pipe_phv_out_data_466,
  output [7:0]   io_pipe_phv_out_data_467,
  output [7:0]   io_pipe_phv_out_data_468,
  output [7:0]   io_pipe_phv_out_data_469,
  output [7:0]   io_pipe_phv_out_data_470,
  output [7:0]   io_pipe_phv_out_data_471,
  output [7:0]   io_pipe_phv_out_data_472,
  output [7:0]   io_pipe_phv_out_data_473,
  output [7:0]   io_pipe_phv_out_data_474,
  output [7:0]   io_pipe_phv_out_data_475,
  output [7:0]   io_pipe_phv_out_data_476,
  output [7:0]   io_pipe_phv_out_data_477,
  output [7:0]   io_pipe_phv_out_data_478,
  output [7:0]   io_pipe_phv_out_data_479,
  output [7:0]   io_pipe_phv_out_data_480,
  output [7:0]   io_pipe_phv_out_data_481,
  output [7:0]   io_pipe_phv_out_data_482,
  output [7:0]   io_pipe_phv_out_data_483,
  output [7:0]   io_pipe_phv_out_data_484,
  output [7:0]   io_pipe_phv_out_data_485,
  output [7:0]   io_pipe_phv_out_data_486,
  output [7:0]   io_pipe_phv_out_data_487,
  output [7:0]   io_pipe_phv_out_data_488,
  output [7:0]   io_pipe_phv_out_data_489,
  output [7:0]   io_pipe_phv_out_data_490,
  output [7:0]   io_pipe_phv_out_data_491,
  output [7:0]   io_pipe_phv_out_data_492,
  output [7:0]   io_pipe_phv_out_data_493,
  output [7:0]   io_pipe_phv_out_data_494,
  output [7:0]   io_pipe_phv_out_data_495,
  output [7:0]   io_pipe_phv_out_data_496,
  output [7:0]   io_pipe_phv_out_data_497,
  output [7:0]   io_pipe_phv_out_data_498,
  output [7:0]   io_pipe_phv_out_data_499,
  output [7:0]   io_pipe_phv_out_data_500,
  output [7:0]   io_pipe_phv_out_data_501,
  output [7:0]   io_pipe_phv_out_data_502,
  output [7:0]   io_pipe_phv_out_data_503,
  output [7:0]   io_pipe_phv_out_data_504,
  output [7:0]   io_pipe_phv_out_data_505,
  output [7:0]   io_pipe_phv_out_data_506,
  output [7:0]   io_pipe_phv_out_data_507,
  output [7:0]   io_pipe_phv_out_data_508,
  output [7:0]   io_pipe_phv_out_data_509,
  output [7:0]   io_pipe_phv_out_data_510,
  output [7:0]   io_pipe_phv_out_data_511,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [191:0] io_sum_in,
  output [191:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [191:0] _RAND_534;
  reg [191:0] _RAND_535;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 41:22]
  reg [7:0] phv_data_1; // @[hash.scala 41:22]
  reg [7:0] phv_data_2; // @[hash.scala 41:22]
  reg [7:0] phv_data_3; // @[hash.scala 41:22]
  reg [7:0] phv_data_4; // @[hash.scala 41:22]
  reg [7:0] phv_data_5; // @[hash.scala 41:22]
  reg [7:0] phv_data_6; // @[hash.scala 41:22]
  reg [7:0] phv_data_7; // @[hash.scala 41:22]
  reg [7:0] phv_data_8; // @[hash.scala 41:22]
  reg [7:0] phv_data_9; // @[hash.scala 41:22]
  reg [7:0] phv_data_10; // @[hash.scala 41:22]
  reg [7:0] phv_data_11; // @[hash.scala 41:22]
  reg [7:0] phv_data_12; // @[hash.scala 41:22]
  reg [7:0] phv_data_13; // @[hash.scala 41:22]
  reg [7:0] phv_data_14; // @[hash.scala 41:22]
  reg [7:0] phv_data_15; // @[hash.scala 41:22]
  reg [7:0] phv_data_16; // @[hash.scala 41:22]
  reg [7:0] phv_data_17; // @[hash.scala 41:22]
  reg [7:0] phv_data_18; // @[hash.scala 41:22]
  reg [7:0] phv_data_19; // @[hash.scala 41:22]
  reg [7:0] phv_data_20; // @[hash.scala 41:22]
  reg [7:0] phv_data_21; // @[hash.scala 41:22]
  reg [7:0] phv_data_22; // @[hash.scala 41:22]
  reg [7:0] phv_data_23; // @[hash.scala 41:22]
  reg [7:0] phv_data_24; // @[hash.scala 41:22]
  reg [7:0] phv_data_25; // @[hash.scala 41:22]
  reg [7:0] phv_data_26; // @[hash.scala 41:22]
  reg [7:0] phv_data_27; // @[hash.scala 41:22]
  reg [7:0] phv_data_28; // @[hash.scala 41:22]
  reg [7:0] phv_data_29; // @[hash.scala 41:22]
  reg [7:0] phv_data_30; // @[hash.scala 41:22]
  reg [7:0] phv_data_31; // @[hash.scala 41:22]
  reg [7:0] phv_data_32; // @[hash.scala 41:22]
  reg [7:0] phv_data_33; // @[hash.scala 41:22]
  reg [7:0] phv_data_34; // @[hash.scala 41:22]
  reg [7:0] phv_data_35; // @[hash.scala 41:22]
  reg [7:0] phv_data_36; // @[hash.scala 41:22]
  reg [7:0] phv_data_37; // @[hash.scala 41:22]
  reg [7:0] phv_data_38; // @[hash.scala 41:22]
  reg [7:0] phv_data_39; // @[hash.scala 41:22]
  reg [7:0] phv_data_40; // @[hash.scala 41:22]
  reg [7:0] phv_data_41; // @[hash.scala 41:22]
  reg [7:0] phv_data_42; // @[hash.scala 41:22]
  reg [7:0] phv_data_43; // @[hash.scala 41:22]
  reg [7:0] phv_data_44; // @[hash.scala 41:22]
  reg [7:0] phv_data_45; // @[hash.scala 41:22]
  reg [7:0] phv_data_46; // @[hash.scala 41:22]
  reg [7:0] phv_data_47; // @[hash.scala 41:22]
  reg [7:0] phv_data_48; // @[hash.scala 41:22]
  reg [7:0] phv_data_49; // @[hash.scala 41:22]
  reg [7:0] phv_data_50; // @[hash.scala 41:22]
  reg [7:0] phv_data_51; // @[hash.scala 41:22]
  reg [7:0] phv_data_52; // @[hash.scala 41:22]
  reg [7:0] phv_data_53; // @[hash.scala 41:22]
  reg [7:0] phv_data_54; // @[hash.scala 41:22]
  reg [7:0] phv_data_55; // @[hash.scala 41:22]
  reg [7:0] phv_data_56; // @[hash.scala 41:22]
  reg [7:0] phv_data_57; // @[hash.scala 41:22]
  reg [7:0] phv_data_58; // @[hash.scala 41:22]
  reg [7:0] phv_data_59; // @[hash.scala 41:22]
  reg [7:0] phv_data_60; // @[hash.scala 41:22]
  reg [7:0] phv_data_61; // @[hash.scala 41:22]
  reg [7:0] phv_data_62; // @[hash.scala 41:22]
  reg [7:0] phv_data_63; // @[hash.scala 41:22]
  reg [7:0] phv_data_64; // @[hash.scala 41:22]
  reg [7:0] phv_data_65; // @[hash.scala 41:22]
  reg [7:0] phv_data_66; // @[hash.scala 41:22]
  reg [7:0] phv_data_67; // @[hash.scala 41:22]
  reg [7:0] phv_data_68; // @[hash.scala 41:22]
  reg [7:0] phv_data_69; // @[hash.scala 41:22]
  reg [7:0] phv_data_70; // @[hash.scala 41:22]
  reg [7:0] phv_data_71; // @[hash.scala 41:22]
  reg [7:0] phv_data_72; // @[hash.scala 41:22]
  reg [7:0] phv_data_73; // @[hash.scala 41:22]
  reg [7:0] phv_data_74; // @[hash.scala 41:22]
  reg [7:0] phv_data_75; // @[hash.scala 41:22]
  reg [7:0] phv_data_76; // @[hash.scala 41:22]
  reg [7:0] phv_data_77; // @[hash.scala 41:22]
  reg [7:0] phv_data_78; // @[hash.scala 41:22]
  reg [7:0] phv_data_79; // @[hash.scala 41:22]
  reg [7:0] phv_data_80; // @[hash.scala 41:22]
  reg [7:0] phv_data_81; // @[hash.scala 41:22]
  reg [7:0] phv_data_82; // @[hash.scala 41:22]
  reg [7:0] phv_data_83; // @[hash.scala 41:22]
  reg [7:0] phv_data_84; // @[hash.scala 41:22]
  reg [7:0] phv_data_85; // @[hash.scala 41:22]
  reg [7:0] phv_data_86; // @[hash.scala 41:22]
  reg [7:0] phv_data_87; // @[hash.scala 41:22]
  reg [7:0] phv_data_88; // @[hash.scala 41:22]
  reg [7:0] phv_data_89; // @[hash.scala 41:22]
  reg [7:0] phv_data_90; // @[hash.scala 41:22]
  reg [7:0] phv_data_91; // @[hash.scala 41:22]
  reg [7:0] phv_data_92; // @[hash.scala 41:22]
  reg [7:0] phv_data_93; // @[hash.scala 41:22]
  reg [7:0] phv_data_94; // @[hash.scala 41:22]
  reg [7:0] phv_data_95; // @[hash.scala 41:22]
  reg [7:0] phv_data_96; // @[hash.scala 41:22]
  reg [7:0] phv_data_97; // @[hash.scala 41:22]
  reg [7:0] phv_data_98; // @[hash.scala 41:22]
  reg [7:0] phv_data_99; // @[hash.scala 41:22]
  reg [7:0] phv_data_100; // @[hash.scala 41:22]
  reg [7:0] phv_data_101; // @[hash.scala 41:22]
  reg [7:0] phv_data_102; // @[hash.scala 41:22]
  reg [7:0] phv_data_103; // @[hash.scala 41:22]
  reg [7:0] phv_data_104; // @[hash.scala 41:22]
  reg [7:0] phv_data_105; // @[hash.scala 41:22]
  reg [7:0] phv_data_106; // @[hash.scala 41:22]
  reg [7:0] phv_data_107; // @[hash.scala 41:22]
  reg [7:0] phv_data_108; // @[hash.scala 41:22]
  reg [7:0] phv_data_109; // @[hash.scala 41:22]
  reg [7:0] phv_data_110; // @[hash.scala 41:22]
  reg [7:0] phv_data_111; // @[hash.scala 41:22]
  reg [7:0] phv_data_112; // @[hash.scala 41:22]
  reg [7:0] phv_data_113; // @[hash.scala 41:22]
  reg [7:0] phv_data_114; // @[hash.scala 41:22]
  reg [7:0] phv_data_115; // @[hash.scala 41:22]
  reg [7:0] phv_data_116; // @[hash.scala 41:22]
  reg [7:0] phv_data_117; // @[hash.scala 41:22]
  reg [7:0] phv_data_118; // @[hash.scala 41:22]
  reg [7:0] phv_data_119; // @[hash.scala 41:22]
  reg [7:0] phv_data_120; // @[hash.scala 41:22]
  reg [7:0] phv_data_121; // @[hash.scala 41:22]
  reg [7:0] phv_data_122; // @[hash.scala 41:22]
  reg [7:0] phv_data_123; // @[hash.scala 41:22]
  reg [7:0] phv_data_124; // @[hash.scala 41:22]
  reg [7:0] phv_data_125; // @[hash.scala 41:22]
  reg [7:0] phv_data_126; // @[hash.scala 41:22]
  reg [7:0] phv_data_127; // @[hash.scala 41:22]
  reg [7:0] phv_data_128; // @[hash.scala 41:22]
  reg [7:0] phv_data_129; // @[hash.scala 41:22]
  reg [7:0] phv_data_130; // @[hash.scala 41:22]
  reg [7:0] phv_data_131; // @[hash.scala 41:22]
  reg [7:0] phv_data_132; // @[hash.scala 41:22]
  reg [7:0] phv_data_133; // @[hash.scala 41:22]
  reg [7:0] phv_data_134; // @[hash.scala 41:22]
  reg [7:0] phv_data_135; // @[hash.scala 41:22]
  reg [7:0] phv_data_136; // @[hash.scala 41:22]
  reg [7:0] phv_data_137; // @[hash.scala 41:22]
  reg [7:0] phv_data_138; // @[hash.scala 41:22]
  reg [7:0] phv_data_139; // @[hash.scala 41:22]
  reg [7:0] phv_data_140; // @[hash.scala 41:22]
  reg [7:0] phv_data_141; // @[hash.scala 41:22]
  reg [7:0] phv_data_142; // @[hash.scala 41:22]
  reg [7:0] phv_data_143; // @[hash.scala 41:22]
  reg [7:0] phv_data_144; // @[hash.scala 41:22]
  reg [7:0] phv_data_145; // @[hash.scala 41:22]
  reg [7:0] phv_data_146; // @[hash.scala 41:22]
  reg [7:0] phv_data_147; // @[hash.scala 41:22]
  reg [7:0] phv_data_148; // @[hash.scala 41:22]
  reg [7:0] phv_data_149; // @[hash.scala 41:22]
  reg [7:0] phv_data_150; // @[hash.scala 41:22]
  reg [7:0] phv_data_151; // @[hash.scala 41:22]
  reg [7:0] phv_data_152; // @[hash.scala 41:22]
  reg [7:0] phv_data_153; // @[hash.scala 41:22]
  reg [7:0] phv_data_154; // @[hash.scala 41:22]
  reg [7:0] phv_data_155; // @[hash.scala 41:22]
  reg [7:0] phv_data_156; // @[hash.scala 41:22]
  reg [7:0] phv_data_157; // @[hash.scala 41:22]
  reg [7:0] phv_data_158; // @[hash.scala 41:22]
  reg [7:0] phv_data_159; // @[hash.scala 41:22]
  reg [7:0] phv_data_160; // @[hash.scala 41:22]
  reg [7:0] phv_data_161; // @[hash.scala 41:22]
  reg [7:0] phv_data_162; // @[hash.scala 41:22]
  reg [7:0] phv_data_163; // @[hash.scala 41:22]
  reg [7:0] phv_data_164; // @[hash.scala 41:22]
  reg [7:0] phv_data_165; // @[hash.scala 41:22]
  reg [7:0] phv_data_166; // @[hash.scala 41:22]
  reg [7:0] phv_data_167; // @[hash.scala 41:22]
  reg [7:0] phv_data_168; // @[hash.scala 41:22]
  reg [7:0] phv_data_169; // @[hash.scala 41:22]
  reg [7:0] phv_data_170; // @[hash.scala 41:22]
  reg [7:0] phv_data_171; // @[hash.scala 41:22]
  reg [7:0] phv_data_172; // @[hash.scala 41:22]
  reg [7:0] phv_data_173; // @[hash.scala 41:22]
  reg [7:0] phv_data_174; // @[hash.scala 41:22]
  reg [7:0] phv_data_175; // @[hash.scala 41:22]
  reg [7:0] phv_data_176; // @[hash.scala 41:22]
  reg [7:0] phv_data_177; // @[hash.scala 41:22]
  reg [7:0] phv_data_178; // @[hash.scala 41:22]
  reg [7:0] phv_data_179; // @[hash.scala 41:22]
  reg [7:0] phv_data_180; // @[hash.scala 41:22]
  reg [7:0] phv_data_181; // @[hash.scala 41:22]
  reg [7:0] phv_data_182; // @[hash.scala 41:22]
  reg [7:0] phv_data_183; // @[hash.scala 41:22]
  reg [7:0] phv_data_184; // @[hash.scala 41:22]
  reg [7:0] phv_data_185; // @[hash.scala 41:22]
  reg [7:0] phv_data_186; // @[hash.scala 41:22]
  reg [7:0] phv_data_187; // @[hash.scala 41:22]
  reg [7:0] phv_data_188; // @[hash.scala 41:22]
  reg [7:0] phv_data_189; // @[hash.scala 41:22]
  reg [7:0] phv_data_190; // @[hash.scala 41:22]
  reg [7:0] phv_data_191; // @[hash.scala 41:22]
  reg [7:0] phv_data_192; // @[hash.scala 41:22]
  reg [7:0] phv_data_193; // @[hash.scala 41:22]
  reg [7:0] phv_data_194; // @[hash.scala 41:22]
  reg [7:0] phv_data_195; // @[hash.scala 41:22]
  reg [7:0] phv_data_196; // @[hash.scala 41:22]
  reg [7:0] phv_data_197; // @[hash.scala 41:22]
  reg [7:0] phv_data_198; // @[hash.scala 41:22]
  reg [7:0] phv_data_199; // @[hash.scala 41:22]
  reg [7:0] phv_data_200; // @[hash.scala 41:22]
  reg [7:0] phv_data_201; // @[hash.scala 41:22]
  reg [7:0] phv_data_202; // @[hash.scala 41:22]
  reg [7:0] phv_data_203; // @[hash.scala 41:22]
  reg [7:0] phv_data_204; // @[hash.scala 41:22]
  reg [7:0] phv_data_205; // @[hash.scala 41:22]
  reg [7:0] phv_data_206; // @[hash.scala 41:22]
  reg [7:0] phv_data_207; // @[hash.scala 41:22]
  reg [7:0] phv_data_208; // @[hash.scala 41:22]
  reg [7:0] phv_data_209; // @[hash.scala 41:22]
  reg [7:0] phv_data_210; // @[hash.scala 41:22]
  reg [7:0] phv_data_211; // @[hash.scala 41:22]
  reg [7:0] phv_data_212; // @[hash.scala 41:22]
  reg [7:0] phv_data_213; // @[hash.scala 41:22]
  reg [7:0] phv_data_214; // @[hash.scala 41:22]
  reg [7:0] phv_data_215; // @[hash.scala 41:22]
  reg [7:0] phv_data_216; // @[hash.scala 41:22]
  reg [7:0] phv_data_217; // @[hash.scala 41:22]
  reg [7:0] phv_data_218; // @[hash.scala 41:22]
  reg [7:0] phv_data_219; // @[hash.scala 41:22]
  reg [7:0] phv_data_220; // @[hash.scala 41:22]
  reg [7:0] phv_data_221; // @[hash.scala 41:22]
  reg [7:0] phv_data_222; // @[hash.scala 41:22]
  reg [7:0] phv_data_223; // @[hash.scala 41:22]
  reg [7:0] phv_data_224; // @[hash.scala 41:22]
  reg [7:0] phv_data_225; // @[hash.scala 41:22]
  reg [7:0] phv_data_226; // @[hash.scala 41:22]
  reg [7:0] phv_data_227; // @[hash.scala 41:22]
  reg [7:0] phv_data_228; // @[hash.scala 41:22]
  reg [7:0] phv_data_229; // @[hash.scala 41:22]
  reg [7:0] phv_data_230; // @[hash.scala 41:22]
  reg [7:0] phv_data_231; // @[hash.scala 41:22]
  reg [7:0] phv_data_232; // @[hash.scala 41:22]
  reg [7:0] phv_data_233; // @[hash.scala 41:22]
  reg [7:0] phv_data_234; // @[hash.scala 41:22]
  reg [7:0] phv_data_235; // @[hash.scala 41:22]
  reg [7:0] phv_data_236; // @[hash.scala 41:22]
  reg [7:0] phv_data_237; // @[hash.scala 41:22]
  reg [7:0] phv_data_238; // @[hash.scala 41:22]
  reg [7:0] phv_data_239; // @[hash.scala 41:22]
  reg [7:0] phv_data_240; // @[hash.scala 41:22]
  reg [7:0] phv_data_241; // @[hash.scala 41:22]
  reg [7:0] phv_data_242; // @[hash.scala 41:22]
  reg [7:0] phv_data_243; // @[hash.scala 41:22]
  reg [7:0] phv_data_244; // @[hash.scala 41:22]
  reg [7:0] phv_data_245; // @[hash.scala 41:22]
  reg [7:0] phv_data_246; // @[hash.scala 41:22]
  reg [7:0] phv_data_247; // @[hash.scala 41:22]
  reg [7:0] phv_data_248; // @[hash.scala 41:22]
  reg [7:0] phv_data_249; // @[hash.scala 41:22]
  reg [7:0] phv_data_250; // @[hash.scala 41:22]
  reg [7:0] phv_data_251; // @[hash.scala 41:22]
  reg [7:0] phv_data_252; // @[hash.scala 41:22]
  reg [7:0] phv_data_253; // @[hash.scala 41:22]
  reg [7:0] phv_data_254; // @[hash.scala 41:22]
  reg [7:0] phv_data_255; // @[hash.scala 41:22]
  reg [7:0] phv_data_256; // @[hash.scala 41:22]
  reg [7:0] phv_data_257; // @[hash.scala 41:22]
  reg [7:0] phv_data_258; // @[hash.scala 41:22]
  reg [7:0] phv_data_259; // @[hash.scala 41:22]
  reg [7:0] phv_data_260; // @[hash.scala 41:22]
  reg [7:0] phv_data_261; // @[hash.scala 41:22]
  reg [7:0] phv_data_262; // @[hash.scala 41:22]
  reg [7:0] phv_data_263; // @[hash.scala 41:22]
  reg [7:0] phv_data_264; // @[hash.scala 41:22]
  reg [7:0] phv_data_265; // @[hash.scala 41:22]
  reg [7:0] phv_data_266; // @[hash.scala 41:22]
  reg [7:0] phv_data_267; // @[hash.scala 41:22]
  reg [7:0] phv_data_268; // @[hash.scala 41:22]
  reg [7:0] phv_data_269; // @[hash.scala 41:22]
  reg [7:0] phv_data_270; // @[hash.scala 41:22]
  reg [7:0] phv_data_271; // @[hash.scala 41:22]
  reg [7:0] phv_data_272; // @[hash.scala 41:22]
  reg [7:0] phv_data_273; // @[hash.scala 41:22]
  reg [7:0] phv_data_274; // @[hash.scala 41:22]
  reg [7:0] phv_data_275; // @[hash.scala 41:22]
  reg [7:0] phv_data_276; // @[hash.scala 41:22]
  reg [7:0] phv_data_277; // @[hash.scala 41:22]
  reg [7:0] phv_data_278; // @[hash.scala 41:22]
  reg [7:0] phv_data_279; // @[hash.scala 41:22]
  reg [7:0] phv_data_280; // @[hash.scala 41:22]
  reg [7:0] phv_data_281; // @[hash.scala 41:22]
  reg [7:0] phv_data_282; // @[hash.scala 41:22]
  reg [7:0] phv_data_283; // @[hash.scala 41:22]
  reg [7:0] phv_data_284; // @[hash.scala 41:22]
  reg [7:0] phv_data_285; // @[hash.scala 41:22]
  reg [7:0] phv_data_286; // @[hash.scala 41:22]
  reg [7:0] phv_data_287; // @[hash.scala 41:22]
  reg [7:0] phv_data_288; // @[hash.scala 41:22]
  reg [7:0] phv_data_289; // @[hash.scala 41:22]
  reg [7:0] phv_data_290; // @[hash.scala 41:22]
  reg [7:0] phv_data_291; // @[hash.scala 41:22]
  reg [7:0] phv_data_292; // @[hash.scala 41:22]
  reg [7:0] phv_data_293; // @[hash.scala 41:22]
  reg [7:0] phv_data_294; // @[hash.scala 41:22]
  reg [7:0] phv_data_295; // @[hash.scala 41:22]
  reg [7:0] phv_data_296; // @[hash.scala 41:22]
  reg [7:0] phv_data_297; // @[hash.scala 41:22]
  reg [7:0] phv_data_298; // @[hash.scala 41:22]
  reg [7:0] phv_data_299; // @[hash.scala 41:22]
  reg [7:0] phv_data_300; // @[hash.scala 41:22]
  reg [7:0] phv_data_301; // @[hash.scala 41:22]
  reg [7:0] phv_data_302; // @[hash.scala 41:22]
  reg [7:0] phv_data_303; // @[hash.scala 41:22]
  reg [7:0] phv_data_304; // @[hash.scala 41:22]
  reg [7:0] phv_data_305; // @[hash.scala 41:22]
  reg [7:0] phv_data_306; // @[hash.scala 41:22]
  reg [7:0] phv_data_307; // @[hash.scala 41:22]
  reg [7:0] phv_data_308; // @[hash.scala 41:22]
  reg [7:0] phv_data_309; // @[hash.scala 41:22]
  reg [7:0] phv_data_310; // @[hash.scala 41:22]
  reg [7:0] phv_data_311; // @[hash.scala 41:22]
  reg [7:0] phv_data_312; // @[hash.scala 41:22]
  reg [7:0] phv_data_313; // @[hash.scala 41:22]
  reg [7:0] phv_data_314; // @[hash.scala 41:22]
  reg [7:0] phv_data_315; // @[hash.scala 41:22]
  reg [7:0] phv_data_316; // @[hash.scala 41:22]
  reg [7:0] phv_data_317; // @[hash.scala 41:22]
  reg [7:0] phv_data_318; // @[hash.scala 41:22]
  reg [7:0] phv_data_319; // @[hash.scala 41:22]
  reg [7:0] phv_data_320; // @[hash.scala 41:22]
  reg [7:0] phv_data_321; // @[hash.scala 41:22]
  reg [7:0] phv_data_322; // @[hash.scala 41:22]
  reg [7:0] phv_data_323; // @[hash.scala 41:22]
  reg [7:0] phv_data_324; // @[hash.scala 41:22]
  reg [7:0] phv_data_325; // @[hash.scala 41:22]
  reg [7:0] phv_data_326; // @[hash.scala 41:22]
  reg [7:0] phv_data_327; // @[hash.scala 41:22]
  reg [7:0] phv_data_328; // @[hash.scala 41:22]
  reg [7:0] phv_data_329; // @[hash.scala 41:22]
  reg [7:0] phv_data_330; // @[hash.scala 41:22]
  reg [7:0] phv_data_331; // @[hash.scala 41:22]
  reg [7:0] phv_data_332; // @[hash.scala 41:22]
  reg [7:0] phv_data_333; // @[hash.scala 41:22]
  reg [7:0] phv_data_334; // @[hash.scala 41:22]
  reg [7:0] phv_data_335; // @[hash.scala 41:22]
  reg [7:0] phv_data_336; // @[hash.scala 41:22]
  reg [7:0] phv_data_337; // @[hash.scala 41:22]
  reg [7:0] phv_data_338; // @[hash.scala 41:22]
  reg [7:0] phv_data_339; // @[hash.scala 41:22]
  reg [7:0] phv_data_340; // @[hash.scala 41:22]
  reg [7:0] phv_data_341; // @[hash.scala 41:22]
  reg [7:0] phv_data_342; // @[hash.scala 41:22]
  reg [7:0] phv_data_343; // @[hash.scala 41:22]
  reg [7:0] phv_data_344; // @[hash.scala 41:22]
  reg [7:0] phv_data_345; // @[hash.scala 41:22]
  reg [7:0] phv_data_346; // @[hash.scala 41:22]
  reg [7:0] phv_data_347; // @[hash.scala 41:22]
  reg [7:0] phv_data_348; // @[hash.scala 41:22]
  reg [7:0] phv_data_349; // @[hash.scala 41:22]
  reg [7:0] phv_data_350; // @[hash.scala 41:22]
  reg [7:0] phv_data_351; // @[hash.scala 41:22]
  reg [7:0] phv_data_352; // @[hash.scala 41:22]
  reg [7:0] phv_data_353; // @[hash.scala 41:22]
  reg [7:0] phv_data_354; // @[hash.scala 41:22]
  reg [7:0] phv_data_355; // @[hash.scala 41:22]
  reg [7:0] phv_data_356; // @[hash.scala 41:22]
  reg [7:0] phv_data_357; // @[hash.scala 41:22]
  reg [7:0] phv_data_358; // @[hash.scala 41:22]
  reg [7:0] phv_data_359; // @[hash.scala 41:22]
  reg [7:0] phv_data_360; // @[hash.scala 41:22]
  reg [7:0] phv_data_361; // @[hash.scala 41:22]
  reg [7:0] phv_data_362; // @[hash.scala 41:22]
  reg [7:0] phv_data_363; // @[hash.scala 41:22]
  reg [7:0] phv_data_364; // @[hash.scala 41:22]
  reg [7:0] phv_data_365; // @[hash.scala 41:22]
  reg [7:0] phv_data_366; // @[hash.scala 41:22]
  reg [7:0] phv_data_367; // @[hash.scala 41:22]
  reg [7:0] phv_data_368; // @[hash.scala 41:22]
  reg [7:0] phv_data_369; // @[hash.scala 41:22]
  reg [7:0] phv_data_370; // @[hash.scala 41:22]
  reg [7:0] phv_data_371; // @[hash.scala 41:22]
  reg [7:0] phv_data_372; // @[hash.scala 41:22]
  reg [7:0] phv_data_373; // @[hash.scala 41:22]
  reg [7:0] phv_data_374; // @[hash.scala 41:22]
  reg [7:0] phv_data_375; // @[hash.scala 41:22]
  reg [7:0] phv_data_376; // @[hash.scala 41:22]
  reg [7:0] phv_data_377; // @[hash.scala 41:22]
  reg [7:0] phv_data_378; // @[hash.scala 41:22]
  reg [7:0] phv_data_379; // @[hash.scala 41:22]
  reg [7:0] phv_data_380; // @[hash.scala 41:22]
  reg [7:0] phv_data_381; // @[hash.scala 41:22]
  reg [7:0] phv_data_382; // @[hash.scala 41:22]
  reg [7:0] phv_data_383; // @[hash.scala 41:22]
  reg [7:0] phv_data_384; // @[hash.scala 41:22]
  reg [7:0] phv_data_385; // @[hash.scala 41:22]
  reg [7:0] phv_data_386; // @[hash.scala 41:22]
  reg [7:0] phv_data_387; // @[hash.scala 41:22]
  reg [7:0] phv_data_388; // @[hash.scala 41:22]
  reg [7:0] phv_data_389; // @[hash.scala 41:22]
  reg [7:0] phv_data_390; // @[hash.scala 41:22]
  reg [7:0] phv_data_391; // @[hash.scala 41:22]
  reg [7:0] phv_data_392; // @[hash.scala 41:22]
  reg [7:0] phv_data_393; // @[hash.scala 41:22]
  reg [7:0] phv_data_394; // @[hash.scala 41:22]
  reg [7:0] phv_data_395; // @[hash.scala 41:22]
  reg [7:0] phv_data_396; // @[hash.scala 41:22]
  reg [7:0] phv_data_397; // @[hash.scala 41:22]
  reg [7:0] phv_data_398; // @[hash.scala 41:22]
  reg [7:0] phv_data_399; // @[hash.scala 41:22]
  reg [7:0] phv_data_400; // @[hash.scala 41:22]
  reg [7:0] phv_data_401; // @[hash.scala 41:22]
  reg [7:0] phv_data_402; // @[hash.scala 41:22]
  reg [7:0] phv_data_403; // @[hash.scala 41:22]
  reg [7:0] phv_data_404; // @[hash.scala 41:22]
  reg [7:0] phv_data_405; // @[hash.scala 41:22]
  reg [7:0] phv_data_406; // @[hash.scala 41:22]
  reg [7:0] phv_data_407; // @[hash.scala 41:22]
  reg [7:0] phv_data_408; // @[hash.scala 41:22]
  reg [7:0] phv_data_409; // @[hash.scala 41:22]
  reg [7:0] phv_data_410; // @[hash.scala 41:22]
  reg [7:0] phv_data_411; // @[hash.scala 41:22]
  reg [7:0] phv_data_412; // @[hash.scala 41:22]
  reg [7:0] phv_data_413; // @[hash.scala 41:22]
  reg [7:0] phv_data_414; // @[hash.scala 41:22]
  reg [7:0] phv_data_415; // @[hash.scala 41:22]
  reg [7:0] phv_data_416; // @[hash.scala 41:22]
  reg [7:0] phv_data_417; // @[hash.scala 41:22]
  reg [7:0] phv_data_418; // @[hash.scala 41:22]
  reg [7:0] phv_data_419; // @[hash.scala 41:22]
  reg [7:0] phv_data_420; // @[hash.scala 41:22]
  reg [7:0] phv_data_421; // @[hash.scala 41:22]
  reg [7:0] phv_data_422; // @[hash.scala 41:22]
  reg [7:0] phv_data_423; // @[hash.scala 41:22]
  reg [7:0] phv_data_424; // @[hash.scala 41:22]
  reg [7:0] phv_data_425; // @[hash.scala 41:22]
  reg [7:0] phv_data_426; // @[hash.scala 41:22]
  reg [7:0] phv_data_427; // @[hash.scala 41:22]
  reg [7:0] phv_data_428; // @[hash.scala 41:22]
  reg [7:0] phv_data_429; // @[hash.scala 41:22]
  reg [7:0] phv_data_430; // @[hash.scala 41:22]
  reg [7:0] phv_data_431; // @[hash.scala 41:22]
  reg [7:0] phv_data_432; // @[hash.scala 41:22]
  reg [7:0] phv_data_433; // @[hash.scala 41:22]
  reg [7:0] phv_data_434; // @[hash.scala 41:22]
  reg [7:0] phv_data_435; // @[hash.scala 41:22]
  reg [7:0] phv_data_436; // @[hash.scala 41:22]
  reg [7:0] phv_data_437; // @[hash.scala 41:22]
  reg [7:0] phv_data_438; // @[hash.scala 41:22]
  reg [7:0] phv_data_439; // @[hash.scala 41:22]
  reg [7:0] phv_data_440; // @[hash.scala 41:22]
  reg [7:0] phv_data_441; // @[hash.scala 41:22]
  reg [7:0] phv_data_442; // @[hash.scala 41:22]
  reg [7:0] phv_data_443; // @[hash.scala 41:22]
  reg [7:0] phv_data_444; // @[hash.scala 41:22]
  reg [7:0] phv_data_445; // @[hash.scala 41:22]
  reg [7:0] phv_data_446; // @[hash.scala 41:22]
  reg [7:0] phv_data_447; // @[hash.scala 41:22]
  reg [7:0] phv_data_448; // @[hash.scala 41:22]
  reg [7:0] phv_data_449; // @[hash.scala 41:22]
  reg [7:0] phv_data_450; // @[hash.scala 41:22]
  reg [7:0] phv_data_451; // @[hash.scala 41:22]
  reg [7:0] phv_data_452; // @[hash.scala 41:22]
  reg [7:0] phv_data_453; // @[hash.scala 41:22]
  reg [7:0] phv_data_454; // @[hash.scala 41:22]
  reg [7:0] phv_data_455; // @[hash.scala 41:22]
  reg [7:0] phv_data_456; // @[hash.scala 41:22]
  reg [7:0] phv_data_457; // @[hash.scala 41:22]
  reg [7:0] phv_data_458; // @[hash.scala 41:22]
  reg [7:0] phv_data_459; // @[hash.scala 41:22]
  reg [7:0] phv_data_460; // @[hash.scala 41:22]
  reg [7:0] phv_data_461; // @[hash.scala 41:22]
  reg [7:0] phv_data_462; // @[hash.scala 41:22]
  reg [7:0] phv_data_463; // @[hash.scala 41:22]
  reg [7:0] phv_data_464; // @[hash.scala 41:22]
  reg [7:0] phv_data_465; // @[hash.scala 41:22]
  reg [7:0] phv_data_466; // @[hash.scala 41:22]
  reg [7:0] phv_data_467; // @[hash.scala 41:22]
  reg [7:0] phv_data_468; // @[hash.scala 41:22]
  reg [7:0] phv_data_469; // @[hash.scala 41:22]
  reg [7:0] phv_data_470; // @[hash.scala 41:22]
  reg [7:0] phv_data_471; // @[hash.scala 41:22]
  reg [7:0] phv_data_472; // @[hash.scala 41:22]
  reg [7:0] phv_data_473; // @[hash.scala 41:22]
  reg [7:0] phv_data_474; // @[hash.scala 41:22]
  reg [7:0] phv_data_475; // @[hash.scala 41:22]
  reg [7:0] phv_data_476; // @[hash.scala 41:22]
  reg [7:0] phv_data_477; // @[hash.scala 41:22]
  reg [7:0] phv_data_478; // @[hash.scala 41:22]
  reg [7:0] phv_data_479; // @[hash.scala 41:22]
  reg [7:0] phv_data_480; // @[hash.scala 41:22]
  reg [7:0] phv_data_481; // @[hash.scala 41:22]
  reg [7:0] phv_data_482; // @[hash.scala 41:22]
  reg [7:0] phv_data_483; // @[hash.scala 41:22]
  reg [7:0] phv_data_484; // @[hash.scala 41:22]
  reg [7:0] phv_data_485; // @[hash.scala 41:22]
  reg [7:0] phv_data_486; // @[hash.scala 41:22]
  reg [7:0] phv_data_487; // @[hash.scala 41:22]
  reg [7:0] phv_data_488; // @[hash.scala 41:22]
  reg [7:0] phv_data_489; // @[hash.scala 41:22]
  reg [7:0] phv_data_490; // @[hash.scala 41:22]
  reg [7:0] phv_data_491; // @[hash.scala 41:22]
  reg [7:0] phv_data_492; // @[hash.scala 41:22]
  reg [7:0] phv_data_493; // @[hash.scala 41:22]
  reg [7:0] phv_data_494; // @[hash.scala 41:22]
  reg [7:0] phv_data_495; // @[hash.scala 41:22]
  reg [7:0] phv_data_496; // @[hash.scala 41:22]
  reg [7:0] phv_data_497; // @[hash.scala 41:22]
  reg [7:0] phv_data_498; // @[hash.scala 41:22]
  reg [7:0] phv_data_499; // @[hash.scala 41:22]
  reg [7:0] phv_data_500; // @[hash.scala 41:22]
  reg [7:0] phv_data_501; // @[hash.scala 41:22]
  reg [7:0] phv_data_502; // @[hash.scala 41:22]
  reg [7:0] phv_data_503; // @[hash.scala 41:22]
  reg [7:0] phv_data_504; // @[hash.scala 41:22]
  reg [7:0] phv_data_505; // @[hash.scala 41:22]
  reg [7:0] phv_data_506; // @[hash.scala 41:22]
  reg [7:0] phv_data_507; // @[hash.scala 41:22]
  reg [7:0] phv_data_508; // @[hash.scala 41:22]
  reg [7:0] phv_data_509; // @[hash.scala 41:22]
  reg [7:0] phv_data_510; // @[hash.scala 41:22]
  reg [7:0] phv_data_511; // @[hash.scala 41:22]
  reg [15:0] phv_header_0; // @[hash.scala 41:22]
  reg [15:0] phv_header_1; // @[hash.scala 41:22]
  reg [15:0] phv_header_2; // @[hash.scala 41:22]
  reg [15:0] phv_header_3; // @[hash.scala 41:22]
  reg [15:0] phv_header_4; // @[hash.scala 41:22]
  reg [15:0] phv_header_5; // @[hash.scala 41:22]
  reg [15:0] phv_header_6; // @[hash.scala 41:22]
  reg [15:0] phv_header_7; // @[hash.scala 41:22]
  reg [15:0] phv_header_8; // @[hash.scala 41:22]
  reg [15:0] phv_header_9; // @[hash.scala 41:22]
  reg [15:0] phv_header_10; // @[hash.scala 41:22]
  reg [15:0] phv_header_11; // @[hash.scala 41:22]
  reg [15:0] phv_header_12; // @[hash.scala 41:22]
  reg [15:0] phv_header_13; // @[hash.scala 41:22]
  reg [15:0] phv_header_14; // @[hash.scala 41:22]
  reg [15:0] phv_header_15; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 41:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 41:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 41:22]
  reg  phv_next_config_id; // @[hash.scala 41:22]
  reg  phv_is_valid_processor; // @[hash.scala 41:22]
  reg [191:0] key; // @[hash.scala 45:22]
  reg [191:0] sum; // @[hash.scala 49:22]
  wire [15:0] sum_temp_0 = sum[15:0]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_1 = sum[31:16]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_2 = sum[47:32]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_3 = sum[63:48]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_4 = sum[79:64]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_5 = sum[95:80]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_6 = sum[111:96]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_7 = sum[127:112]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_8 = sum[143:128]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_9 = sum[159:144]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_10 = sum[175:160]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_11 = sum[191:176]; // @[hash.scala 64:35]
  wire [15:0] out_temp_0 = sum_temp_0 + sum_temp_1; // @[hash.scala 70:51]
  wire [15:0] out_temp_1 = sum_temp_2 + sum_temp_3; // @[hash.scala 70:51]
  wire [15:0] out_temp_2 = sum_temp_4 + sum_temp_5; // @[hash.scala 70:51]
  wire [15:0] out_temp_3 = sum_temp_6 + sum_temp_7; // @[hash.scala 70:51]
  wire [15:0] out_temp_4 = sum_temp_8 + sum_temp_9; // @[hash.scala 70:51]
  wire [15:0] out_temp_5 = sum_temp_10 + sum_temp_11; // @[hash.scala 70:51]
  wire [95:0] _io_sum_out_T = {out_temp_0,out_temp_1,out_temp_2,out_temp_3,out_temp_4,out_temp_5}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_160 = phv_data_160; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_161 = phv_data_161; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_162 = phv_data_162; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_163 = phv_data_163; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_164 = phv_data_164; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_165 = phv_data_165; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_166 = phv_data_166; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_167 = phv_data_167; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_168 = phv_data_168; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_169 = phv_data_169; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_170 = phv_data_170; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_171 = phv_data_171; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_172 = phv_data_172; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_173 = phv_data_173; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_174 = phv_data_174; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_175 = phv_data_175; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_176 = phv_data_176; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_177 = phv_data_177; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_178 = phv_data_178; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_179 = phv_data_179; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_180 = phv_data_180; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_181 = phv_data_181; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_182 = phv_data_182; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_183 = phv_data_183; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_184 = phv_data_184; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_185 = phv_data_185; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_186 = phv_data_186; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_187 = phv_data_187; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_188 = phv_data_188; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_189 = phv_data_189; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_190 = phv_data_190; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_191 = phv_data_191; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_192 = phv_data_192; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_193 = phv_data_193; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_194 = phv_data_194; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_195 = phv_data_195; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_196 = phv_data_196; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_197 = phv_data_197; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_198 = phv_data_198; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_199 = phv_data_199; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_200 = phv_data_200; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_201 = phv_data_201; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_202 = phv_data_202; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_203 = phv_data_203; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_204 = phv_data_204; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_205 = phv_data_205; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_206 = phv_data_206; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_207 = phv_data_207; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_208 = phv_data_208; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_209 = phv_data_209; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_210 = phv_data_210; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_211 = phv_data_211; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_212 = phv_data_212; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_213 = phv_data_213; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_214 = phv_data_214; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_215 = phv_data_215; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_216 = phv_data_216; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_217 = phv_data_217; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_218 = phv_data_218; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_219 = phv_data_219; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_220 = phv_data_220; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_221 = phv_data_221; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_222 = phv_data_222; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_223 = phv_data_223; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_224 = phv_data_224; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_225 = phv_data_225; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_226 = phv_data_226; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_227 = phv_data_227; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_228 = phv_data_228; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_229 = phv_data_229; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_230 = phv_data_230; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_231 = phv_data_231; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_232 = phv_data_232; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_233 = phv_data_233; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_234 = phv_data_234; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_235 = phv_data_235; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_236 = phv_data_236; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_237 = phv_data_237; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_238 = phv_data_238; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_239 = phv_data_239; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_240 = phv_data_240; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_241 = phv_data_241; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_242 = phv_data_242; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_243 = phv_data_243; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_244 = phv_data_244; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_245 = phv_data_245; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_246 = phv_data_246; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_247 = phv_data_247; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_248 = phv_data_248; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_249 = phv_data_249; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_250 = phv_data_250; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_251 = phv_data_251; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_252 = phv_data_252; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_253 = phv_data_253; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_254 = phv_data_254; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_255 = phv_data_255; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_256 = phv_data_256; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_257 = phv_data_257; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_258 = phv_data_258; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_259 = phv_data_259; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_260 = phv_data_260; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_261 = phv_data_261; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_262 = phv_data_262; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_263 = phv_data_263; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_264 = phv_data_264; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_265 = phv_data_265; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_266 = phv_data_266; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_267 = phv_data_267; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_268 = phv_data_268; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_269 = phv_data_269; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_270 = phv_data_270; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_271 = phv_data_271; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_272 = phv_data_272; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_273 = phv_data_273; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_274 = phv_data_274; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_275 = phv_data_275; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_276 = phv_data_276; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_277 = phv_data_277; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_278 = phv_data_278; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_279 = phv_data_279; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_280 = phv_data_280; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_281 = phv_data_281; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_282 = phv_data_282; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_283 = phv_data_283; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_284 = phv_data_284; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_285 = phv_data_285; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_286 = phv_data_286; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_287 = phv_data_287; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_288 = phv_data_288; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_289 = phv_data_289; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_290 = phv_data_290; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_291 = phv_data_291; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_292 = phv_data_292; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_293 = phv_data_293; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_294 = phv_data_294; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_295 = phv_data_295; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_296 = phv_data_296; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_297 = phv_data_297; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_298 = phv_data_298; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_299 = phv_data_299; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_300 = phv_data_300; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_301 = phv_data_301; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_302 = phv_data_302; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_303 = phv_data_303; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_304 = phv_data_304; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_305 = phv_data_305; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_306 = phv_data_306; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_307 = phv_data_307; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_308 = phv_data_308; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_309 = phv_data_309; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_310 = phv_data_310; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_311 = phv_data_311; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_312 = phv_data_312; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_313 = phv_data_313; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_314 = phv_data_314; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_315 = phv_data_315; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_316 = phv_data_316; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_317 = phv_data_317; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_318 = phv_data_318; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_319 = phv_data_319; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_320 = phv_data_320; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_321 = phv_data_321; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_322 = phv_data_322; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_323 = phv_data_323; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_324 = phv_data_324; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_325 = phv_data_325; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_326 = phv_data_326; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_327 = phv_data_327; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_328 = phv_data_328; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_329 = phv_data_329; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_330 = phv_data_330; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_331 = phv_data_331; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_332 = phv_data_332; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_333 = phv_data_333; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_334 = phv_data_334; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_335 = phv_data_335; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_336 = phv_data_336; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_337 = phv_data_337; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_338 = phv_data_338; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_339 = phv_data_339; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_340 = phv_data_340; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_341 = phv_data_341; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_342 = phv_data_342; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_343 = phv_data_343; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_344 = phv_data_344; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_345 = phv_data_345; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_346 = phv_data_346; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_347 = phv_data_347; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_348 = phv_data_348; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_349 = phv_data_349; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_350 = phv_data_350; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_351 = phv_data_351; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_352 = phv_data_352; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_353 = phv_data_353; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_354 = phv_data_354; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_355 = phv_data_355; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_356 = phv_data_356; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_357 = phv_data_357; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_358 = phv_data_358; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_359 = phv_data_359; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_360 = phv_data_360; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_361 = phv_data_361; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_362 = phv_data_362; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_363 = phv_data_363; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_364 = phv_data_364; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_365 = phv_data_365; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_366 = phv_data_366; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_367 = phv_data_367; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_368 = phv_data_368; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_369 = phv_data_369; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_370 = phv_data_370; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_371 = phv_data_371; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_372 = phv_data_372; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_373 = phv_data_373; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_374 = phv_data_374; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_375 = phv_data_375; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_376 = phv_data_376; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_377 = phv_data_377; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_378 = phv_data_378; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_379 = phv_data_379; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_380 = phv_data_380; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_381 = phv_data_381; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_382 = phv_data_382; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_383 = phv_data_383; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_384 = phv_data_384; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_385 = phv_data_385; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_386 = phv_data_386; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_387 = phv_data_387; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_388 = phv_data_388; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_389 = phv_data_389; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_390 = phv_data_390; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_391 = phv_data_391; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_392 = phv_data_392; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_393 = phv_data_393; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_394 = phv_data_394; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_395 = phv_data_395; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_396 = phv_data_396; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_397 = phv_data_397; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_398 = phv_data_398; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_399 = phv_data_399; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_400 = phv_data_400; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_401 = phv_data_401; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_402 = phv_data_402; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_403 = phv_data_403; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_404 = phv_data_404; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_405 = phv_data_405; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_406 = phv_data_406; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_407 = phv_data_407; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_408 = phv_data_408; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_409 = phv_data_409; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_410 = phv_data_410; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_411 = phv_data_411; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_412 = phv_data_412; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_413 = phv_data_413; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_414 = phv_data_414; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_415 = phv_data_415; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_416 = phv_data_416; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_417 = phv_data_417; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_418 = phv_data_418; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_419 = phv_data_419; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_420 = phv_data_420; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_421 = phv_data_421; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_422 = phv_data_422; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_423 = phv_data_423; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_424 = phv_data_424; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_425 = phv_data_425; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_426 = phv_data_426; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_427 = phv_data_427; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_428 = phv_data_428; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_429 = phv_data_429; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_430 = phv_data_430; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_431 = phv_data_431; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_432 = phv_data_432; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_433 = phv_data_433; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_434 = phv_data_434; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_435 = phv_data_435; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_436 = phv_data_436; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_437 = phv_data_437; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_438 = phv_data_438; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_439 = phv_data_439; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_440 = phv_data_440; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_441 = phv_data_441; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_442 = phv_data_442; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_443 = phv_data_443; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_444 = phv_data_444; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_445 = phv_data_445; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_446 = phv_data_446; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_447 = phv_data_447; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_448 = phv_data_448; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_449 = phv_data_449; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_450 = phv_data_450; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_451 = phv_data_451; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_452 = phv_data_452; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_453 = phv_data_453; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_454 = phv_data_454; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_455 = phv_data_455; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_456 = phv_data_456; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_457 = phv_data_457; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_458 = phv_data_458; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_459 = phv_data_459; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_460 = phv_data_460; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_461 = phv_data_461; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_462 = phv_data_462; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_463 = phv_data_463; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_464 = phv_data_464; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_465 = phv_data_465; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_466 = phv_data_466; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_467 = phv_data_467; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_468 = phv_data_468; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_469 = phv_data_469; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_470 = phv_data_470; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_471 = phv_data_471; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_472 = phv_data_472; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_473 = phv_data_473; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_474 = phv_data_474; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_475 = phv_data_475; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_476 = phv_data_476; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_477 = phv_data_477; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_478 = phv_data_478; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_479 = phv_data_479; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_480 = phv_data_480; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_481 = phv_data_481; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_482 = phv_data_482; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_483 = phv_data_483; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_484 = phv_data_484; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_485 = phv_data_485; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_486 = phv_data_486; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_487 = phv_data_487; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_488 = phv_data_488; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_489 = phv_data_489; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_490 = phv_data_490; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_491 = phv_data_491; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_492 = phv_data_492; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_493 = phv_data_493; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_494 = phv_data_494; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_495 = phv_data_495; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_496 = phv_data_496; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_497 = phv_data_497; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_498 = phv_data_498; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_499 = phv_data_499; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_500 = phv_data_500; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_501 = phv_data_501; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_502 = phv_data_502; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_503 = phv_data_503; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_504 = phv_data_504; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_505 = phv_data_505; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_506 = phv_data_506; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_507 = phv_data_507; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_508 = phv_data_508; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_509 = phv_data_509; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_510 = phv_data_510; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_511 = phv_data_511; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 43:25]
  assign io_key_out = key; // @[hash.scala 47:20]
  assign io_sum_out = phv_is_valid_processor ? {{96'd0}, _io_sum_out_T} : sum; // @[hash.scala 52:39 hash.scala 75:24 hash.scala 77:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 42:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 42:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 42:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 42:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 42:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 42:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 42:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 42:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 42:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 42:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 42:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 42:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 42:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 42:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 42:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 42:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 42:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 42:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 42:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 42:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 42:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 42:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 42:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 42:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 42:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 42:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 42:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 42:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 42:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 42:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 42:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 42:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 42:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 42:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 42:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 42:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 42:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 42:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 42:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 42:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 42:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 42:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 42:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 42:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 42:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 42:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 42:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 42:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 42:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 42:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 42:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 42:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 42:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 42:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 42:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 42:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 42:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 42:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 42:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 42:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 42:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 42:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 42:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 42:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 42:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 42:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 42:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 42:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 42:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 42:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 42:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 42:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 42:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 42:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 42:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 42:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 42:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 42:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 42:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 42:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 42:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 42:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 42:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 42:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 42:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 42:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 42:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 42:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 42:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 42:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 42:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 42:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 42:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 42:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 42:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 42:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 42:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 42:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 42:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 42:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 42:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 42:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 42:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 42:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 42:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 42:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 42:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 42:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 42:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 42:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 42:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 42:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 42:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 42:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 42:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 42:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 42:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 42:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 42:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 42:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 42:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 42:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 42:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 42:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 42:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 42:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 42:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 42:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 42:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 42:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 42:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 42:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 42:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 42:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 42:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 42:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 42:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 42:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 42:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 42:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 42:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 42:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 42:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 42:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 42:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 42:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 42:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 42:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 42:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 42:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 42:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 42:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 42:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 42:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 42:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 42:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 42:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 42:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 42:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 42:13]
    phv_data_160 <= io_pipe_phv_in_data_160; // @[hash.scala 42:13]
    phv_data_161 <= io_pipe_phv_in_data_161; // @[hash.scala 42:13]
    phv_data_162 <= io_pipe_phv_in_data_162; // @[hash.scala 42:13]
    phv_data_163 <= io_pipe_phv_in_data_163; // @[hash.scala 42:13]
    phv_data_164 <= io_pipe_phv_in_data_164; // @[hash.scala 42:13]
    phv_data_165 <= io_pipe_phv_in_data_165; // @[hash.scala 42:13]
    phv_data_166 <= io_pipe_phv_in_data_166; // @[hash.scala 42:13]
    phv_data_167 <= io_pipe_phv_in_data_167; // @[hash.scala 42:13]
    phv_data_168 <= io_pipe_phv_in_data_168; // @[hash.scala 42:13]
    phv_data_169 <= io_pipe_phv_in_data_169; // @[hash.scala 42:13]
    phv_data_170 <= io_pipe_phv_in_data_170; // @[hash.scala 42:13]
    phv_data_171 <= io_pipe_phv_in_data_171; // @[hash.scala 42:13]
    phv_data_172 <= io_pipe_phv_in_data_172; // @[hash.scala 42:13]
    phv_data_173 <= io_pipe_phv_in_data_173; // @[hash.scala 42:13]
    phv_data_174 <= io_pipe_phv_in_data_174; // @[hash.scala 42:13]
    phv_data_175 <= io_pipe_phv_in_data_175; // @[hash.scala 42:13]
    phv_data_176 <= io_pipe_phv_in_data_176; // @[hash.scala 42:13]
    phv_data_177 <= io_pipe_phv_in_data_177; // @[hash.scala 42:13]
    phv_data_178 <= io_pipe_phv_in_data_178; // @[hash.scala 42:13]
    phv_data_179 <= io_pipe_phv_in_data_179; // @[hash.scala 42:13]
    phv_data_180 <= io_pipe_phv_in_data_180; // @[hash.scala 42:13]
    phv_data_181 <= io_pipe_phv_in_data_181; // @[hash.scala 42:13]
    phv_data_182 <= io_pipe_phv_in_data_182; // @[hash.scala 42:13]
    phv_data_183 <= io_pipe_phv_in_data_183; // @[hash.scala 42:13]
    phv_data_184 <= io_pipe_phv_in_data_184; // @[hash.scala 42:13]
    phv_data_185 <= io_pipe_phv_in_data_185; // @[hash.scala 42:13]
    phv_data_186 <= io_pipe_phv_in_data_186; // @[hash.scala 42:13]
    phv_data_187 <= io_pipe_phv_in_data_187; // @[hash.scala 42:13]
    phv_data_188 <= io_pipe_phv_in_data_188; // @[hash.scala 42:13]
    phv_data_189 <= io_pipe_phv_in_data_189; // @[hash.scala 42:13]
    phv_data_190 <= io_pipe_phv_in_data_190; // @[hash.scala 42:13]
    phv_data_191 <= io_pipe_phv_in_data_191; // @[hash.scala 42:13]
    phv_data_192 <= io_pipe_phv_in_data_192; // @[hash.scala 42:13]
    phv_data_193 <= io_pipe_phv_in_data_193; // @[hash.scala 42:13]
    phv_data_194 <= io_pipe_phv_in_data_194; // @[hash.scala 42:13]
    phv_data_195 <= io_pipe_phv_in_data_195; // @[hash.scala 42:13]
    phv_data_196 <= io_pipe_phv_in_data_196; // @[hash.scala 42:13]
    phv_data_197 <= io_pipe_phv_in_data_197; // @[hash.scala 42:13]
    phv_data_198 <= io_pipe_phv_in_data_198; // @[hash.scala 42:13]
    phv_data_199 <= io_pipe_phv_in_data_199; // @[hash.scala 42:13]
    phv_data_200 <= io_pipe_phv_in_data_200; // @[hash.scala 42:13]
    phv_data_201 <= io_pipe_phv_in_data_201; // @[hash.scala 42:13]
    phv_data_202 <= io_pipe_phv_in_data_202; // @[hash.scala 42:13]
    phv_data_203 <= io_pipe_phv_in_data_203; // @[hash.scala 42:13]
    phv_data_204 <= io_pipe_phv_in_data_204; // @[hash.scala 42:13]
    phv_data_205 <= io_pipe_phv_in_data_205; // @[hash.scala 42:13]
    phv_data_206 <= io_pipe_phv_in_data_206; // @[hash.scala 42:13]
    phv_data_207 <= io_pipe_phv_in_data_207; // @[hash.scala 42:13]
    phv_data_208 <= io_pipe_phv_in_data_208; // @[hash.scala 42:13]
    phv_data_209 <= io_pipe_phv_in_data_209; // @[hash.scala 42:13]
    phv_data_210 <= io_pipe_phv_in_data_210; // @[hash.scala 42:13]
    phv_data_211 <= io_pipe_phv_in_data_211; // @[hash.scala 42:13]
    phv_data_212 <= io_pipe_phv_in_data_212; // @[hash.scala 42:13]
    phv_data_213 <= io_pipe_phv_in_data_213; // @[hash.scala 42:13]
    phv_data_214 <= io_pipe_phv_in_data_214; // @[hash.scala 42:13]
    phv_data_215 <= io_pipe_phv_in_data_215; // @[hash.scala 42:13]
    phv_data_216 <= io_pipe_phv_in_data_216; // @[hash.scala 42:13]
    phv_data_217 <= io_pipe_phv_in_data_217; // @[hash.scala 42:13]
    phv_data_218 <= io_pipe_phv_in_data_218; // @[hash.scala 42:13]
    phv_data_219 <= io_pipe_phv_in_data_219; // @[hash.scala 42:13]
    phv_data_220 <= io_pipe_phv_in_data_220; // @[hash.scala 42:13]
    phv_data_221 <= io_pipe_phv_in_data_221; // @[hash.scala 42:13]
    phv_data_222 <= io_pipe_phv_in_data_222; // @[hash.scala 42:13]
    phv_data_223 <= io_pipe_phv_in_data_223; // @[hash.scala 42:13]
    phv_data_224 <= io_pipe_phv_in_data_224; // @[hash.scala 42:13]
    phv_data_225 <= io_pipe_phv_in_data_225; // @[hash.scala 42:13]
    phv_data_226 <= io_pipe_phv_in_data_226; // @[hash.scala 42:13]
    phv_data_227 <= io_pipe_phv_in_data_227; // @[hash.scala 42:13]
    phv_data_228 <= io_pipe_phv_in_data_228; // @[hash.scala 42:13]
    phv_data_229 <= io_pipe_phv_in_data_229; // @[hash.scala 42:13]
    phv_data_230 <= io_pipe_phv_in_data_230; // @[hash.scala 42:13]
    phv_data_231 <= io_pipe_phv_in_data_231; // @[hash.scala 42:13]
    phv_data_232 <= io_pipe_phv_in_data_232; // @[hash.scala 42:13]
    phv_data_233 <= io_pipe_phv_in_data_233; // @[hash.scala 42:13]
    phv_data_234 <= io_pipe_phv_in_data_234; // @[hash.scala 42:13]
    phv_data_235 <= io_pipe_phv_in_data_235; // @[hash.scala 42:13]
    phv_data_236 <= io_pipe_phv_in_data_236; // @[hash.scala 42:13]
    phv_data_237 <= io_pipe_phv_in_data_237; // @[hash.scala 42:13]
    phv_data_238 <= io_pipe_phv_in_data_238; // @[hash.scala 42:13]
    phv_data_239 <= io_pipe_phv_in_data_239; // @[hash.scala 42:13]
    phv_data_240 <= io_pipe_phv_in_data_240; // @[hash.scala 42:13]
    phv_data_241 <= io_pipe_phv_in_data_241; // @[hash.scala 42:13]
    phv_data_242 <= io_pipe_phv_in_data_242; // @[hash.scala 42:13]
    phv_data_243 <= io_pipe_phv_in_data_243; // @[hash.scala 42:13]
    phv_data_244 <= io_pipe_phv_in_data_244; // @[hash.scala 42:13]
    phv_data_245 <= io_pipe_phv_in_data_245; // @[hash.scala 42:13]
    phv_data_246 <= io_pipe_phv_in_data_246; // @[hash.scala 42:13]
    phv_data_247 <= io_pipe_phv_in_data_247; // @[hash.scala 42:13]
    phv_data_248 <= io_pipe_phv_in_data_248; // @[hash.scala 42:13]
    phv_data_249 <= io_pipe_phv_in_data_249; // @[hash.scala 42:13]
    phv_data_250 <= io_pipe_phv_in_data_250; // @[hash.scala 42:13]
    phv_data_251 <= io_pipe_phv_in_data_251; // @[hash.scala 42:13]
    phv_data_252 <= io_pipe_phv_in_data_252; // @[hash.scala 42:13]
    phv_data_253 <= io_pipe_phv_in_data_253; // @[hash.scala 42:13]
    phv_data_254 <= io_pipe_phv_in_data_254; // @[hash.scala 42:13]
    phv_data_255 <= io_pipe_phv_in_data_255; // @[hash.scala 42:13]
    phv_data_256 <= io_pipe_phv_in_data_256; // @[hash.scala 42:13]
    phv_data_257 <= io_pipe_phv_in_data_257; // @[hash.scala 42:13]
    phv_data_258 <= io_pipe_phv_in_data_258; // @[hash.scala 42:13]
    phv_data_259 <= io_pipe_phv_in_data_259; // @[hash.scala 42:13]
    phv_data_260 <= io_pipe_phv_in_data_260; // @[hash.scala 42:13]
    phv_data_261 <= io_pipe_phv_in_data_261; // @[hash.scala 42:13]
    phv_data_262 <= io_pipe_phv_in_data_262; // @[hash.scala 42:13]
    phv_data_263 <= io_pipe_phv_in_data_263; // @[hash.scala 42:13]
    phv_data_264 <= io_pipe_phv_in_data_264; // @[hash.scala 42:13]
    phv_data_265 <= io_pipe_phv_in_data_265; // @[hash.scala 42:13]
    phv_data_266 <= io_pipe_phv_in_data_266; // @[hash.scala 42:13]
    phv_data_267 <= io_pipe_phv_in_data_267; // @[hash.scala 42:13]
    phv_data_268 <= io_pipe_phv_in_data_268; // @[hash.scala 42:13]
    phv_data_269 <= io_pipe_phv_in_data_269; // @[hash.scala 42:13]
    phv_data_270 <= io_pipe_phv_in_data_270; // @[hash.scala 42:13]
    phv_data_271 <= io_pipe_phv_in_data_271; // @[hash.scala 42:13]
    phv_data_272 <= io_pipe_phv_in_data_272; // @[hash.scala 42:13]
    phv_data_273 <= io_pipe_phv_in_data_273; // @[hash.scala 42:13]
    phv_data_274 <= io_pipe_phv_in_data_274; // @[hash.scala 42:13]
    phv_data_275 <= io_pipe_phv_in_data_275; // @[hash.scala 42:13]
    phv_data_276 <= io_pipe_phv_in_data_276; // @[hash.scala 42:13]
    phv_data_277 <= io_pipe_phv_in_data_277; // @[hash.scala 42:13]
    phv_data_278 <= io_pipe_phv_in_data_278; // @[hash.scala 42:13]
    phv_data_279 <= io_pipe_phv_in_data_279; // @[hash.scala 42:13]
    phv_data_280 <= io_pipe_phv_in_data_280; // @[hash.scala 42:13]
    phv_data_281 <= io_pipe_phv_in_data_281; // @[hash.scala 42:13]
    phv_data_282 <= io_pipe_phv_in_data_282; // @[hash.scala 42:13]
    phv_data_283 <= io_pipe_phv_in_data_283; // @[hash.scala 42:13]
    phv_data_284 <= io_pipe_phv_in_data_284; // @[hash.scala 42:13]
    phv_data_285 <= io_pipe_phv_in_data_285; // @[hash.scala 42:13]
    phv_data_286 <= io_pipe_phv_in_data_286; // @[hash.scala 42:13]
    phv_data_287 <= io_pipe_phv_in_data_287; // @[hash.scala 42:13]
    phv_data_288 <= io_pipe_phv_in_data_288; // @[hash.scala 42:13]
    phv_data_289 <= io_pipe_phv_in_data_289; // @[hash.scala 42:13]
    phv_data_290 <= io_pipe_phv_in_data_290; // @[hash.scala 42:13]
    phv_data_291 <= io_pipe_phv_in_data_291; // @[hash.scala 42:13]
    phv_data_292 <= io_pipe_phv_in_data_292; // @[hash.scala 42:13]
    phv_data_293 <= io_pipe_phv_in_data_293; // @[hash.scala 42:13]
    phv_data_294 <= io_pipe_phv_in_data_294; // @[hash.scala 42:13]
    phv_data_295 <= io_pipe_phv_in_data_295; // @[hash.scala 42:13]
    phv_data_296 <= io_pipe_phv_in_data_296; // @[hash.scala 42:13]
    phv_data_297 <= io_pipe_phv_in_data_297; // @[hash.scala 42:13]
    phv_data_298 <= io_pipe_phv_in_data_298; // @[hash.scala 42:13]
    phv_data_299 <= io_pipe_phv_in_data_299; // @[hash.scala 42:13]
    phv_data_300 <= io_pipe_phv_in_data_300; // @[hash.scala 42:13]
    phv_data_301 <= io_pipe_phv_in_data_301; // @[hash.scala 42:13]
    phv_data_302 <= io_pipe_phv_in_data_302; // @[hash.scala 42:13]
    phv_data_303 <= io_pipe_phv_in_data_303; // @[hash.scala 42:13]
    phv_data_304 <= io_pipe_phv_in_data_304; // @[hash.scala 42:13]
    phv_data_305 <= io_pipe_phv_in_data_305; // @[hash.scala 42:13]
    phv_data_306 <= io_pipe_phv_in_data_306; // @[hash.scala 42:13]
    phv_data_307 <= io_pipe_phv_in_data_307; // @[hash.scala 42:13]
    phv_data_308 <= io_pipe_phv_in_data_308; // @[hash.scala 42:13]
    phv_data_309 <= io_pipe_phv_in_data_309; // @[hash.scala 42:13]
    phv_data_310 <= io_pipe_phv_in_data_310; // @[hash.scala 42:13]
    phv_data_311 <= io_pipe_phv_in_data_311; // @[hash.scala 42:13]
    phv_data_312 <= io_pipe_phv_in_data_312; // @[hash.scala 42:13]
    phv_data_313 <= io_pipe_phv_in_data_313; // @[hash.scala 42:13]
    phv_data_314 <= io_pipe_phv_in_data_314; // @[hash.scala 42:13]
    phv_data_315 <= io_pipe_phv_in_data_315; // @[hash.scala 42:13]
    phv_data_316 <= io_pipe_phv_in_data_316; // @[hash.scala 42:13]
    phv_data_317 <= io_pipe_phv_in_data_317; // @[hash.scala 42:13]
    phv_data_318 <= io_pipe_phv_in_data_318; // @[hash.scala 42:13]
    phv_data_319 <= io_pipe_phv_in_data_319; // @[hash.scala 42:13]
    phv_data_320 <= io_pipe_phv_in_data_320; // @[hash.scala 42:13]
    phv_data_321 <= io_pipe_phv_in_data_321; // @[hash.scala 42:13]
    phv_data_322 <= io_pipe_phv_in_data_322; // @[hash.scala 42:13]
    phv_data_323 <= io_pipe_phv_in_data_323; // @[hash.scala 42:13]
    phv_data_324 <= io_pipe_phv_in_data_324; // @[hash.scala 42:13]
    phv_data_325 <= io_pipe_phv_in_data_325; // @[hash.scala 42:13]
    phv_data_326 <= io_pipe_phv_in_data_326; // @[hash.scala 42:13]
    phv_data_327 <= io_pipe_phv_in_data_327; // @[hash.scala 42:13]
    phv_data_328 <= io_pipe_phv_in_data_328; // @[hash.scala 42:13]
    phv_data_329 <= io_pipe_phv_in_data_329; // @[hash.scala 42:13]
    phv_data_330 <= io_pipe_phv_in_data_330; // @[hash.scala 42:13]
    phv_data_331 <= io_pipe_phv_in_data_331; // @[hash.scala 42:13]
    phv_data_332 <= io_pipe_phv_in_data_332; // @[hash.scala 42:13]
    phv_data_333 <= io_pipe_phv_in_data_333; // @[hash.scala 42:13]
    phv_data_334 <= io_pipe_phv_in_data_334; // @[hash.scala 42:13]
    phv_data_335 <= io_pipe_phv_in_data_335; // @[hash.scala 42:13]
    phv_data_336 <= io_pipe_phv_in_data_336; // @[hash.scala 42:13]
    phv_data_337 <= io_pipe_phv_in_data_337; // @[hash.scala 42:13]
    phv_data_338 <= io_pipe_phv_in_data_338; // @[hash.scala 42:13]
    phv_data_339 <= io_pipe_phv_in_data_339; // @[hash.scala 42:13]
    phv_data_340 <= io_pipe_phv_in_data_340; // @[hash.scala 42:13]
    phv_data_341 <= io_pipe_phv_in_data_341; // @[hash.scala 42:13]
    phv_data_342 <= io_pipe_phv_in_data_342; // @[hash.scala 42:13]
    phv_data_343 <= io_pipe_phv_in_data_343; // @[hash.scala 42:13]
    phv_data_344 <= io_pipe_phv_in_data_344; // @[hash.scala 42:13]
    phv_data_345 <= io_pipe_phv_in_data_345; // @[hash.scala 42:13]
    phv_data_346 <= io_pipe_phv_in_data_346; // @[hash.scala 42:13]
    phv_data_347 <= io_pipe_phv_in_data_347; // @[hash.scala 42:13]
    phv_data_348 <= io_pipe_phv_in_data_348; // @[hash.scala 42:13]
    phv_data_349 <= io_pipe_phv_in_data_349; // @[hash.scala 42:13]
    phv_data_350 <= io_pipe_phv_in_data_350; // @[hash.scala 42:13]
    phv_data_351 <= io_pipe_phv_in_data_351; // @[hash.scala 42:13]
    phv_data_352 <= io_pipe_phv_in_data_352; // @[hash.scala 42:13]
    phv_data_353 <= io_pipe_phv_in_data_353; // @[hash.scala 42:13]
    phv_data_354 <= io_pipe_phv_in_data_354; // @[hash.scala 42:13]
    phv_data_355 <= io_pipe_phv_in_data_355; // @[hash.scala 42:13]
    phv_data_356 <= io_pipe_phv_in_data_356; // @[hash.scala 42:13]
    phv_data_357 <= io_pipe_phv_in_data_357; // @[hash.scala 42:13]
    phv_data_358 <= io_pipe_phv_in_data_358; // @[hash.scala 42:13]
    phv_data_359 <= io_pipe_phv_in_data_359; // @[hash.scala 42:13]
    phv_data_360 <= io_pipe_phv_in_data_360; // @[hash.scala 42:13]
    phv_data_361 <= io_pipe_phv_in_data_361; // @[hash.scala 42:13]
    phv_data_362 <= io_pipe_phv_in_data_362; // @[hash.scala 42:13]
    phv_data_363 <= io_pipe_phv_in_data_363; // @[hash.scala 42:13]
    phv_data_364 <= io_pipe_phv_in_data_364; // @[hash.scala 42:13]
    phv_data_365 <= io_pipe_phv_in_data_365; // @[hash.scala 42:13]
    phv_data_366 <= io_pipe_phv_in_data_366; // @[hash.scala 42:13]
    phv_data_367 <= io_pipe_phv_in_data_367; // @[hash.scala 42:13]
    phv_data_368 <= io_pipe_phv_in_data_368; // @[hash.scala 42:13]
    phv_data_369 <= io_pipe_phv_in_data_369; // @[hash.scala 42:13]
    phv_data_370 <= io_pipe_phv_in_data_370; // @[hash.scala 42:13]
    phv_data_371 <= io_pipe_phv_in_data_371; // @[hash.scala 42:13]
    phv_data_372 <= io_pipe_phv_in_data_372; // @[hash.scala 42:13]
    phv_data_373 <= io_pipe_phv_in_data_373; // @[hash.scala 42:13]
    phv_data_374 <= io_pipe_phv_in_data_374; // @[hash.scala 42:13]
    phv_data_375 <= io_pipe_phv_in_data_375; // @[hash.scala 42:13]
    phv_data_376 <= io_pipe_phv_in_data_376; // @[hash.scala 42:13]
    phv_data_377 <= io_pipe_phv_in_data_377; // @[hash.scala 42:13]
    phv_data_378 <= io_pipe_phv_in_data_378; // @[hash.scala 42:13]
    phv_data_379 <= io_pipe_phv_in_data_379; // @[hash.scala 42:13]
    phv_data_380 <= io_pipe_phv_in_data_380; // @[hash.scala 42:13]
    phv_data_381 <= io_pipe_phv_in_data_381; // @[hash.scala 42:13]
    phv_data_382 <= io_pipe_phv_in_data_382; // @[hash.scala 42:13]
    phv_data_383 <= io_pipe_phv_in_data_383; // @[hash.scala 42:13]
    phv_data_384 <= io_pipe_phv_in_data_384; // @[hash.scala 42:13]
    phv_data_385 <= io_pipe_phv_in_data_385; // @[hash.scala 42:13]
    phv_data_386 <= io_pipe_phv_in_data_386; // @[hash.scala 42:13]
    phv_data_387 <= io_pipe_phv_in_data_387; // @[hash.scala 42:13]
    phv_data_388 <= io_pipe_phv_in_data_388; // @[hash.scala 42:13]
    phv_data_389 <= io_pipe_phv_in_data_389; // @[hash.scala 42:13]
    phv_data_390 <= io_pipe_phv_in_data_390; // @[hash.scala 42:13]
    phv_data_391 <= io_pipe_phv_in_data_391; // @[hash.scala 42:13]
    phv_data_392 <= io_pipe_phv_in_data_392; // @[hash.scala 42:13]
    phv_data_393 <= io_pipe_phv_in_data_393; // @[hash.scala 42:13]
    phv_data_394 <= io_pipe_phv_in_data_394; // @[hash.scala 42:13]
    phv_data_395 <= io_pipe_phv_in_data_395; // @[hash.scala 42:13]
    phv_data_396 <= io_pipe_phv_in_data_396; // @[hash.scala 42:13]
    phv_data_397 <= io_pipe_phv_in_data_397; // @[hash.scala 42:13]
    phv_data_398 <= io_pipe_phv_in_data_398; // @[hash.scala 42:13]
    phv_data_399 <= io_pipe_phv_in_data_399; // @[hash.scala 42:13]
    phv_data_400 <= io_pipe_phv_in_data_400; // @[hash.scala 42:13]
    phv_data_401 <= io_pipe_phv_in_data_401; // @[hash.scala 42:13]
    phv_data_402 <= io_pipe_phv_in_data_402; // @[hash.scala 42:13]
    phv_data_403 <= io_pipe_phv_in_data_403; // @[hash.scala 42:13]
    phv_data_404 <= io_pipe_phv_in_data_404; // @[hash.scala 42:13]
    phv_data_405 <= io_pipe_phv_in_data_405; // @[hash.scala 42:13]
    phv_data_406 <= io_pipe_phv_in_data_406; // @[hash.scala 42:13]
    phv_data_407 <= io_pipe_phv_in_data_407; // @[hash.scala 42:13]
    phv_data_408 <= io_pipe_phv_in_data_408; // @[hash.scala 42:13]
    phv_data_409 <= io_pipe_phv_in_data_409; // @[hash.scala 42:13]
    phv_data_410 <= io_pipe_phv_in_data_410; // @[hash.scala 42:13]
    phv_data_411 <= io_pipe_phv_in_data_411; // @[hash.scala 42:13]
    phv_data_412 <= io_pipe_phv_in_data_412; // @[hash.scala 42:13]
    phv_data_413 <= io_pipe_phv_in_data_413; // @[hash.scala 42:13]
    phv_data_414 <= io_pipe_phv_in_data_414; // @[hash.scala 42:13]
    phv_data_415 <= io_pipe_phv_in_data_415; // @[hash.scala 42:13]
    phv_data_416 <= io_pipe_phv_in_data_416; // @[hash.scala 42:13]
    phv_data_417 <= io_pipe_phv_in_data_417; // @[hash.scala 42:13]
    phv_data_418 <= io_pipe_phv_in_data_418; // @[hash.scala 42:13]
    phv_data_419 <= io_pipe_phv_in_data_419; // @[hash.scala 42:13]
    phv_data_420 <= io_pipe_phv_in_data_420; // @[hash.scala 42:13]
    phv_data_421 <= io_pipe_phv_in_data_421; // @[hash.scala 42:13]
    phv_data_422 <= io_pipe_phv_in_data_422; // @[hash.scala 42:13]
    phv_data_423 <= io_pipe_phv_in_data_423; // @[hash.scala 42:13]
    phv_data_424 <= io_pipe_phv_in_data_424; // @[hash.scala 42:13]
    phv_data_425 <= io_pipe_phv_in_data_425; // @[hash.scala 42:13]
    phv_data_426 <= io_pipe_phv_in_data_426; // @[hash.scala 42:13]
    phv_data_427 <= io_pipe_phv_in_data_427; // @[hash.scala 42:13]
    phv_data_428 <= io_pipe_phv_in_data_428; // @[hash.scala 42:13]
    phv_data_429 <= io_pipe_phv_in_data_429; // @[hash.scala 42:13]
    phv_data_430 <= io_pipe_phv_in_data_430; // @[hash.scala 42:13]
    phv_data_431 <= io_pipe_phv_in_data_431; // @[hash.scala 42:13]
    phv_data_432 <= io_pipe_phv_in_data_432; // @[hash.scala 42:13]
    phv_data_433 <= io_pipe_phv_in_data_433; // @[hash.scala 42:13]
    phv_data_434 <= io_pipe_phv_in_data_434; // @[hash.scala 42:13]
    phv_data_435 <= io_pipe_phv_in_data_435; // @[hash.scala 42:13]
    phv_data_436 <= io_pipe_phv_in_data_436; // @[hash.scala 42:13]
    phv_data_437 <= io_pipe_phv_in_data_437; // @[hash.scala 42:13]
    phv_data_438 <= io_pipe_phv_in_data_438; // @[hash.scala 42:13]
    phv_data_439 <= io_pipe_phv_in_data_439; // @[hash.scala 42:13]
    phv_data_440 <= io_pipe_phv_in_data_440; // @[hash.scala 42:13]
    phv_data_441 <= io_pipe_phv_in_data_441; // @[hash.scala 42:13]
    phv_data_442 <= io_pipe_phv_in_data_442; // @[hash.scala 42:13]
    phv_data_443 <= io_pipe_phv_in_data_443; // @[hash.scala 42:13]
    phv_data_444 <= io_pipe_phv_in_data_444; // @[hash.scala 42:13]
    phv_data_445 <= io_pipe_phv_in_data_445; // @[hash.scala 42:13]
    phv_data_446 <= io_pipe_phv_in_data_446; // @[hash.scala 42:13]
    phv_data_447 <= io_pipe_phv_in_data_447; // @[hash.scala 42:13]
    phv_data_448 <= io_pipe_phv_in_data_448; // @[hash.scala 42:13]
    phv_data_449 <= io_pipe_phv_in_data_449; // @[hash.scala 42:13]
    phv_data_450 <= io_pipe_phv_in_data_450; // @[hash.scala 42:13]
    phv_data_451 <= io_pipe_phv_in_data_451; // @[hash.scala 42:13]
    phv_data_452 <= io_pipe_phv_in_data_452; // @[hash.scala 42:13]
    phv_data_453 <= io_pipe_phv_in_data_453; // @[hash.scala 42:13]
    phv_data_454 <= io_pipe_phv_in_data_454; // @[hash.scala 42:13]
    phv_data_455 <= io_pipe_phv_in_data_455; // @[hash.scala 42:13]
    phv_data_456 <= io_pipe_phv_in_data_456; // @[hash.scala 42:13]
    phv_data_457 <= io_pipe_phv_in_data_457; // @[hash.scala 42:13]
    phv_data_458 <= io_pipe_phv_in_data_458; // @[hash.scala 42:13]
    phv_data_459 <= io_pipe_phv_in_data_459; // @[hash.scala 42:13]
    phv_data_460 <= io_pipe_phv_in_data_460; // @[hash.scala 42:13]
    phv_data_461 <= io_pipe_phv_in_data_461; // @[hash.scala 42:13]
    phv_data_462 <= io_pipe_phv_in_data_462; // @[hash.scala 42:13]
    phv_data_463 <= io_pipe_phv_in_data_463; // @[hash.scala 42:13]
    phv_data_464 <= io_pipe_phv_in_data_464; // @[hash.scala 42:13]
    phv_data_465 <= io_pipe_phv_in_data_465; // @[hash.scala 42:13]
    phv_data_466 <= io_pipe_phv_in_data_466; // @[hash.scala 42:13]
    phv_data_467 <= io_pipe_phv_in_data_467; // @[hash.scala 42:13]
    phv_data_468 <= io_pipe_phv_in_data_468; // @[hash.scala 42:13]
    phv_data_469 <= io_pipe_phv_in_data_469; // @[hash.scala 42:13]
    phv_data_470 <= io_pipe_phv_in_data_470; // @[hash.scala 42:13]
    phv_data_471 <= io_pipe_phv_in_data_471; // @[hash.scala 42:13]
    phv_data_472 <= io_pipe_phv_in_data_472; // @[hash.scala 42:13]
    phv_data_473 <= io_pipe_phv_in_data_473; // @[hash.scala 42:13]
    phv_data_474 <= io_pipe_phv_in_data_474; // @[hash.scala 42:13]
    phv_data_475 <= io_pipe_phv_in_data_475; // @[hash.scala 42:13]
    phv_data_476 <= io_pipe_phv_in_data_476; // @[hash.scala 42:13]
    phv_data_477 <= io_pipe_phv_in_data_477; // @[hash.scala 42:13]
    phv_data_478 <= io_pipe_phv_in_data_478; // @[hash.scala 42:13]
    phv_data_479 <= io_pipe_phv_in_data_479; // @[hash.scala 42:13]
    phv_data_480 <= io_pipe_phv_in_data_480; // @[hash.scala 42:13]
    phv_data_481 <= io_pipe_phv_in_data_481; // @[hash.scala 42:13]
    phv_data_482 <= io_pipe_phv_in_data_482; // @[hash.scala 42:13]
    phv_data_483 <= io_pipe_phv_in_data_483; // @[hash.scala 42:13]
    phv_data_484 <= io_pipe_phv_in_data_484; // @[hash.scala 42:13]
    phv_data_485 <= io_pipe_phv_in_data_485; // @[hash.scala 42:13]
    phv_data_486 <= io_pipe_phv_in_data_486; // @[hash.scala 42:13]
    phv_data_487 <= io_pipe_phv_in_data_487; // @[hash.scala 42:13]
    phv_data_488 <= io_pipe_phv_in_data_488; // @[hash.scala 42:13]
    phv_data_489 <= io_pipe_phv_in_data_489; // @[hash.scala 42:13]
    phv_data_490 <= io_pipe_phv_in_data_490; // @[hash.scala 42:13]
    phv_data_491 <= io_pipe_phv_in_data_491; // @[hash.scala 42:13]
    phv_data_492 <= io_pipe_phv_in_data_492; // @[hash.scala 42:13]
    phv_data_493 <= io_pipe_phv_in_data_493; // @[hash.scala 42:13]
    phv_data_494 <= io_pipe_phv_in_data_494; // @[hash.scala 42:13]
    phv_data_495 <= io_pipe_phv_in_data_495; // @[hash.scala 42:13]
    phv_data_496 <= io_pipe_phv_in_data_496; // @[hash.scala 42:13]
    phv_data_497 <= io_pipe_phv_in_data_497; // @[hash.scala 42:13]
    phv_data_498 <= io_pipe_phv_in_data_498; // @[hash.scala 42:13]
    phv_data_499 <= io_pipe_phv_in_data_499; // @[hash.scala 42:13]
    phv_data_500 <= io_pipe_phv_in_data_500; // @[hash.scala 42:13]
    phv_data_501 <= io_pipe_phv_in_data_501; // @[hash.scala 42:13]
    phv_data_502 <= io_pipe_phv_in_data_502; // @[hash.scala 42:13]
    phv_data_503 <= io_pipe_phv_in_data_503; // @[hash.scala 42:13]
    phv_data_504 <= io_pipe_phv_in_data_504; // @[hash.scala 42:13]
    phv_data_505 <= io_pipe_phv_in_data_505; // @[hash.scala 42:13]
    phv_data_506 <= io_pipe_phv_in_data_506; // @[hash.scala 42:13]
    phv_data_507 <= io_pipe_phv_in_data_507; // @[hash.scala 42:13]
    phv_data_508 <= io_pipe_phv_in_data_508; // @[hash.scala 42:13]
    phv_data_509 <= io_pipe_phv_in_data_509; // @[hash.scala 42:13]
    phv_data_510 <= io_pipe_phv_in_data_510; // @[hash.scala 42:13]
    phv_data_511 <= io_pipe_phv_in_data_511; // @[hash.scala 42:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 42:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 42:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 42:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 42:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 42:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 42:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 42:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 42:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 42:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 42:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 42:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 42:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 42:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 42:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 42:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 42:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 42:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 42:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 42:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 42:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 42:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 42:13]
    key <= io_key_in; // @[hash.scala 46:13]
    sum <= io_sum_in; // @[hash.scala 50:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_data_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  phv_data_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  phv_data_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  phv_data_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  phv_data_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  phv_data_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  phv_data_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  phv_data_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  phv_data_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  phv_data_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  phv_data_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  phv_data_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  phv_data_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  phv_data_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  phv_data_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  phv_data_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  phv_data_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_data_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_data_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  phv_data_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  phv_data_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  phv_data_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  phv_data_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  phv_data_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  phv_data_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  phv_data_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  phv_data_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  phv_data_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  phv_data_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  phv_data_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  phv_data_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  phv_data_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  phv_data_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  phv_data_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  phv_data_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  phv_data_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  phv_data_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  phv_data_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  phv_data_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  phv_data_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  phv_data_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  phv_data_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  phv_data_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  phv_data_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  phv_data_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  phv_data_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  phv_data_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  phv_data_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  phv_data_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  phv_data_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  phv_data_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  phv_data_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  phv_data_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  phv_data_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  phv_data_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  phv_data_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  phv_data_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  phv_data_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  phv_data_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  phv_data_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  phv_data_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  phv_data_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  phv_data_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  phv_data_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  phv_data_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  phv_data_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  phv_data_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  phv_data_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  phv_data_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  phv_data_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  phv_data_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  phv_data_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  phv_data_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  phv_data_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  phv_data_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  phv_data_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  phv_data_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  phv_data_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  phv_data_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  phv_data_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  phv_data_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  phv_data_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  phv_data_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  phv_data_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  phv_data_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  phv_data_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  phv_data_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  phv_data_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  phv_data_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  phv_data_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  phv_data_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  phv_data_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  phv_data_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  phv_data_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  phv_data_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  phv_data_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  phv_data_256 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  phv_data_257 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  phv_data_258 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  phv_data_259 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  phv_data_260 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  phv_data_261 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  phv_data_262 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  phv_data_263 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  phv_data_264 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  phv_data_265 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  phv_data_266 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  phv_data_267 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  phv_data_268 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  phv_data_269 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  phv_data_270 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  phv_data_271 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  phv_data_272 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  phv_data_273 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  phv_data_274 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  phv_data_275 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  phv_data_276 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  phv_data_277 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  phv_data_278 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  phv_data_279 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  phv_data_280 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  phv_data_281 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  phv_data_282 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  phv_data_283 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  phv_data_284 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  phv_data_285 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  phv_data_286 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  phv_data_287 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  phv_data_288 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  phv_data_289 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  phv_data_290 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  phv_data_291 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  phv_data_292 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  phv_data_293 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  phv_data_294 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  phv_data_295 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  phv_data_296 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  phv_data_297 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  phv_data_298 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  phv_data_299 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  phv_data_300 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  phv_data_301 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  phv_data_302 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  phv_data_303 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  phv_data_304 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  phv_data_305 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  phv_data_306 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  phv_data_307 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  phv_data_308 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  phv_data_309 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  phv_data_310 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  phv_data_311 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  phv_data_312 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  phv_data_313 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  phv_data_314 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  phv_data_315 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  phv_data_316 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  phv_data_317 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  phv_data_318 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  phv_data_319 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  phv_data_320 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  phv_data_321 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  phv_data_322 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  phv_data_323 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  phv_data_324 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  phv_data_325 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  phv_data_326 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  phv_data_327 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  phv_data_328 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  phv_data_329 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  phv_data_330 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  phv_data_331 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  phv_data_332 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  phv_data_333 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  phv_data_334 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  phv_data_335 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  phv_data_336 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  phv_data_337 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  phv_data_338 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  phv_data_339 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  phv_data_340 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  phv_data_341 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  phv_data_342 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  phv_data_343 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  phv_data_344 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  phv_data_345 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  phv_data_346 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  phv_data_347 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  phv_data_348 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  phv_data_349 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  phv_data_350 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  phv_data_351 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  phv_data_352 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  phv_data_353 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  phv_data_354 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  phv_data_355 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  phv_data_356 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  phv_data_357 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  phv_data_358 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  phv_data_359 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  phv_data_360 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  phv_data_361 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  phv_data_362 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  phv_data_363 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  phv_data_364 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  phv_data_365 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  phv_data_366 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  phv_data_367 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  phv_data_368 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  phv_data_369 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  phv_data_370 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  phv_data_371 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  phv_data_372 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  phv_data_373 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  phv_data_374 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  phv_data_375 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  phv_data_376 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  phv_data_377 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  phv_data_378 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  phv_data_379 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  phv_data_380 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  phv_data_381 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  phv_data_382 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  phv_data_383 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  phv_data_384 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  phv_data_385 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  phv_data_386 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  phv_data_387 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  phv_data_388 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  phv_data_389 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  phv_data_390 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  phv_data_391 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  phv_data_392 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  phv_data_393 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  phv_data_394 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  phv_data_395 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  phv_data_396 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  phv_data_397 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  phv_data_398 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  phv_data_399 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  phv_data_400 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  phv_data_401 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  phv_data_402 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  phv_data_403 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  phv_data_404 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  phv_data_405 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  phv_data_406 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  phv_data_407 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  phv_data_408 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  phv_data_409 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  phv_data_410 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  phv_data_411 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  phv_data_412 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  phv_data_413 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  phv_data_414 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  phv_data_415 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  phv_data_416 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  phv_data_417 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  phv_data_418 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  phv_data_419 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  phv_data_420 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  phv_data_421 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  phv_data_422 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  phv_data_423 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  phv_data_424 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  phv_data_425 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  phv_data_426 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  phv_data_427 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  phv_data_428 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  phv_data_429 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  phv_data_430 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  phv_data_431 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  phv_data_432 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  phv_data_433 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  phv_data_434 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  phv_data_435 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  phv_data_436 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  phv_data_437 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  phv_data_438 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  phv_data_439 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  phv_data_440 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  phv_data_441 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  phv_data_442 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  phv_data_443 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  phv_data_444 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  phv_data_445 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  phv_data_446 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  phv_data_447 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  phv_data_448 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  phv_data_449 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  phv_data_450 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  phv_data_451 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  phv_data_452 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  phv_data_453 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  phv_data_454 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  phv_data_455 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  phv_data_456 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  phv_data_457 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  phv_data_458 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  phv_data_459 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  phv_data_460 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  phv_data_461 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  phv_data_462 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  phv_data_463 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  phv_data_464 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  phv_data_465 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  phv_data_466 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  phv_data_467 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  phv_data_468 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  phv_data_469 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  phv_data_470 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  phv_data_471 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  phv_data_472 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  phv_data_473 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  phv_data_474 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  phv_data_475 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  phv_data_476 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  phv_data_477 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  phv_data_478 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  phv_data_479 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  phv_data_480 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  phv_data_481 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  phv_data_482 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  phv_data_483 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  phv_data_484 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  phv_data_485 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  phv_data_486 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  phv_data_487 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  phv_data_488 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  phv_data_489 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  phv_data_490 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  phv_data_491 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  phv_data_492 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  phv_data_493 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  phv_data_494 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  phv_data_495 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  phv_data_496 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  phv_data_497 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  phv_data_498 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  phv_data_499 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  phv_data_500 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  phv_data_501 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  phv_data_502 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  phv_data_503 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  phv_data_504 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  phv_data_505 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  phv_data_506 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  phv_data_507 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  phv_data_508 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  phv_data_509 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  phv_data_510 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  phv_data_511 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  phv_header_0 = _RAND_512[15:0];
  _RAND_513 = {1{`RANDOM}};
  phv_header_1 = _RAND_513[15:0];
  _RAND_514 = {1{`RANDOM}};
  phv_header_2 = _RAND_514[15:0];
  _RAND_515 = {1{`RANDOM}};
  phv_header_3 = _RAND_515[15:0];
  _RAND_516 = {1{`RANDOM}};
  phv_header_4 = _RAND_516[15:0];
  _RAND_517 = {1{`RANDOM}};
  phv_header_5 = _RAND_517[15:0];
  _RAND_518 = {1{`RANDOM}};
  phv_header_6 = _RAND_518[15:0];
  _RAND_519 = {1{`RANDOM}};
  phv_header_7 = _RAND_519[15:0];
  _RAND_520 = {1{`RANDOM}};
  phv_header_8 = _RAND_520[15:0];
  _RAND_521 = {1{`RANDOM}};
  phv_header_9 = _RAND_521[15:0];
  _RAND_522 = {1{`RANDOM}};
  phv_header_10 = _RAND_522[15:0];
  _RAND_523 = {1{`RANDOM}};
  phv_header_11 = _RAND_523[15:0];
  _RAND_524 = {1{`RANDOM}};
  phv_header_12 = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  phv_header_13 = _RAND_525[15:0];
  _RAND_526 = {1{`RANDOM}};
  phv_header_14 = _RAND_526[15:0];
  _RAND_527 = {1{`RANDOM}};
  phv_header_15 = _RAND_527[15:0];
  _RAND_528 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_530[15:0];
  _RAND_531 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  phv_next_config_id = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_533[0:0];
  _RAND_534 = {6{`RANDOM}};
  key = _RAND_534[191:0];
  _RAND_535 = {6{`RANDOM}};
  sum = _RAND_535[191:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
