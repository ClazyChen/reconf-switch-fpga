module MatchGetKeyPISA(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [1:0]   io_key_config_0_field_config_0,
  input  [1:0]   io_key_config_0_field_config_1,
  input  [1:0]   io_key_config_0_field_config_2,
  input  [1:0]   io_key_config_0_field_config_3,
  input  [1:0]   io_key_config_0_field_config_4,
  input  [1:0]   io_key_config_0_field_config_5,
  input          io_key_config_0_field_mask_0_0,
  input          io_key_config_0_field_mask_0_1,
  input          io_key_config_0_field_mask_0_2,
  input          io_key_config_0_field_mask_0_3,
  input          io_key_config_0_field_mask_1_0,
  input          io_key_config_0_field_mask_1_1,
  input          io_key_config_0_field_mask_1_2,
  input          io_key_config_0_field_mask_1_3,
  input          io_key_config_0_field_mask_2_0,
  input          io_key_config_0_field_mask_2_1,
  input          io_key_config_0_field_mask_2_2,
  input          io_key_config_0_field_mask_2_3,
  input          io_key_config_0_field_mask_3_0,
  input          io_key_config_0_field_mask_3_1,
  input          io_key_config_0_field_mask_3_2,
  input          io_key_config_0_field_mask_3_3,
  input          io_key_config_0_field_mask_4_0,
  input          io_key_config_0_field_mask_4_1,
  input          io_key_config_0_field_mask_4_2,
  input          io_key_config_0_field_mask_4_3,
  input          io_key_config_0_field_mask_5_0,
  input          io_key_config_0_field_mask_5_1,
  input          io_key_config_0_field_mask_5_2,
  input          io_key_config_0_field_mask_5_3,
  input  [6:0]   io_key_config_0_field_id_0_0,
  input  [6:0]   io_key_config_0_field_id_0_1,
  input  [6:0]   io_key_config_0_field_id_0_2,
  input  [6:0]   io_key_config_0_field_id_0_3,
  input  [6:0]   io_key_config_0_field_id_1_0,
  input  [6:0]   io_key_config_0_field_id_1_1,
  input  [6:0]   io_key_config_0_field_id_1_2,
  input  [6:0]   io_key_config_0_field_id_1_3,
  input  [6:0]   io_key_config_0_field_id_2_0,
  input  [6:0]   io_key_config_0_field_id_2_1,
  input  [6:0]   io_key_config_0_field_id_2_2,
  input  [6:0]   io_key_config_0_field_id_2_3,
  input  [6:0]   io_key_config_0_field_id_3_0,
  input  [6:0]   io_key_config_0_field_id_3_1,
  input  [6:0]   io_key_config_0_field_id_3_2,
  input  [6:0]   io_key_config_0_field_id_3_3,
  input  [6:0]   io_key_config_0_field_id_4_0,
  input  [6:0]   io_key_config_0_field_id_4_1,
  input  [6:0]   io_key_config_0_field_id_4_2,
  input  [6:0]   io_key_config_0_field_id_4_3,
  input  [6:0]   io_key_config_0_field_id_5_0,
  input  [6:0]   io_key_config_0_field_id_5_1,
  input  [6:0]   io_key_config_0_field_id_5_2,
  input  [6:0]   io_key_config_0_field_id_5_3,
  input  [1:0]   io_key_config_1_field_config_0,
  input  [1:0]   io_key_config_1_field_config_1,
  input  [1:0]   io_key_config_1_field_config_2,
  input  [1:0]   io_key_config_1_field_config_3,
  input  [1:0]   io_key_config_1_field_config_4,
  input  [1:0]   io_key_config_1_field_config_5,
  input          io_key_config_1_field_mask_0_0,
  input          io_key_config_1_field_mask_0_1,
  input          io_key_config_1_field_mask_0_2,
  input          io_key_config_1_field_mask_0_3,
  input          io_key_config_1_field_mask_1_0,
  input          io_key_config_1_field_mask_1_1,
  input          io_key_config_1_field_mask_1_2,
  input          io_key_config_1_field_mask_1_3,
  input          io_key_config_1_field_mask_2_0,
  input          io_key_config_1_field_mask_2_1,
  input          io_key_config_1_field_mask_2_2,
  input          io_key_config_1_field_mask_2_3,
  input          io_key_config_1_field_mask_3_0,
  input          io_key_config_1_field_mask_3_1,
  input          io_key_config_1_field_mask_3_2,
  input          io_key_config_1_field_mask_3_3,
  input          io_key_config_1_field_mask_4_0,
  input          io_key_config_1_field_mask_4_1,
  input          io_key_config_1_field_mask_4_2,
  input          io_key_config_1_field_mask_4_3,
  input          io_key_config_1_field_mask_5_0,
  input          io_key_config_1_field_mask_5_1,
  input          io_key_config_1_field_mask_5_2,
  input          io_key_config_1_field_mask_5_3,
  input  [6:0]   io_key_config_1_field_id_0_0,
  input  [6:0]   io_key_config_1_field_id_0_1,
  input  [6:0]   io_key_config_1_field_id_0_2,
  input  [6:0]   io_key_config_1_field_id_0_3,
  input  [6:0]   io_key_config_1_field_id_1_0,
  input  [6:0]   io_key_config_1_field_id_1_1,
  input  [6:0]   io_key_config_1_field_id_1_2,
  input  [6:0]   io_key_config_1_field_id_1_3,
  input  [6:0]   io_key_config_1_field_id_2_0,
  input  [6:0]   io_key_config_1_field_id_2_1,
  input  [6:0]   io_key_config_1_field_id_2_2,
  input  [6:0]   io_key_config_1_field_id_2_3,
  input  [6:0]   io_key_config_1_field_id_3_0,
  input  [6:0]   io_key_config_1_field_id_3_1,
  input  [6:0]   io_key_config_1_field_id_3_2,
  input  [6:0]   io_key_config_1_field_id_3_3,
  input  [6:0]   io_key_config_1_field_id_4_0,
  input  [6:0]   io_key_config_1_field_id_4_1,
  input  [6:0]   io_key_config_1_field_id_4_2,
  input  [6:0]   io_key_config_1_field_id_4_3,
  input  [6:0]   io_key_config_1_field_id_5_0,
  input  [6:0]   io_key_config_1_field_id_5_1,
  input  [6:0]   io_key_config_1_field_id_5_2,
  input  [6:0]   io_key_config_1_field_id_5_3,
  output [191:0] io_match_key
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_1; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_2; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_3; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_4; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_5; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_6; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_7; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_8; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_9; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_10; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_11; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_12; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_13; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_14; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_15; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_16; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_17; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_18; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_19; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_20; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_21; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_22; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_23; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_24; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_25; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_26; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_27; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_28; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_29; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_30; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_31; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_32; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_33; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_34; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_35; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_36; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_37; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_38; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_39; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_40; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_41; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_42; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_43; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_44; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_45; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_46; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_47; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_48; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_49; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_50; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_51; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_52; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_53; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_54; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_55; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_56; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_57; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_58; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_59; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_60; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_61; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_62; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_63; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_64; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_65; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_66; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_67; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_68; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_69; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_70; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_71; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_72; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_73; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_74; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_75; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_76; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_77; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_78; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_79; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_80; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_81; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_82; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_83; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_84; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_85; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_86; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_87; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_88; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_89; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_90; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_91; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_92; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_93; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_94; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_95; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_96; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_97; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_98; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_99; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_100; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_101; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_102; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_103; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_104; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_105; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_106; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_107; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_108; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_109; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_110; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_111; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_112; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_113; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_114; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_115; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_116; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_117; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_118; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_119; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_120; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_121; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_122; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_123; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_124; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_125; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_126; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_127; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_128; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_129; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_130; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_131; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_132; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_133; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_134; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_135; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_136; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_137; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_138; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_139; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_140; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_141; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_142; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_143; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_144; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_145; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_146; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_147; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_148; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_149; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_150; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_151; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_152; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_153; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_154; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_155; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_156; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_157; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_158; // @[matcher_pisa.scala 102:22]
  reg [7:0] phv_data_159; // @[matcher_pisa.scala 102:22]
  reg  phv_next_config_id; // @[matcher_pisa.scala 102:22]
  reg  phv_is_valid_processor; // @[matcher_pisa.scala 102:22]
  wire [1:0] _GEN_56 = phv_next_config_id ? io_key_config_1_field_config_0 : io_key_config_0_field_config_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [1:0] _GEN_57 = phv_next_config_id ? io_key_config_1_field_config_1 : io_key_config_0_field_config_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [1:0] _GEN_58 = phv_next_config_id ? io_key_config_1_field_config_2 : io_key_config_0_field_config_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [1:0] _GEN_59 = phv_next_config_id ? io_key_config_1_field_config_3 : io_key_config_0_field_config_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [1:0] _GEN_60 = phv_next_config_id ? io_key_config_1_field_config_4 : io_key_config_0_field_config_4; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [1:0] _GEN_61 = phv_next_config_id ? io_key_config_1_field_config_5 : io_key_config_0_field_config_5; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_62 = phv_next_config_id ? io_key_config_1_field_mask_0_0 : io_key_config_0_field_mask_0_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_63 = phv_next_config_id ? io_key_config_1_field_mask_0_1 : io_key_config_0_field_mask_0_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_64 = phv_next_config_id ? io_key_config_1_field_mask_0_2 : io_key_config_0_field_mask_0_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_65 = phv_next_config_id ? io_key_config_1_field_mask_0_3 : io_key_config_0_field_mask_0_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_66 = phv_next_config_id ? io_key_config_1_field_mask_1_0 : io_key_config_0_field_mask_1_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_67 = phv_next_config_id ? io_key_config_1_field_mask_1_1 : io_key_config_0_field_mask_1_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_68 = phv_next_config_id ? io_key_config_1_field_mask_1_2 : io_key_config_0_field_mask_1_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_69 = phv_next_config_id ? io_key_config_1_field_mask_1_3 : io_key_config_0_field_mask_1_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_70 = phv_next_config_id ? io_key_config_1_field_mask_2_0 : io_key_config_0_field_mask_2_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_71 = phv_next_config_id ? io_key_config_1_field_mask_2_1 : io_key_config_0_field_mask_2_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_72 = phv_next_config_id ? io_key_config_1_field_mask_2_2 : io_key_config_0_field_mask_2_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_73 = phv_next_config_id ? io_key_config_1_field_mask_2_3 : io_key_config_0_field_mask_2_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_74 = phv_next_config_id ? io_key_config_1_field_mask_3_0 : io_key_config_0_field_mask_3_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_75 = phv_next_config_id ? io_key_config_1_field_mask_3_1 : io_key_config_0_field_mask_3_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_76 = phv_next_config_id ? io_key_config_1_field_mask_3_2 : io_key_config_0_field_mask_3_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_77 = phv_next_config_id ? io_key_config_1_field_mask_3_3 : io_key_config_0_field_mask_3_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_78 = phv_next_config_id ? io_key_config_1_field_mask_4_0 : io_key_config_0_field_mask_4_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_79 = phv_next_config_id ? io_key_config_1_field_mask_4_1 : io_key_config_0_field_mask_4_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_80 = phv_next_config_id ? io_key_config_1_field_mask_4_2 : io_key_config_0_field_mask_4_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_81 = phv_next_config_id ? io_key_config_1_field_mask_4_3 : io_key_config_0_field_mask_4_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_82 = phv_next_config_id ? io_key_config_1_field_mask_5_0 : io_key_config_0_field_mask_5_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_83 = phv_next_config_id ? io_key_config_1_field_mask_5_1 : io_key_config_0_field_mask_5_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_84 = phv_next_config_id ? io_key_config_1_field_mask_5_2 : io_key_config_0_field_mask_5_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire  _GEN_85 = phv_next_config_id ? io_key_config_1_field_mask_5_3 : io_key_config_0_field_mask_5_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_86 = phv_next_config_id ? io_key_config_1_field_id_0_0 : io_key_config_0_field_id_0_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_87 = phv_next_config_id ? io_key_config_1_field_id_0_1 : io_key_config_0_field_id_0_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_88 = phv_next_config_id ? io_key_config_1_field_id_0_2 : io_key_config_0_field_id_0_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_89 = phv_next_config_id ? io_key_config_1_field_id_0_3 : io_key_config_0_field_id_0_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_90 = phv_next_config_id ? io_key_config_1_field_id_1_0 : io_key_config_0_field_id_1_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_91 = phv_next_config_id ? io_key_config_1_field_id_1_1 : io_key_config_0_field_id_1_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_92 = phv_next_config_id ? io_key_config_1_field_id_1_2 : io_key_config_0_field_id_1_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_93 = phv_next_config_id ? io_key_config_1_field_id_1_3 : io_key_config_0_field_id_1_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_94 = phv_next_config_id ? io_key_config_1_field_id_2_0 : io_key_config_0_field_id_2_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_95 = phv_next_config_id ? io_key_config_1_field_id_2_1 : io_key_config_0_field_id_2_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_96 = phv_next_config_id ? io_key_config_1_field_id_2_2 : io_key_config_0_field_id_2_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_97 = phv_next_config_id ? io_key_config_1_field_id_2_3 : io_key_config_0_field_id_2_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_98 = phv_next_config_id ? io_key_config_1_field_id_3_0 : io_key_config_0_field_id_3_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_99 = phv_next_config_id ? io_key_config_1_field_id_3_1 : io_key_config_0_field_id_3_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_100 = phv_next_config_id ? io_key_config_1_field_id_3_2 : io_key_config_0_field_id_3_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_101 = phv_next_config_id ? io_key_config_1_field_id_3_3 : io_key_config_0_field_id_3_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_102 = phv_next_config_id ? io_key_config_1_field_id_4_0 : io_key_config_0_field_id_4_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_103 = phv_next_config_id ? io_key_config_1_field_id_4_1 : io_key_config_0_field_id_4_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_104 = phv_next_config_id ? io_key_config_1_field_id_4_2 : io_key_config_0_field_id_4_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_105 = phv_next_config_id ? io_key_config_1_field_id_4_3 : io_key_config_0_field_id_4_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_106 = phv_next_config_id ? io_key_config_1_field_id_5_0 : io_key_config_0_field_id_5_0; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_107 = phv_next_config_id ? io_key_config_1_field_id_5_1 : io_key_config_0_field_id_5_1; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_108 = phv_next_config_id ? io_key_config_1_field_id_5_2 : io_key_config_0_field_id_5_2; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [6:0] _GEN_109 = phv_next_config_id ? io_key_config_1_field_id_5_3 : io_key_config_0_field_id_5_3; // @[matcher_pisa.scala 115:36 matcher_pisa.scala 115:36]
  wire [7:0] _GEN_110 = 7'h0 == _GEN_86 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_111 = 7'h1 == _GEN_86 ? phv_data_1 : _GEN_110; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_112 = 7'h2 == _GEN_86 ? phv_data_2 : _GEN_111; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_113 = 7'h3 == _GEN_86 ? phv_data_3 : _GEN_112; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_114 = 7'h4 == _GEN_86 ? phv_data_4 : _GEN_113; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_115 = 7'h5 == _GEN_86 ? phv_data_5 : _GEN_114; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_116 = 7'h6 == _GEN_86 ? phv_data_6 : _GEN_115; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_117 = 7'h7 == _GEN_86 ? phv_data_7 : _GEN_116; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_118 = 7'h8 == _GEN_86 ? phv_data_8 : _GEN_117; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_119 = 7'h9 == _GEN_86 ? phv_data_9 : _GEN_118; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_120 = 7'ha == _GEN_86 ? phv_data_10 : _GEN_119; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_121 = 7'hb == _GEN_86 ? phv_data_11 : _GEN_120; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_122 = 7'hc == _GEN_86 ? phv_data_12 : _GEN_121; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_123 = 7'hd == _GEN_86 ? phv_data_13 : _GEN_122; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_124 = 7'he == _GEN_86 ? phv_data_14 : _GEN_123; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_125 = 7'hf == _GEN_86 ? phv_data_15 : _GEN_124; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_126 = 7'h10 == _GEN_86 ? phv_data_16 : _GEN_125; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_127 = 7'h11 == _GEN_86 ? phv_data_17 : _GEN_126; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_128 = 7'h12 == _GEN_86 ? phv_data_18 : _GEN_127; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_129 = 7'h13 == _GEN_86 ? phv_data_19 : _GEN_128; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes__0 = _GEN_62 ? _GEN_129 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_131 = 7'h0 == _GEN_87 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_132 = 7'h1 == _GEN_87 ? phv_data_1 : _GEN_131; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_133 = 7'h2 == _GEN_87 ? phv_data_2 : _GEN_132; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_134 = 7'h3 == _GEN_87 ? phv_data_3 : _GEN_133; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_135 = 7'h4 == _GEN_87 ? phv_data_4 : _GEN_134; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_136 = 7'h5 == _GEN_87 ? phv_data_5 : _GEN_135; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_137 = 7'h6 == _GEN_87 ? phv_data_6 : _GEN_136; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_138 = 7'h7 == _GEN_87 ? phv_data_7 : _GEN_137; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_139 = 7'h8 == _GEN_87 ? phv_data_8 : _GEN_138; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_140 = 7'h9 == _GEN_87 ? phv_data_9 : _GEN_139; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_141 = 7'ha == _GEN_87 ? phv_data_10 : _GEN_140; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_142 = 7'hb == _GEN_87 ? phv_data_11 : _GEN_141; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_143 = 7'hc == _GEN_87 ? phv_data_12 : _GEN_142; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_144 = 7'hd == _GEN_87 ? phv_data_13 : _GEN_143; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_145 = 7'he == _GEN_87 ? phv_data_14 : _GEN_144; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_146 = 7'hf == _GEN_87 ? phv_data_15 : _GEN_145; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_147 = 7'h10 == _GEN_87 ? phv_data_16 : _GEN_146; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_148 = 7'h11 == _GEN_87 ? phv_data_17 : _GEN_147; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_149 = 7'h12 == _GEN_87 ? phv_data_18 : _GEN_148; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_150 = 7'h13 == _GEN_87 ? phv_data_19 : _GEN_149; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes__1 = _GEN_63 ? _GEN_150 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_152 = 7'h0 == _GEN_88 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_153 = 7'h1 == _GEN_88 ? phv_data_1 : _GEN_152; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_154 = 7'h2 == _GEN_88 ? phv_data_2 : _GEN_153; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_155 = 7'h3 == _GEN_88 ? phv_data_3 : _GEN_154; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_156 = 7'h4 == _GEN_88 ? phv_data_4 : _GEN_155; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_157 = 7'h5 == _GEN_88 ? phv_data_5 : _GEN_156; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_158 = 7'h6 == _GEN_88 ? phv_data_6 : _GEN_157; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_159 = 7'h7 == _GEN_88 ? phv_data_7 : _GEN_158; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_160 = 7'h8 == _GEN_88 ? phv_data_8 : _GEN_159; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_161 = 7'h9 == _GEN_88 ? phv_data_9 : _GEN_160; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_162 = 7'ha == _GEN_88 ? phv_data_10 : _GEN_161; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_163 = 7'hb == _GEN_88 ? phv_data_11 : _GEN_162; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_164 = 7'hc == _GEN_88 ? phv_data_12 : _GEN_163; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_165 = 7'hd == _GEN_88 ? phv_data_13 : _GEN_164; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_166 = 7'he == _GEN_88 ? phv_data_14 : _GEN_165; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_167 = 7'hf == _GEN_88 ? phv_data_15 : _GEN_166; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_168 = 7'h10 == _GEN_88 ? phv_data_16 : _GEN_167; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_169 = 7'h11 == _GEN_88 ? phv_data_17 : _GEN_168; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_170 = 7'h12 == _GEN_88 ? phv_data_18 : _GEN_169; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_171 = 7'h13 == _GEN_88 ? phv_data_19 : _GEN_170; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes__2 = _GEN_64 ? _GEN_171 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_173 = 7'h0 == _GEN_89 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_174 = 7'h1 == _GEN_89 ? phv_data_1 : _GEN_173; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_175 = 7'h2 == _GEN_89 ? phv_data_2 : _GEN_174; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_176 = 7'h3 == _GEN_89 ? phv_data_3 : _GEN_175; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_177 = 7'h4 == _GEN_89 ? phv_data_4 : _GEN_176; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_178 = 7'h5 == _GEN_89 ? phv_data_5 : _GEN_177; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_179 = 7'h6 == _GEN_89 ? phv_data_6 : _GEN_178; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_180 = 7'h7 == _GEN_89 ? phv_data_7 : _GEN_179; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_181 = 7'h8 == _GEN_89 ? phv_data_8 : _GEN_180; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_182 = 7'h9 == _GEN_89 ? phv_data_9 : _GEN_181; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_183 = 7'ha == _GEN_89 ? phv_data_10 : _GEN_182; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_184 = 7'hb == _GEN_89 ? phv_data_11 : _GEN_183; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_185 = 7'hc == _GEN_89 ? phv_data_12 : _GEN_184; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_186 = 7'hd == _GEN_89 ? phv_data_13 : _GEN_185; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_187 = 7'he == _GEN_89 ? phv_data_14 : _GEN_186; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_188 = 7'hf == _GEN_89 ? phv_data_15 : _GEN_187; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_189 = 7'h10 == _GEN_89 ? phv_data_16 : _GEN_188; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_190 = 7'h11 == _GEN_89 ? phv_data_17 : _GEN_189; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_191 = 7'h12 == _GEN_89 ? phv_data_18 : _GEN_190; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_192 = 7'h13 == _GEN_89 ? phv_data_19 : _GEN_191; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes__3 = _GEN_65 ? _GEN_192 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [31:0] _groups_0_T = {bytes__0,bytes__1,bytes__2,bytes__3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_194 = _GEN_56 == 2'h1 ? _groups_0_T : 32'h0; // @[matcher_pisa.scala 115:50 matcher_pisa.scala 129:31 matcher_pisa.scala 114:27]
  wire [15:0] _double_bytes_0_T = {phv_data_20,phv_data_21}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_195 = 7'h14 == _GEN_86 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _double_bytes_0_T_1 = {phv_data_22,phv_data_23}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_196 = 7'h15 == _GEN_86 ? _double_bytes_0_T_1 : _GEN_195; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_2 = {phv_data_24,phv_data_25}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_197 = 7'h16 == _GEN_86 ? _double_bytes_0_T_2 : _GEN_196; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_3 = {phv_data_26,phv_data_27}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_198 = 7'h17 == _GEN_86 ? _double_bytes_0_T_3 : _GEN_197; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_4 = {phv_data_28,phv_data_29}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_199 = 7'h18 == _GEN_86 ? _double_bytes_0_T_4 : _GEN_198; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_5 = {phv_data_30,phv_data_31}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_200 = 7'h19 == _GEN_86 ? _double_bytes_0_T_5 : _GEN_199; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_6 = {phv_data_32,phv_data_33}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_201 = 7'h1a == _GEN_86 ? _double_bytes_0_T_6 : _GEN_200; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_7 = {phv_data_34,phv_data_35}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_202 = 7'h1b == _GEN_86 ? _double_bytes_0_T_7 : _GEN_201; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_8 = {phv_data_36,phv_data_37}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_203 = 7'h1c == _GEN_86 ? _double_bytes_0_T_8 : _GEN_202; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_9 = {phv_data_38,phv_data_39}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_204 = 7'h1d == _GEN_86 ? _double_bytes_0_T_9 : _GEN_203; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_10 = {phv_data_40,phv_data_41}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_205 = 7'h1e == _GEN_86 ? _double_bytes_0_T_10 : _GEN_204; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_11 = {phv_data_42,phv_data_43}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_206 = 7'h1f == _GEN_86 ? _double_bytes_0_T_11 : _GEN_205; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_12 = {phv_data_44,phv_data_45}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_207 = 7'h20 == _GEN_86 ? _double_bytes_0_T_12 : _GEN_206; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_13 = {phv_data_46,phv_data_47}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_208 = 7'h21 == _GEN_86 ? _double_bytes_0_T_13 : _GEN_207; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_14 = {phv_data_48,phv_data_49}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_209 = 7'h22 == _GEN_86 ? _double_bytes_0_T_14 : _GEN_208; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_15 = {phv_data_50,phv_data_51}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_210 = 7'h23 == _GEN_86 ? _double_bytes_0_T_15 : _GEN_209; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_16 = {phv_data_52,phv_data_53}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_211 = 7'h24 == _GEN_86 ? _double_bytes_0_T_16 : _GEN_210; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_17 = {phv_data_54,phv_data_55}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_212 = 7'h25 == _GEN_86 ? _double_bytes_0_T_17 : _GEN_211; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_18 = {phv_data_56,phv_data_57}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_213 = 7'h26 == _GEN_86 ? _double_bytes_0_T_18 : _GEN_212; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_19 = {phv_data_58,phv_data_59}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_214 = 7'h27 == _GEN_86 ? _double_bytes_0_T_19 : _GEN_213; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_20 = {phv_data_60,phv_data_61}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_215 = 7'h28 == _GEN_86 ? _double_bytes_0_T_20 : _GEN_214; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_21 = {phv_data_62,phv_data_63}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_216 = 7'h29 == _GEN_86 ? _double_bytes_0_T_21 : _GEN_215; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_22 = {phv_data_64,phv_data_65}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_217 = 7'h2a == _GEN_86 ? _double_bytes_0_T_22 : _GEN_216; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_23 = {phv_data_66,phv_data_67}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_218 = 7'h2b == _GEN_86 ? _double_bytes_0_T_23 : _GEN_217; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_24 = {phv_data_68,phv_data_69}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_219 = 7'h2c == _GEN_86 ? _double_bytes_0_T_24 : _GEN_218; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_25 = {phv_data_70,phv_data_71}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_220 = 7'h2d == _GEN_86 ? _double_bytes_0_T_25 : _GEN_219; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_26 = {phv_data_72,phv_data_73}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_221 = 7'h2e == _GEN_86 ? _double_bytes_0_T_26 : _GEN_220; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_27 = {phv_data_74,phv_data_75}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_222 = 7'h2f == _GEN_86 ? _double_bytes_0_T_27 : _GEN_221; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_28 = {phv_data_76,phv_data_77}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_223 = 7'h30 == _GEN_86 ? _double_bytes_0_T_28 : _GEN_222; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _double_bytes_0_T_29 = {phv_data_78,phv_data_79}; // @[Cat.scala 30:58]
  wire [15:0] _GEN_224 = 7'h31 == _GEN_86 ? _double_bytes_0_T_29 : _GEN_223; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes__0 = _GEN_62 ? _GEN_224 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_226 = 7'h14 == _GEN_87 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_227 = 7'h15 == _GEN_87 ? _double_bytes_0_T_1 : _GEN_226; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_228 = 7'h16 == _GEN_87 ? _double_bytes_0_T_2 : _GEN_227; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_229 = 7'h17 == _GEN_87 ? _double_bytes_0_T_3 : _GEN_228; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_230 = 7'h18 == _GEN_87 ? _double_bytes_0_T_4 : _GEN_229; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_231 = 7'h19 == _GEN_87 ? _double_bytes_0_T_5 : _GEN_230; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_232 = 7'h1a == _GEN_87 ? _double_bytes_0_T_6 : _GEN_231; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_233 = 7'h1b == _GEN_87 ? _double_bytes_0_T_7 : _GEN_232; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_234 = 7'h1c == _GEN_87 ? _double_bytes_0_T_8 : _GEN_233; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_235 = 7'h1d == _GEN_87 ? _double_bytes_0_T_9 : _GEN_234; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_236 = 7'h1e == _GEN_87 ? _double_bytes_0_T_10 : _GEN_235; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_237 = 7'h1f == _GEN_87 ? _double_bytes_0_T_11 : _GEN_236; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_238 = 7'h20 == _GEN_87 ? _double_bytes_0_T_12 : _GEN_237; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_239 = 7'h21 == _GEN_87 ? _double_bytes_0_T_13 : _GEN_238; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_240 = 7'h22 == _GEN_87 ? _double_bytes_0_T_14 : _GEN_239; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_241 = 7'h23 == _GEN_87 ? _double_bytes_0_T_15 : _GEN_240; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_242 = 7'h24 == _GEN_87 ? _double_bytes_0_T_16 : _GEN_241; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_243 = 7'h25 == _GEN_87 ? _double_bytes_0_T_17 : _GEN_242; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_244 = 7'h26 == _GEN_87 ? _double_bytes_0_T_18 : _GEN_243; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_245 = 7'h27 == _GEN_87 ? _double_bytes_0_T_19 : _GEN_244; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_246 = 7'h28 == _GEN_87 ? _double_bytes_0_T_20 : _GEN_245; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_247 = 7'h29 == _GEN_87 ? _double_bytes_0_T_21 : _GEN_246; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_248 = 7'h2a == _GEN_87 ? _double_bytes_0_T_22 : _GEN_247; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_249 = 7'h2b == _GEN_87 ? _double_bytes_0_T_23 : _GEN_248; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_250 = 7'h2c == _GEN_87 ? _double_bytes_0_T_24 : _GEN_249; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_251 = 7'h2d == _GEN_87 ? _double_bytes_0_T_25 : _GEN_250; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_252 = 7'h2e == _GEN_87 ? _double_bytes_0_T_26 : _GEN_251; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_253 = 7'h2f == _GEN_87 ? _double_bytes_0_T_27 : _GEN_252; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_254 = 7'h30 == _GEN_87 ? _double_bytes_0_T_28 : _GEN_253; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_255 = 7'h31 == _GEN_87 ? _double_bytes_0_T_29 : _GEN_254; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes__1 = _GEN_63 ? _GEN_255 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [31:0] _groups_0_T_1 = {double_bytes__0,double_bytes__1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_257 = _GEN_56 == 2'h2 ? _groups_0_T_1 : _GEN_194; // @[matcher_pisa.scala 131:50 matcher_pisa.scala 145:31]
  wire [31:0] _groups_0_T_2 = {phv_data_80,phv_data_81,phv_data_82,phv_data_83}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_258 = 7'h32 == _GEN_86 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39 matcher_pisa.scala 150:31]
  wire [31:0] _groups_0_T_3 = {phv_data_84,phv_data_85,phv_data_86,phv_data_87}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_259 = 7'h33 == _GEN_86 ? _groups_0_T_3 : _GEN_258; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_4 = {phv_data_88,phv_data_89,phv_data_90,phv_data_91}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_260 = 7'h34 == _GEN_86 ? _groups_0_T_4 : _GEN_259; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_5 = {phv_data_92,phv_data_93,phv_data_94,phv_data_95}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_261 = 7'h35 == _GEN_86 ? _groups_0_T_5 : _GEN_260; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_6 = {phv_data_96,phv_data_97,phv_data_98,phv_data_99}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_262 = 7'h36 == _GEN_86 ? _groups_0_T_6 : _GEN_261; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_7 = {phv_data_100,phv_data_101,phv_data_102,phv_data_103}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_263 = 7'h37 == _GEN_86 ? _groups_0_T_7 : _GEN_262; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_8 = {phv_data_104,phv_data_105,phv_data_106,phv_data_107}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_264 = 7'h38 == _GEN_86 ? _groups_0_T_8 : _GEN_263; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_9 = {phv_data_108,phv_data_109,phv_data_110,phv_data_111}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_265 = 7'h39 == _GEN_86 ? _groups_0_T_9 : _GEN_264; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_10 = {phv_data_112,phv_data_113,phv_data_114,phv_data_115}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_266 = 7'h3a == _GEN_86 ? _groups_0_T_10 : _GEN_265; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_11 = {phv_data_116,phv_data_117,phv_data_118,phv_data_119}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_267 = 7'h3b == _GEN_86 ? _groups_0_T_11 : _GEN_266; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_12 = {phv_data_120,phv_data_121,phv_data_122,phv_data_123}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_268 = 7'h3c == _GEN_86 ? _groups_0_T_12 : _GEN_267; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_13 = {phv_data_124,phv_data_125,phv_data_126,phv_data_127}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_269 = 7'h3d == _GEN_86 ? _groups_0_T_13 : _GEN_268; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_14 = {phv_data_128,phv_data_129,phv_data_130,phv_data_131}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_270 = 7'h3e == _GEN_86 ? _groups_0_T_14 : _GEN_269; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_15 = {phv_data_132,phv_data_133,phv_data_134,phv_data_135}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_271 = 7'h3f == _GEN_86 ? _groups_0_T_15 : _GEN_270; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_16 = {phv_data_136,phv_data_137,phv_data_138,phv_data_139}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_272 = 7'h40 == _GEN_86 ? _groups_0_T_16 : _GEN_271; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_17 = {phv_data_140,phv_data_141,phv_data_142,phv_data_143}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_273 = 7'h41 == _GEN_86 ? _groups_0_T_17 : _GEN_272; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_18 = {phv_data_144,phv_data_145,phv_data_146,phv_data_147}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_274 = 7'h42 == _GEN_86 ? _groups_0_T_18 : _GEN_273; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_19 = {phv_data_148,phv_data_149,phv_data_150,phv_data_151}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_275 = 7'h43 == _GEN_86 ? _groups_0_T_19 : _GEN_274; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_20 = {phv_data_152,phv_data_153,phv_data_154,phv_data_155}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_276 = 7'h44 == _GEN_86 ? _groups_0_T_20 : _GEN_275; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _groups_0_T_21 = {phv_data_156,phv_data_157,phv_data_158,phv_data_159}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_277 = 7'h45 == _GEN_86 ? _groups_0_T_21 : _GEN_276; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] groups_0 = _GEN_56 == 2'h3 ? _GEN_277 : _GEN_257; // @[matcher_pisa.scala 147:50]
  wire [7:0] _GEN_279 = 7'h0 == _GEN_90 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_280 = 7'h1 == _GEN_90 ? phv_data_1 : _GEN_279; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_281 = 7'h2 == _GEN_90 ? phv_data_2 : _GEN_280; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_282 = 7'h3 == _GEN_90 ? phv_data_3 : _GEN_281; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_283 = 7'h4 == _GEN_90 ? phv_data_4 : _GEN_282; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_284 = 7'h5 == _GEN_90 ? phv_data_5 : _GEN_283; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_285 = 7'h6 == _GEN_90 ? phv_data_6 : _GEN_284; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_286 = 7'h7 == _GEN_90 ? phv_data_7 : _GEN_285; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_287 = 7'h8 == _GEN_90 ? phv_data_8 : _GEN_286; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_288 = 7'h9 == _GEN_90 ? phv_data_9 : _GEN_287; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_289 = 7'ha == _GEN_90 ? phv_data_10 : _GEN_288; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_290 = 7'hb == _GEN_90 ? phv_data_11 : _GEN_289; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_291 = 7'hc == _GEN_90 ? phv_data_12 : _GEN_290; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_292 = 7'hd == _GEN_90 ? phv_data_13 : _GEN_291; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_293 = 7'he == _GEN_90 ? phv_data_14 : _GEN_292; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_294 = 7'hf == _GEN_90 ? phv_data_15 : _GEN_293; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_295 = 7'h10 == _GEN_90 ? phv_data_16 : _GEN_294; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_296 = 7'h11 == _GEN_90 ? phv_data_17 : _GEN_295; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_297 = 7'h12 == _GEN_90 ? phv_data_18 : _GEN_296; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_298 = 7'h13 == _GEN_90 ? phv_data_19 : _GEN_297; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_1_0 = _GEN_66 ? _GEN_298 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_300 = 7'h0 == _GEN_91 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_301 = 7'h1 == _GEN_91 ? phv_data_1 : _GEN_300; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_302 = 7'h2 == _GEN_91 ? phv_data_2 : _GEN_301; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_303 = 7'h3 == _GEN_91 ? phv_data_3 : _GEN_302; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_304 = 7'h4 == _GEN_91 ? phv_data_4 : _GEN_303; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_305 = 7'h5 == _GEN_91 ? phv_data_5 : _GEN_304; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_306 = 7'h6 == _GEN_91 ? phv_data_6 : _GEN_305; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_307 = 7'h7 == _GEN_91 ? phv_data_7 : _GEN_306; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_308 = 7'h8 == _GEN_91 ? phv_data_8 : _GEN_307; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_309 = 7'h9 == _GEN_91 ? phv_data_9 : _GEN_308; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_310 = 7'ha == _GEN_91 ? phv_data_10 : _GEN_309; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_311 = 7'hb == _GEN_91 ? phv_data_11 : _GEN_310; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_312 = 7'hc == _GEN_91 ? phv_data_12 : _GEN_311; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_313 = 7'hd == _GEN_91 ? phv_data_13 : _GEN_312; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_314 = 7'he == _GEN_91 ? phv_data_14 : _GEN_313; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_315 = 7'hf == _GEN_91 ? phv_data_15 : _GEN_314; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_316 = 7'h10 == _GEN_91 ? phv_data_16 : _GEN_315; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_317 = 7'h11 == _GEN_91 ? phv_data_17 : _GEN_316; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_318 = 7'h12 == _GEN_91 ? phv_data_18 : _GEN_317; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_319 = 7'h13 == _GEN_91 ? phv_data_19 : _GEN_318; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_1_1 = _GEN_67 ? _GEN_319 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_321 = 7'h0 == _GEN_92 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_322 = 7'h1 == _GEN_92 ? phv_data_1 : _GEN_321; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_323 = 7'h2 == _GEN_92 ? phv_data_2 : _GEN_322; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_324 = 7'h3 == _GEN_92 ? phv_data_3 : _GEN_323; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_325 = 7'h4 == _GEN_92 ? phv_data_4 : _GEN_324; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_326 = 7'h5 == _GEN_92 ? phv_data_5 : _GEN_325; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_327 = 7'h6 == _GEN_92 ? phv_data_6 : _GEN_326; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_328 = 7'h7 == _GEN_92 ? phv_data_7 : _GEN_327; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_329 = 7'h8 == _GEN_92 ? phv_data_8 : _GEN_328; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_330 = 7'h9 == _GEN_92 ? phv_data_9 : _GEN_329; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_331 = 7'ha == _GEN_92 ? phv_data_10 : _GEN_330; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_332 = 7'hb == _GEN_92 ? phv_data_11 : _GEN_331; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_333 = 7'hc == _GEN_92 ? phv_data_12 : _GEN_332; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_334 = 7'hd == _GEN_92 ? phv_data_13 : _GEN_333; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_335 = 7'he == _GEN_92 ? phv_data_14 : _GEN_334; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_336 = 7'hf == _GEN_92 ? phv_data_15 : _GEN_335; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_337 = 7'h10 == _GEN_92 ? phv_data_16 : _GEN_336; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_338 = 7'h11 == _GEN_92 ? phv_data_17 : _GEN_337; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_339 = 7'h12 == _GEN_92 ? phv_data_18 : _GEN_338; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_340 = 7'h13 == _GEN_92 ? phv_data_19 : _GEN_339; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_1_2 = _GEN_68 ? _GEN_340 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_342 = 7'h0 == _GEN_93 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_343 = 7'h1 == _GEN_93 ? phv_data_1 : _GEN_342; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_344 = 7'h2 == _GEN_93 ? phv_data_2 : _GEN_343; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_345 = 7'h3 == _GEN_93 ? phv_data_3 : _GEN_344; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_346 = 7'h4 == _GEN_93 ? phv_data_4 : _GEN_345; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_347 = 7'h5 == _GEN_93 ? phv_data_5 : _GEN_346; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_348 = 7'h6 == _GEN_93 ? phv_data_6 : _GEN_347; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_349 = 7'h7 == _GEN_93 ? phv_data_7 : _GEN_348; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_350 = 7'h8 == _GEN_93 ? phv_data_8 : _GEN_349; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_351 = 7'h9 == _GEN_93 ? phv_data_9 : _GEN_350; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_352 = 7'ha == _GEN_93 ? phv_data_10 : _GEN_351; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_353 = 7'hb == _GEN_93 ? phv_data_11 : _GEN_352; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_354 = 7'hc == _GEN_93 ? phv_data_12 : _GEN_353; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_355 = 7'hd == _GEN_93 ? phv_data_13 : _GEN_354; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_356 = 7'he == _GEN_93 ? phv_data_14 : _GEN_355; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_357 = 7'hf == _GEN_93 ? phv_data_15 : _GEN_356; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_358 = 7'h10 == _GEN_93 ? phv_data_16 : _GEN_357; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_359 = 7'h11 == _GEN_93 ? phv_data_17 : _GEN_358; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_360 = 7'h12 == _GEN_93 ? phv_data_18 : _GEN_359; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_361 = 7'h13 == _GEN_93 ? phv_data_19 : _GEN_360; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_1_3 = _GEN_69 ? _GEN_361 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [31:0] _groups_1_T = {bytes_1_0,bytes_1_1,bytes_1_2,bytes_1_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_363 = _GEN_57 == 2'h1 ? _groups_1_T : 32'h0; // @[matcher_pisa.scala 115:50 matcher_pisa.scala 129:31 matcher_pisa.scala 114:27]
  wire [15:0] _GEN_364 = 7'h14 == _GEN_90 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_365 = 7'h15 == _GEN_90 ? _double_bytes_0_T_1 : _GEN_364; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_366 = 7'h16 == _GEN_90 ? _double_bytes_0_T_2 : _GEN_365; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_367 = 7'h17 == _GEN_90 ? _double_bytes_0_T_3 : _GEN_366; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_368 = 7'h18 == _GEN_90 ? _double_bytes_0_T_4 : _GEN_367; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_369 = 7'h19 == _GEN_90 ? _double_bytes_0_T_5 : _GEN_368; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_370 = 7'h1a == _GEN_90 ? _double_bytes_0_T_6 : _GEN_369; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_371 = 7'h1b == _GEN_90 ? _double_bytes_0_T_7 : _GEN_370; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_372 = 7'h1c == _GEN_90 ? _double_bytes_0_T_8 : _GEN_371; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_373 = 7'h1d == _GEN_90 ? _double_bytes_0_T_9 : _GEN_372; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_374 = 7'h1e == _GEN_90 ? _double_bytes_0_T_10 : _GEN_373; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_375 = 7'h1f == _GEN_90 ? _double_bytes_0_T_11 : _GEN_374; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_376 = 7'h20 == _GEN_90 ? _double_bytes_0_T_12 : _GEN_375; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_377 = 7'h21 == _GEN_90 ? _double_bytes_0_T_13 : _GEN_376; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_378 = 7'h22 == _GEN_90 ? _double_bytes_0_T_14 : _GEN_377; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_379 = 7'h23 == _GEN_90 ? _double_bytes_0_T_15 : _GEN_378; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_380 = 7'h24 == _GEN_90 ? _double_bytes_0_T_16 : _GEN_379; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_381 = 7'h25 == _GEN_90 ? _double_bytes_0_T_17 : _GEN_380; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_382 = 7'h26 == _GEN_90 ? _double_bytes_0_T_18 : _GEN_381; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_383 = 7'h27 == _GEN_90 ? _double_bytes_0_T_19 : _GEN_382; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_384 = 7'h28 == _GEN_90 ? _double_bytes_0_T_20 : _GEN_383; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_385 = 7'h29 == _GEN_90 ? _double_bytes_0_T_21 : _GEN_384; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_386 = 7'h2a == _GEN_90 ? _double_bytes_0_T_22 : _GEN_385; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_387 = 7'h2b == _GEN_90 ? _double_bytes_0_T_23 : _GEN_386; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_388 = 7'h2c == _GEN_90 ? _double_bytes_0_T_24 : _GEN_387; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_389 = 7'h2d == _GEN_90 ? _double_bytes_0_T_25 : _GEN_388; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_390 = 7'h2e == _GEN_90 ? _double_bytes_0_T_26 : _GEN_389; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_391 = 7'h2f == _GEN_90 ? _double_bytes_0_T_27 : _GEN_390; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_392 = 7'h30 == _GEN_90 ? _double_bytes_0_T_28 : _GEN_391; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_393 = 7'h31 == _GEN_90 ? _double_bytes_0_T_29 : _GEN_392; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_1_0 = _GEN_66 ? _GEN_393 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_395 = 7'h14 == _GEN_91 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_396 = 7'h15 == _GEN_91 ? _double_bytes_0_T_1 : _GEN_395; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_397 = 7'h16 == _GEN_91 ? _double_bytes_0_T_2 : _GEN_396; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_398 = 7'h17 == _GEN_91 ? _double_bytes_0_T_3 : _GEN_397; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_399 = 7'h18 == _GEN_91 ? _double_bytes_0_T_4 : _GEN_398; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_400 = 7'h19 == _GEN_91 ? _double_bytes_0_T_5 : _GEN_399; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_401 = 7'h1a == _GEN_91 ? _double_bytes_0_T_6 : _GEN_400; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_402 = 7'h1b == _GEN_91 ? _double_bytes_0_T_7 : _GEN_401; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_403 = 7'h1c == _GEN_91 ? _double_bytes_0_T_8 : _GEN_402; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_404 = 7'h1d == _GEN_91 ? _double_bytes_0_T_9 : _GEN_403; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_405 = 7'h1e == _GEN_91 ? _double_bytes_0_T_10 : _GEN_404; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_406 = 7'h1f == _GEN_91 ? _double_bytes_0_T_11 : _GEN_405; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_407 = 7'h20 == _GEN_91 ? _double_bytes_0_T_12 : _GEN_406; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_408 = 7'h21 == _GEN_91 ? _double_bytes_0_T_13 : _GEN_407; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_409 = 7'h22 == _GEN_91 ? _double_bytes_0_T_14 : _GEN_408; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_410 = 7'h23 == _GEN_91 ? _double_bytes_0_T_15 : _GEN_409; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_411 = 7'h24 == _GEN_91 ? _double_bytes_0_T_16 : _GEN_410; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_412 = 7'h25 == _GEN_91 ? _double_bytes_0_T_17 : _GEN_411; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_413 = 7'h26 == _GEN_91 ? _double_bytes_0_T_18 : _GEN_412; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_414 = 7'h27 == _GEN_91 ? _double_bytes_0_T_19 : _GEN_413; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_415 = 7'h28 == _GEN_91 ? _double_bytes_0_T_20 : _GEN_414; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_416 = 7'h29 == _GEN_91 ? _double_bytes_0_T_21 : _GEN_415; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_417 = 7'h2a == _GEN_91 ? _double_bytes_0_T_22 : _GEN_416; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_418 = 7'h2b == _GEN_91 ? _double_bytes_0_T_23 : _GEN_417; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_419 = 7'h2c == _GEN_91 ? _double_bytes_0_T_24 : _GEN_418; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_420 = 7'h2d == _GEN_91 ? _double_bytes_0_T_25 : _GEN_419; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_421 = 7'h2e == _GEN_91 ? _double_bytes_0_T_26 : _GEN_420; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_422 = 7'h2f == _GEN_91 ? _double_bytes_0_T_27 : _GEN_421; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_423 = 7'h30 == _GEN_91 ? _double_bytes_0_T_28 : _GEN_422; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_424 = 7'h31 == _GEN_91 ? _double_bytes_0_T_29 : _GEN_423; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_1_1 = _GEN_67 ? _GEN_424 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [31:0] _groups_1_T_1 = {double_bytes_1_0,double_bytes_1_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_426 = _GEN_57 == 2'h2 ? _groups_1_T_1 : _GEN_363; // @[matcher_pisa.scala 131:50 matcher_pisa.scala 145:31]
  wire [31:0] _GEN_427 = 7'h32 == _GEN_90 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39 matcher_pisa.scala 150:31]
  wire [31:0] _GEN_428 = 7'h33 == _GEN_90 ? _groups_0_T_3 : _GEN_427; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_429 = 7'h34 == _GEN_90 ? _groups_0_T_4 : _GEN_428; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_430 = 7'h35 == _GEN_90 ? _groups_0_T_5 : _GEN_429; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_431 = 7'h36 == _GEN_90 ? _groups_0_T_6 : _GEN_430; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_432 = 7'h37 == _GEN_90 ? _groups_0_T_7 : _GEN_431; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_433 = 7'h38 == _GEN_90 ? _groups_0_T_8 : _GEN_432; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_434 = 7'h39 == _GEN_90 ? _groups_0_T_9 : _GEN_433; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_435 = 7'h3a == _GEN_90 ? _groups_0_T_10 : _GEN_434; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_436 = 7'h3b == _GEN_90 ? _groups_0_T_11 : _GEN_435; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_437 = 7'h3c == _GEN_90 ? _groups_0_T_12 : _GEN_436; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_438 = 7'h3d == _GEN_90 ? _groups_0_T_13 : _GEN_437; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_439 = 7'h3e == _GEN_90 ? _groups_0_T_14 : _GEN_438; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_440 = 7'h3f == _GEN_90 ? _groups_0_T_15 : _GEN_439; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_441 = 7'h40 == _GEN_90 ? _groups_0_T_16 : _GEN_440; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_442 = 7'h41 == _GEN_90 ? _groups_0_T_17 : _GEN_441; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_443 = 7'h42 == _GEN_90 ? _groups_0_T_18 : _GEN_442; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_444 = 7'h43 == _GEN_90 ? _groups_0_T_19 : _GEN_443; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_445 = 7'h44 == _GEN_90 ? _groups_0_T_20 : _GEN_444; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_446 = 7'h45 == _GEN_90 ? _groups_0_T_21 : _GEN_445; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] groups_1 = _GEN_57 == 2'h3 ? _GEN_446 : _GEN_426; // @[matcher_pisa.scala 147:50]
  wire [7:0] _GEN_448 = 7'h0 == _GEN_94 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_449 = 7'h1 == _GEN_94 ? phv_data_1 : _GEN_448; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_450 = 7'h2 == _GEN_94 ? phv_data_2 : _GEN_449; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_451 = 7'h3 == _GEN_94 ? phv_data_3 : _GEN_450; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_452 = 7'h4 == _GEN_94 ? phv_data_4 : _GEN_451; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_453 = 7'h5 == _GEN_94 ? phv_data_5 : _GEN_452; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_454 = 7'h6 == _GEN_94 ? phv_data_6 : _GEN_453; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_455 = 7'h7 == _GEN_94 ? phv_data_7 : _GEN_454; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_456 = 7'h8 == _GEN_94 ? phv_data_8 : _GEN_455; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_457 = 7'h9 == _GEN_94 ? phv_data_9 : _GEN_456; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_458 = 7'ha == _GEN_94 ? phv_data_10 : _GEN_457; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_459 = 7'hb == _GEN_94 ? phv_data_11 : _GEN_458; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_460 = 7'hc == _GEN_94 ? phv_data_12 : _GEN_459; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_461 = 7'hd == _GEN_94 ? phv_data_13 : _GEN_460; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_462 = 7'he == _GEN_94 ? phv_data_14 : _GEN_461; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_463 = 7'hf == _GEN_94 ? phv_data_15 : _GEN_462; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_464 = 7'h10 == _GEN_94 ? phv_data_16 : _GEN_463; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_465 = 7'h11 == _GEN_94 ? phv_data_17 : _GEN_464; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_466 = 7'h12 == _GEN_94 ? phv_data_18 : _GEN_465; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_467 = 7'h13 == _GEN_94 ? phv_data_19 : _GEN_466; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_2_0 = _GEN_70 ? _GEN_467 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_469 = 7'h0 == _GEN_95 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_470 = 7'h1 == _GEN_95 ? phv_data_1 : _GEN_469; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_471 = 7'h2 == _GEN_95 ? phv_data_2 : _GEN_470; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_472 = 7'h3 == _GEN_95 ? phv_data_3 : _GEN_471; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_473 = 7'h4 == _GEN_95 ? phv_data_4 : _GEN_472; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_474 = 7'h5 == _GEN_95 ? phv_data_5 : _GEN_473; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_475 = 7'h6 == _GEN_95 ? phv_data_6 : _GEN_474; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_476 = 7'h7 == _GEN_95 ? phv_data_7 : _GEN_475; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_477 = 7'h8 == _GEN_95 ? phv_data_8 : _GEN_476; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_478 = 7'h9 == _GEN_95 ? phv_data_9 : _GEN_477; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_479 = 7'ha == _GEN_95 ? phv_data_10 : _GEN_478; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_480 = 7'hb == _GEN_95 ? phv_data_11 : _GEN_479; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_481 = 7'hc == _GEN_95 ? phv_data_12 : _GEN_480; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_482 = 7'hd == _GEN_95 ? phv_data_13 : _GEN_481; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_483 = 7'he == _GEN_95 ? phv_data_14 : _GEN_482; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_484 = 7'hf == _GEN_95 ? phv_data_15 : _GEN_483; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_485 = 7'h10 == _GEN_95 ? phv_data_16 : _GEN_484; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_486 = 7'h11 == _GEN_95 ? phv_data_17 : _GEN_485; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_487 = 7'h12 == _GEN_95 ? phv_data_18 : _GEN_486; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_488 = 7'h13 == _GEN_95 ? phv_data_19 : _GEN_487; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_2_1 = _GEN_71 ? _GEN_488 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_490 = 7'h0 == _GEN_96 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_491 = 7'h1 == _GEN_96 ? phv_data_1 : _GEN_490; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_492 = 7'h2 == _GEN_96 ? phv_data_2 : _GEN_491; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_493 = 7'h3 == _GEN_96 ? phv_data_3 : _GEN_492; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_494 = 7'h4 == _GEN_96 ? phv_data_4 : _GEN_493; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_495 = 7'h5 == _GEN_96 ? phv_data_5 : _GEN_494; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_496 = 7'h6 == _GEN_96 ? phv_data_6 : _GEN_495; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_497 = 7'h7 == _GEN_96 ? phv_data_7 : _GEN_496; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_498 = 7'h8 == _GEN_96 ? phv_data_8 : _GEN_497; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_499 = 7'h9 == _GEN_96 ? phv_data_9 : _GEN_498; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_500 = 7'ha == _GEN_96 ? phv_data_10 : _GEN_499; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_501 = 7'hb == _GEN_96 ? phv_data_11 : _GEN_500; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_502 = 7'hc == _GEN_96 ? phv_data_12 : _GEN_501; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_503 = 7'hd == _GEN_96 ? phv_data_13 : _GEN_502; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_504 = 7'he == _GEN_96 ? phv_data_14 : _GEN_503; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_505 = 7'hf == _GEN_96 ? phv_data_15 : _GEN_504; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_506 = 7'h10 == _GEN_96 ? phv_data_16 : _GEN_505; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_507 = 7'h11 == _GEN_96 ? phv_data_17 : _GEN_506; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_508 = 7'h12 == _GEN_96 ? phv_data_18 : _GEN_507; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_509 = 7'h13 == _GEN_96 ? phv_data_19 : _GEN_508; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_2_2 = _GEN_72 ? _GEN_509 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_511 = 7'h0 == _GEN_97 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_512 = 7'h1 == _GEN_97 ? phv_data_1 : _GEN_511; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_513 = 7'h2 == _GEN_97 ? phv_data_2 : _GEN_512; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_514 = 7'h3 == _GEN_97 ? phv_data_3 : _GEN_513; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_515 = 7'h4 == _GEN_97 ? phv_data_4 : _GEN_514; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_516 = 7'h5 == _GEN_97 ? phv_data_5 : _GEN_515; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_517 = 7'h6 == _GEN_97 ? phv_data_6 : _GEN_516; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_518 = 7'h7 == _GEN_97 ? phv_data_7 : _GEN_517; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_519 = 7'h8 == _GEN_97 ? phv_data_8 : _GEN_518; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_520 = 7'h9 == _GEN_97 ? phv_data_9 : _GEN_519; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_521 = 7'ha == _GEN_97 ? phv_data_10 : _GEN_520; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_522 = 7'hb == _GEN_97 ? phv_data_11 : _GEN_521; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_523 = 7'hc == _GEN_97 ? phv_data_12 : _GEN_522; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_524 = 7'hd == _GEN_97 ? phv_data_13 : _GEN_523; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_525 = 7'he == _GEN_97 ? phv_data_14 : _GEN_524; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_526 = 7'hf == _GEN_97 ? phv_data_15 : _GEN_525; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_527 = 7'h10 == _GEN_97 ? phv_data_16 : _GEN_526; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_528 = 7'h11 == _GEN_97 ? phv_data_17 : _GEN_527; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_529 = 7'h12 == _GEN_97 ? phv_data_18 : _GEN_528; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_530 = 7'h13 == _GEN_97 ? phv_data_19 : _GEN_529; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_2_3 = _GEN_73 ? _GEN_530 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [31:0] _groups_2_T = {bytes_2_0,bytes_2_1,bytes_2_2,bytes_2_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_532 = _GEN_58 == 2'h1 ? _groups_2_T : 32'h0; // @[matcher_pisa.scala 115:50 matcher_pisa.scala 129:31 matcher_pisa.scala 114:27]
  wire [15:0] _GEN_533 = 7'h14 == _GEN_94 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_534 = 7'h15 == _GEN_94 ? _double_bytes_0_T_1 : _GEN_533; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_535 = 7'h16 == _GEN_94 ? _double_bytes_0_T_2 : _GEN_534; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_536 = 7'h17 == _GEN_94 ? _double_bytes_0_T_3 : _GEN_535; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_537 = 7'h18 == _GEN_94 ? _double_bytes_0_T_4 : _GEN_536; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_538 = 7'h19 == _GEN_94 ? _double_bytes_0_T_5 : _GEN_537; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_539 = 7'h1a == _GEN_94 ? _double_bytes_0_T_6 : _GEN_538; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_540 = 7'h1b == _GEN_94 ? _double_bytes_0_T_7 : _GEN_539; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_541 = 7'h1c == _GEN_94 ? _double_bytes_0_T_8 : _GEN_540; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_542 = 7'h1d == _GEN_94 ? _double_bytes_0_T_9 : _GEN_541; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_543 = 7'h1e == _GEN_94 ? _double_bytes_0_T_10 : _GEN_542; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_544 = 7'h1f == _GEN_94 ? _double_bytes_0_T_11 : _GEN_543; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_545 = 7'h20 == _GEN_94 ? _double_bytes_0_T_12 : _GEN_544; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_546 = 7'h21 == _GEN_94 ? _double_bytes_0_T_13 : _GEN_545; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_547 = 7'h22 == _GEN_94 ? _double_bytes_0_T_14 : _GEN_546; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_548 = 7'h23 == _GEN_94 ? _double_bytes_0_T_15 : _GEN_547; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_549 = 7'h24 == _GEN_94 ? _double_bytes_0_T_16 : _GEN_548; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_550 = 7'h25 == _GEN_94 ? _double_bytes_0_T_17 : _GEN_549; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_551 = 7'h26 == _GEN_94 ? _double_bytes_0_T_18 : _GEN_550; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_552 = 7'h27 == _GEN_94 ? _double_bytes_0_T_19 : _GEN_551; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_553 = 7'h28 == _GEN_94 ? _double_bytes_0_T_20 : _GEN_552; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_554 = 7'h29 == _GEN_94 ? _double_bytes_0_T_21 : _GEN_553; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_555 = 7'h2a == _GEN_94 ? _double_bytes_0_T_22 : _GEN_554; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_556 = 7'h2b == _GEN_94 ? _double_bytes_0_T_23 : _GEN_555; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_557 = 7'h2c == _GEN_94 ? _double_bytes_0_T_24 : _GEN_556; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_558 = 7'h2d == _GEN_94 ? _double_bytes_0_T_25 : _GEN_557; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_559 = 7'h2e == _GEN_94 ? _double_bytes_0_T_26 : _GEN_558; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_560 = 7'h2f == _GEN_94 ? _double_bytes_0_T_27 : _GEN_559; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_561 = 7'h30 == _GEN_94 ? _double_bytes_0_T_28 : _GEN_560; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_562 = 7'h31 == _GEN_94 ? _double_bytes_0_T_29 : _GEN_561; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_2_0 = _GEN_70 ? _GEN_562 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_564 = 7'h14 == _GEN_95 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_565 = 7'h15 == _GEN_95 ? _double_bytes_0_T_1 : _GEN_564; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_566 = 7'h16 == _GEN_95 ? _double_bytes_0_T_2 : _GEN_565; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_567 = 7'h17 == _GEN_95 ? _double_bytes_0_T_3 : _GEN_566; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_568 = 7'h18 == _GEN_95 ? _double_bytes_0_T_4 : _GEN_567; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_569 = 7'h19 == _GEN_95 ? _double_bytes_0_T_5 : _GEN_568; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_570 = 7'h1a == _GEN_95 ? _double_bytes_0_T_6 : _GEN_569; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_571 = 7'h1b == _GEN_95 ? _double_bytes_0_T_7 : _GEN_570; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_572 = 7'h1c == _GEN_95 ? _double_bytes_0_T_8 : _GEN_571; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_573 = 7'h1d == _GEN_95 ? _double_bytes_0_T_9 : _GEN_572; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_574 = 7'h1e == _GEN_95 ? _double_bytes_0_T_10 : _GEN_573; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_575 = 7'h1f == _GEN_95 ? _double_bytes_0_T_11 : _GEN_574; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_576 = 7'h20 == _GEN_95 ? _double_bytes_0_T_12 : _GEN_575; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_577 = 7'h21 == _GEN_95 ? _double_bytes_0_T_13 : _GEN_576; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_578 = 7'h22 == _GEN_95 ? _double_bytes_0_T_14 : _GEN_577; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_579 = 7'h23 == _GEN_95 ? _double_bytes_0_T_15 : _GEN_578; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_580 = 7'h24 == _GEN_95 ? _double_bytes_0_T_16 : _GEN_579; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_581 = 7'h25 == _GEN_95 ? _double_bytes_0_T_17 : _GEN_580; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_582 = 7'h26 == _GEN_95 ? _double_bytes_0_T_18 : _GEN_581; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_583 = 7'h27 == _GEN_95 ? _double_bytes_0_T_19 : _GEN_582; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_584 = 7'h28 == _GEN_95 ? _double_bytes_0_T_20 : _GEN_583; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_585 = 7'h29 == _GEN_95 ? _double_bytes_0_T_21 : _GEN_584; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_586 = 7'h2a == _GEN_95 ? _double_bytes_0_T_22 : _GEN_585; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_587 = 7'h2b == _GEN_95 ? _double_bytes_0_T_23 : _GEN_586; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_588 = 7'h2c == _GEN_95 ? _double_bytes_0_T_24 : _GEN_587; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_589 = 7'h2d == _GEN_95 ? _double_bytes_0_T_25 : _GEN_588; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_590 = 7'h2e == _GEN_95 ? _double_bytes_0_T_26 : _GEN_589; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_591 = 7'h2f == _GEN_95 ? _double_bytes_0_T_27 : _GEN_590; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_592 = 7'h30 == _GEN_95 ? _double_bytes_0_T_28 : _GEN_591; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_593 = 7'h31 == _GEN_95 ? _double_bytes_0_T_29 : _GEN_592; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_2_1 = _GEN_71 ? _GEN_593 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [31:0] _groups_2_T_1 = {double_bytes_2_0,double_bytes_2_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_595 = _GEN_58 == 2'h2 ? _groups_2_T_1 : _GEN_532; // @[matcher_pisa.scala 131:50 matcher_pisa.scala 145:31]
  wire [31:0] _GEN_596 = 7'h32 == _GEN_94 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39 matcher_pisa.scala 150:31]
  wire [31:0] _GEN_597 = 7'h33 == _GEN_94 ? _groups_0_T_3 : _GEN_596; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_598 = 7'h34 == _GEN_94 ? _groups_0_T_4 : _GEN_597; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_599 = 7'h35 == _GEN_94 ? _groups_0_T_5 : _GEN_598; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_600 = 7'h36 == _GEN_94 ? _groups_0_T_6 : _GEN_599; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_601 = 7'h37 == _GEN_94 ? _groups_0_T_7 : _GEN_600; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_602 = 7'h38 == _GEN_94 ? _groups_0_T_8 : _GEN_601; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_603 = 7'h39 == _GEN_94 ? _groups_0_T_9 : _GEN_602; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_604 = 7'h3a == _GEN_94 ? _groups_0_T_10 : _GEN_603; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_605 = 7'h3b == _GEN_94 ? _groups_0_T_11 : _GEN_604; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_606 = 7'h3c == _GEN_94 ? _groups_0_T_12 : _GEN_605; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_607 = 7'h3d == _GEN_94 ? _groups_0_T_13 : _GEN_606; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_608 = 7'h3e == _GEN_94 ? _groups_0_T_14 : _GEN_607; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_609 = 7'h3f == _GEN_94 ? _groups_0_T_15 : _GEN_608; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_610 = 7'h40 == _GEN_94 ? _groups_0_T_16 : _GEN_609; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_611 = 7'h41 == _GEN_94 ? _groups_0_T_17 : _GEN_610; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_612 = 7'h42 == _GEN_94 ? _groups_0_T_18 : _GEN_611; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_613 = 7'h43 == _GEN_94 ? _groups_0_T_19 : _GEN_612; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_614 = 7'h44 == _GEN_94 ? _groups_0_T_20 : _GEN_613; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_615 = 7'h45 == _GEN_94 ? _groups_0_T_21 : _GEN_614; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] groups_2 = _GEN_58 == 2'h3 ? _GEN_615 : _GEN_595; // @[matcher_pisa.scala 147:50]
  wire [7:0] _GEN_617 = 7'h0 == _GEN_98 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_618 = 7'h1 == _GEN_98 ? phv_data_1 : _GEN_617; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_619 = 7'h2 == _GEN_98 ? phv_data_2 : _GEN_618; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_620 = 7'h3 == _GEN_98 ? phv_data_3 : _GEN_619; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_621 = 7'h4 == _GEN_98 ? phv_data_4 : _GEN_620; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_622 = 7'h5 == _GEN_98 ? phv_data_5 : _GEN_621; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_623 = 7'h6 == _GEN_98 ? phv_data_6 : _GEN_622; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_624 = 7'h7 == _GEN_98 ? phv_data_7 : _GEN_623; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_625 = 7'h8 == _GEN_98 ? phv_data_8 : _GEN_624; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_626 = 7'h9 == _GEN_98 ? phv_data_9 : _GEN_625; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_627 = 7'ha == _GEN_98 ? phv_data_10 : _GEN_626; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_628 = 7'hb == _GEN_98 ? phv_data_11 : _GEN_627; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_629 = 7'hc == _GEN_98 ? phv_data_12 : _GEN_628; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_630 = 7'hd == _GEN_98 ? phv_data_13 : _GEN_629; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_631 = 7'he == _GEN_98 ? phv_data_14 : _GEN_630; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_632 = 7'hf == _GEN_98 ? phv_data_15 : _GEN_631; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_633 = 7'h10 == _GEN_98 ? phv_data_16 : _GEN_632; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_634 = 7'h11 == _GEN_98 ? phv_data_17 : _GEN_633; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_635 = 7'h12 == _GEN_98 ? phv_data_18 : _GEN_634; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_636 = 7'h13 == _GEN_98 ? phv_data_19 : _GEN_635; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_3_0 = _GEN_74 ? _GEN_636 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_638 = 7'h0 == _GEN_99 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_639 = 7'h1 == _GEN_99 ? phv_data_1 : _GEN_638; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_640 = 7'h2 == _GEN_99 ? phv_data_2 : _GEN_639; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_641 = 7'h3 == _GEN_99 ? phv_data_3 : _GEN_640; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_642 = 7'h4 == _GEN_99 ? phv_data_4 : _GEN_641; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_643 = 7'h5 == _GEN_99 ? phv_data_5 : _GEN_642; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_644 = 7'h6 == _GEN_99 ? phv_data_6 : _GEN_643; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_645 = 7'h7 == _GEN_99 ? phv_data_7 : _GEN_644; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_646 = 7'h8 == _GEN_99 ? phv_data_8 : _GEN_645; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_647 = 7'h9 == _GEN_99 ? phv_data_9 : _GEN_646; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_648 = 7'ha == _GEN_99 ? phv_data_10 : _GEN_647; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_649 = 7'hb == _GEN_99 ? phv_data_11 : _GEN_648; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_650 = 7'hc == _GEN_99 ? phv_data_12 : _GEN_649; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_651 = 7'hd == _GEN_99 ? phv_data_13 : _GEN_650; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_652 = 7'he == _GEN_99 ? phv_data_14 : _GEN_651; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_653 = 7'hf == _GEN_99 ? phv_data_15 : _GEN_652; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_654 = 7'h10 == _GEN_99 ? phv_data_16 : _GEN_653; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_655 = 7'h11 == _GEN_99 ? phv_data_17 : _GEN_654; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_656 = 7'h12 == _GEN_99 ? phv_data_18 : _GEN_655; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_657 = 7'h13 == _GEN_99 ? phv_data_19 : _GEN_656; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_3_1 = _GEN_75 ? _GEN_657 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_659 = 7'h0 == _GEN_100 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_660 = 7'h1 == _GEN_100 ? phv_data_1 : _GEN_659; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_661 = 7'h2 == _GEN_100 ? phv_data_2 : _GEN_660; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_662 = 7'h3 == _GEN_100 ? phv_data_3 : _GEN_661; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_663 = 7'h4 == _GEN_100 ? phv_data_4 : _GEN_662; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_664 = 7'h5 == _GEN_100 ? phv_data_5 : _GEN_663; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_665 = 7'h6 == _GEN_100 ? phv_data_6 : _GEN_664; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_666 = 7'h7 == _GEN_100 ? phv_data_7 : _GEN_665; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_667 = 7'h8 == _GEN_100 ? phv_data_8 : _GEN_666; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_668 = 7'h9 == _GEN_100 ? phv_data_9 : _GEN_667; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_669 = 7'ha == _GEN_100 ? phv_data_10 : _GEN_668; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_670 = 7'hb == _GEN_100 ? phv_data_11 : _GEN_669; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_671 = 7'hc == _GEN_100 ? phv_data_12 : _GEN_670; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_672 = 7'hd == _GEN_100 ? phv_data_13 : _GEN_671; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_673 = 7'he == _GEN_100 ? phv_data_14 : _GEN_672; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_674 = 7'hf == _GEN_100 ? phv_data_15 : _GEN_673; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_675 = 7'h10 == _GEN_100 ? phv_data_16 : _GEN_674; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_676 = 7'h11 == _GEN_100 ? phv_data_17 : _GEN_675; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_677 = 7'h12 == _GEN_100 ? phv_data_18 : _GEN_676; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_678 = 7'h13 == _GEN_100 ? phv_data_19 : _GEN_677; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_3_2 = _GEN_76 ? _GEN_678 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_680 = 7'h0 == _GEN_101 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_681 = 7'h1 == _GEN_101 ? phv_data_1 : _GEN_680; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_682 = 7'h2 == _GEN_101 ? phv_data_2 : _GEN_681; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_683 = 7'h3 == _GEN_101 ? phv_data_3 : _GEN_682; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_684 = 7'h4 == _GEN_101 ? phv_data_4 : _GEN_683; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_685 = 7'h5 == _GEN_101 ? phv_data_5 : _GEN_684; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_686 = 7'h6 == _GEN_101 ? phv_data_6 : _GEN_685; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_687 = 7'h7 == _GEN_101 ? phv_data_7 : _GEN_686; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_688 = 7'h8 == _GEN_101 ? phv_data_8 : _GEN_687; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_689 = 7'h9 == _GEN_101 ? phv_data_9 : _GEN_688; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_690 = 7'ha == _GEN_101 ? phv_data_10 : _GEN_689; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_691 = 7'hb == _GEN_101 ? phv_data_11 : _GEN_690; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_692 = 7'hc == _GEN_101 ? phv_data_12 : _GEN_691; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_693 = 7'hd == _GEN_101 ? phv_data_13 : _GEN_692; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_694 = 7'he == _GEN_101 ? phv_data_14 : _GEN_693; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_695 = 7'hf == _GEN_101 ? phv_data_15 : _GEN_694; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_696 = 7'h10 == _GEN_101 ? phv_data_16 : _GEN_695; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_697 = 7'h11 == _GEN_101 ? phv_data_17 : _GEN_696; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_698 = 7'h12 == _GEN_101 ? phv_data_18 : _GEN_697; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_699 = 7'h13 == _GEN_101 ? phv_data_19 : _GEN_698; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_3_3 = _GEN_77 ? _GEN_699 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [31:0] _groups_3_T = {bytes_3_0,bytes_3_1,bytes_3_2,bytes_3_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_701 = _GEN_59 == 2'h1 ? _groups_3_T : 32'h0; // @[matcher_pisa.scala 115:50 matcher_pisa.scala 129:31 matcher_pisa.scala 114:27]
  wire [15:0] _GEN_702 = 7'h14 == _GEN_98 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_703 = 7'h15 == _GEN_98 ? _double_bytes_0_T_1 : _GEN_702; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_704 = 7'h16 == _GEN_98 ? _double_bytes_0_T_2 : _GEN_703; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_705 = 7'h17 == _GEN_98 ? _double_bytes_0_T_3 : _GEN_704; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_706 = 7'h18 == _GEN_98 ? _double_bytes_0_T_4 : _GEN_705; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_707 = 7'h19 == _GEN_98 ? _double_bytes_0_T_5 : _GEN_706; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_708 = 7'h1a == _GEN_98 ? _double_bytes_0_T_6 : _GEN_707; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_709 = 7'h1b == _GEN_98 ? _double_bytes_0_T_7 : _GEN_708; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_710 = 7'h1c == _GEN_98 ? _double_bytes_0_T_8 : _GEN_709; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_711 = 7'h1d == _GEN_98 ? _double_bytes_0_T_9 : _GEN_710; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_712 = 7'h1e == _GEN_98 ? _double_bytes_0_T_10 : _GEN_711; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_713 = 7'h1f == _GEN_98 ? _double_bytes_0_T_11 : _GEN_712; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_714 = 7'h20 == _GEN_98 ? _double_bytes_0_T_12 : _GEN_713; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_715 = 7'h21 == _GEN_98 ? _double_bytes_0_T_13 : _GEN_714; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_716 = 7'h22 == _GEN_98 ? _double_bytes_0_T_14 : _GEN_715; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_717 = 7'h23 == _GEN_98 ? _double_bytes_0_T_15 : _GEN_716; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_718 = 7'h24 == _GEN_98 ? _double_bytes_0_T_16 : _GEN_717; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_719 = 7'h25 == _GEN_98 ? _double_bytes_0_T_17 : _GEN_718; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_720 = 7'h26 == _GEN_98 ? _double_bytes_0_T_18 : _GEN_719; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_721 = 7'h27 == _GEN_98 ? _double_bytes_0_T_19 : _GEN_720; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_722 = 7'h28 == _GEN_98 ? _double_bytes_0_T_20 : _GEN_721; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_723 = 7'h29 == _GEN_98 ? _double_bytes_0_T_21 : _GEN_722; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_724 = 7'h2a == _GEN_98 ? _double_bytes_0_T_22 : _GEN_723; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_725 = 7'h2b == _GEN_98 ? _double_bytes_0_T_23 : _GEN_724; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_726 = 7'h2c == _GEN_98 ? _double_bytes_0_T_24 : _GEN_725; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_727 = 7'h2d == _GEN_98 ? _double_bytes_0_T_25 : _GEN_726; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_728 = 7'h2e == _GEN_98 ? _double_bytes_0_T_26 : _GEN_727; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_729 = 7'h2f == _GEN_98 ? _double_bytes_0_T_27 : _GEN_728; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_730 = 7'h30 == _GEN_98 ? _double_bytes_0_T_28 : _GEN_729; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_731 = 7'h31 == _GEN_98 ? _double_bytes_0_T_29 : _GEN_730; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_3_0 = _GEN_74 ? _GEN_731 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_733 = 7'h14 == _GEN_99 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_734 = 7'h15 == _GEN_99 ? _double_bytes_0_T_1 : _GEN_733; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_735 = 7'h16 == _GEN_99 ? _double_bytes_0_T_2 : _GEN_734; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_736 = 7'h17 == _GEN_99 ? _double_bytes_0_T_3 : _GEN_735; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_737 = 7'h18 == _GEN_99 ? _double_bytes_0_T_4 : _GEN_736; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_738 = 7'h19 == _GEN_99 ? _double_bytes_0_T_5 : _GEN_737; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_739 = 7'h1a == _GEN_99 ? _double_bytes_0_T_6 : _GEN_738; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_740 = 7'h1b == _GEN_99 ? _double_bytes_0_T_7 : _GEN_739; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_741 = 7'h1c == _GEN_99 ? _double_bytes_0_T_8 : _GEN_740; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_742 = 7'h1d == _GEN_99 ? _double_bytes_0_T_9 : _GEN_741; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_743 = 7'h1e == _GEN_99 ? _double_bytes_0_T_10 : _GEN_742; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_744 = 7'h1f == _GEN_99 ? _double_bytes_0_T_11 : _GEN_743; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_745 = 7'h20 == _GEN_99 ? _double_bytes_0_T_12 : _GEN_744; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_746 = 7'h21 == _GEN_99 ? _double_bytes_0_T_13 : _GEN_745; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_747 = 7'h22 == _GEN_99 ? _double_bytes_0_T_14 : _GEN_746; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_748 = 7'h23 == _GEN_99 ? _double_bytes_0_T_15 : _GEN_747; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_749 = 7'h24 == _GEN_99 ? _double_bytes_0_T_16 : _GEN_748; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_750 = 7'h25 == _GEN_99 ? _double_bytes_0_T_17 : _GEN_749; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_751 = 7'h26 == _GEN_99 ? _double_bytes_0_T_18 : _GEN_750; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_752 = 7'h27 == _GEN_99 ? _double_bytes_0_T_19 : _GEN_751; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_753 = 7'h28 == _GEN_99 ? _double_bytes_0_T_20 : _GEN_752; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_754 = 7'h29 == _GEN_99 ? _double_bytes_0_T_21 : _GEN_753; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_755 = 7'h2a == _GEN_99 ? _double_bytes_0_T_22 : _GEN_754; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_756 = 7'h2b == _GEN_99 ? _double_bytes_0_T_23 : _GEN_755; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_757 = 7'h2c == _GEN_99 ? _double_bytes_0_T_24 : _GEN_756; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_758 = 7'h2d == _GEN_99 ? _double_bytes_0_T_25 : _GEN_757; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_759 = 7'h2e == _GEN_99 ? _double_bytes_0_T_26 : _GEN_758; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_760 = 7'h2f == _GEN_99 ? _double_bytes_0_T_27 : _GEN_759; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_761 = 7'h30 == _GEN_99 ? _double_bytes_0_T_28 : _GEN_760; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_762 = 7'h31 == _GEN_99 ? _double_bytes_0_T_29 : _GEN_761; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_3_1 = _GEN_75 ? _GEN_762 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [31:0] _groups_3_T_1 = {double_bytes_3_0,double_bytes_3_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_764 = _GEN_59 == 2'h2 ? _groups_3_T_1 : _GEN_701; // @[matcher_pisa.scala 131:50 matcher_pisa.scala 145:31]
  wire [31:0] _GEN_765 = 7'h32 == _GEN_98 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39 matcher_pisa.scala 150:31]
  wire [31:0] _GEN_766 = 7'h33 == _GEN_98 ? _groups_0_T_3 : _GEN_765; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_767 = 7'h34 == _GEN_98 ? _groups_0_T_4 : _GEN_766; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_768 = 7'h35 == _GEN_98 ? _groups_0_T_5 : _GEN_767; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_769 = 7'h36 == _GEN_98 ? _groups_0_T_6 : _GEN_768; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_770 = 7'h37 == _GEN_98 ? _groups_0_T_7 : _GEN_769; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_771 = 7'h38 == _GEN_98 ? _groups_0_T_8 : _GEN_770; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_772 = 7'h39 == _GEN_98 ? _groups_0_T_9 : _GEN_771; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_773 = 7'h3a == _GEN_98 ? _groups_0_T_10 : _GEN_772; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_774 = 7'h3b == _GEN_98 ? _groups_0_T_11 : _GEN_773; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_775 = 7'h3c == _GEN_98 ? _groups_0_T_12 : _GEN_774; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_776 = 7'h3d == _GEN_98 ? _groups_0_T_13 : _GEN_775; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_777 = 7'h3e == _GEN_98 ? _groups_0_T_14 : _GEN_776; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_778 = 7'h3f == _GEN_98 ? _groups_0_T_15 : _GEN_777; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_779 = 7'h40 == _GEN_98 ? _groups_0_T_16 : _GEN_778; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_780 = 7'h41 == _GEN_98 ? _groups_0_T_17 : _GEN_779; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_781 = 7'h42 == _GEN_98 ? _groups_0_T_18 : _GEN_780; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_782 = 7'h43 == _GEN_98 ? _groups_0_T_19 : _GEN_781; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_783 = 7'h44 == _GEN_98 ? _groups_0_T_20 : _GEN_782; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_784 = 7'h45 == _GEN_98 ? _groups_0_T_21 : _GEN_783; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] groups_3 = _GEN_59 == 2'h3 ? _GEN_784 : _GEN_764; // @[matcher_pisa.scala 147:50]
  wire [7:0] _GEN_786 = 7'h0 == _GEN_102 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_787 = 7'h1 == _GEN_102 ? phv_data_1 : _GEN_786; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_788 = 7'h2 == _GEN_102 ? phv_data_2 : _GEN_787; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_789 = 7'h3 == _GEN_102 ? phv_data_3 : _GEN_788; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_790 = 7'h4 == _GEN_102 ? phv_data_4 : _GEN_789; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_791 = 7'h5 == _GEN_102 ? phv_data_5 : _GEN_790; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_792 = 7'h6 == _GEN_102 ? phv_data_6 : _GEN_791; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_793 = 7'h7 == _GEN_102 ? phv_data_7 : _GEN_792; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_794 = 7'h8 == _GEN_102 ? phv_data_8 : _GEN_793; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_795 = 7'h9 == _GEN_102 ? phv_data_9 : _GEN_794; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_796 = 7'ha == _GEN_102 ? phv_data_10 : _GEN_795; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_797 = 7'hb == _GEN_102 ? phv_data_11 : _GEN_796; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_798 = 7'hc == _GEN_102 ? phv_data_12 : _GEN_797; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_799 = 7'hd == _GEN_102 ? phv_data_13 : _GEN_798; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_800 = 7'he == _GEN_102 ? phv_data_14 : _GEN_799; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_801 = 7'hf == _GEN_102 ? phv_data_15 : _GEN_800; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_802 = 7'h10 == _GEN_102 ? phv_data_16 : _GEN_801; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_803 = 7'h11 == _GEN_102 ? phv_data_17 : _GEN_802; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_804 = 7'h12 == _GEN_102 ? phv_data_18 : _GEN_803; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_805 = 7'h13 == _GEN_102 ? phv_data_19 : _GEN_804; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_4_0 = _GEN_78 ? _GEN_805 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_807 = 7'h0 == _GEN_103 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_808 = 7'h1 == _GEN_103 ? phv_data_1 : _GEN_807; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_809 = 7'h2 == _GEN_103 ? phv_data_2 : _GEN_808; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_810 = 7'h3 == _GEN_103 ? phv_data_3 : _GEN_809; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_811 = 7'h4 == _GEN_103 ? phv_data_4 : _GEN_810; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_812 = 7'h5 == _GEN_103 ? phv_data_5 : _GEN_811; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_813 = 7'h6 == _GEN_103 ? phv_data_6 : _GEN_812; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_814 = 7'h7 == _GEN_103 ? phv_data_7 : _GEN_813; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_815 = 7'h8 == _GEN_103 ? phv_data_8 : _GEN_814; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_816 = 7'h9 == _GEN_103 ? phv_data_9 : _GEN_815; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_817 = 7'ha == _GEN_103 ? phv_data_10 : _GEN_816; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_818 = 7'hb == _GEN_103 ? phv_data_11 : _GEN_817; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_819 = 7'hc == _GEN_103 ? phv_data_12 : _GEN_818; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_820 = 7'hd == _GEN_103 ? phv_data_13 : _GEN_819; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_821 = 7'he == _GEN_103 ? phv_data_14 : _GEN_820; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_822 = 7'hf == _GEN_103 ? phv_data_15 : _GEN_821; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_823 = 7'h10 == _GEN_103 ? phv_data_16 : _GEN_822; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_824 = 7'h11 == _GEN_103 ? phv_data_17 : _GEN_823; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_825 = 7'h12 == _GEN_103 ? phv_data_18 : _GEN_824; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_826 = 7'h13 == _GEN_103 ? phv_data_19 : _GEN_825; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_4_1 = _GEN_79 ? _GEN_826 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_828 = 7'h0 == _GEN_104 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_829 = 7'h1 == _GEN_104 ? phv_data_1 : _GEN_828; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_830 = 7'h2 == _GEN_104 ? phv_data_2 : _GEN_829; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_831 = 7'h3 == _GEN_104 ? phv_data_3 : _GEN_830; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_832 = 7'h4 == _GEN_104 ? phv_data_4 : _GEN_831; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_833 = 7'h5 == _GEN_104 ? phv_data_5 : _GEN_832; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_834 = 7'h6 == _GEN_104 ? phv_data_6 : _GEN_833; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_835 = 7'h7 == _GEN_104 ? phv_data_7 : _GEN_834; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_836 = 7'h8 == _GEN_104 ? phv_data_8 : _GEN_835; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_837 = 7'h9 == _GEN_104 ? phv_data_9 : _GEN_836; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_838 = 7'ha == _GEN_104 ? phv_data_10 : _GEN_837; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_839 = 7'hb == _GEN_104 ? phv_data_11 : _GEN_838; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_840 = 7'hc == _GEN_104 ? phv_data_12 : _GEN_839; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_841 = 7'hd == _GEN_104 ? phv_data_13 : _GEN_840; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_842 = 7'he == _GEN_104 ? phv_data_14 : _GEN_841; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_843 = 7'hf == _GEN_104 ? phv_data_15 : _GEN_842; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_844 = 7'h10 == _GEN_104 ? phv_data_16 : _GEN_843; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_845 = 7'h11 == _GEN_104 ? phv_data_17 : _GEN_844; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_846 = 7'h12 == _GEN_104 ? phv_data_18 : _GEN_845; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_847 = 7'h13 == _GEN_104 ? phv_data_19 : _GEN_846; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_4_2 = _GEN_80 ? _GEN_847 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_849 = 7'h0 == _GEN_105 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_850 = 7'h1 == _GEN_105 ? phv_data_1 : _GEN_849; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_851 = 7'h2 == _GEN_105 ? phv_data_2 : _GEN_850; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_852 = 7'h3 == _GEN_105 ? phv_data_3 : _GEN_851; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_853 = 7'h4 == _GEN_105 ? phv_data_4 : _GEN_852; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_854 = 7'h5 == _GEN_105 ? phv_data_5 : _GEN_853; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_855 = 7'h6 == _GEN_105 ? phv_data_6 : _GEN_854; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_856 = 7'h7 == _GEN_105 ? phv_data_7 : _GEN_855; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_857 = 7'h8 == _GEN_105 ? phv_data_8 : _GEN_856; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_858 = 7'h9 == _GEN_105 ? phv_data_9 : _GEN_857; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_859 = 7'ha == _GEN_105 ? phv_data_10 : _GEN_858; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_860 = 7'hb == _GEN_105 ? phv_data_11 : _GEN_859; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_861 = 7'hc == _GEN_105 ? phv_data_12 : _GEN_860; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_862 = 7'hd == _GEN_105 ? phv_data_13 : _GEN_861; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_863 = 7'he == _GEN_105 ? phv_data_14 : _GEN_862; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_864 = 7'hf == _GEN_105 ? phv_data_15 : _GEN_863; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_865 = 7'h10 == _GEN_105 ? phv_data_16 : _GEN_864; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_866 = 7'h11 == _GEN_105 ? phv_data_17 : _GEN_865; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_867 = 7'h12 == _GEN_105 ? phv_data_18 : _GEN_866; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_868 = 7'h13 == _GEN_105 ? phv_data_19 : _GEN_867; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_4_3 = _GEN_81 ? _GEN_868 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [31:0] _groups_4_T = {bytes_4_0,bytes_4_1,bytes_4_2,bytes_4_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_870 = _GEN_60 == 2'h1 ? _groups_4_T : 32'h0; // @[matcher_pisa.scala 115:50 matcher_pisa.scala 129:31 matcher_pisa.scala 114:27]
  wire [15:0] _GEN_871 = 7'h14 == _GEN_102 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_872 = 7'h15 == _GEN_102 ? _double_bytes_0_T_1 : _GEN_871; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_873 = 7'h16 == _GEN_102 ? _double_bytes_0_T_2 : _GEN_872; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_874 = 7'h17 == _GEN_102 ? _double_bytes_0_T_3 : _GEN_873; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_875 = 7'h18 == _GEN_102 ? _double_bytes_0_T_4 : _GEN_874; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_876 = 7'h19 == _GEN_102 ? _double_bytes_0_T_5 : _GEN_875; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_877 = 7'h1a == _GEN_102 ? _double_bytes_0_T_6 : _GEN_876; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_878 = 7'h1b == _GEN_102 ? _double_bytes_0_T_7 : _GEN_877; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_879 = 7'h1c == _GEN_102 ? _double_bytes_0_T_8 : _GEN_878; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_880 = 7'h1d == _GEN_102 ? _double_bytes_0_T_9 : _GEN_879; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_881 = 7'h1e == _GEN_102 ? _double_bytes_0_T_10 : _GEN_880; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_882 = 7'h1f == _GEN_102 ? _double_bytes_0_T_11 : _GEN_881; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_883 = 7'h20 == _GEN_102 ? _double_bytes_0_T_12 : _GEN_882; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_884 = 7'h21 == _GEN_102 ? _double_bytes_0_T_13 : _GEN_883; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_885 = 7'h22 == _GEN_102 ? _double_bytes_0_T_14 : _GEN_884; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_886 = 7'h23 == _GEN_102 ? _double_bytes_0_T_15 : _GEN_885; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_887 = 7'h24 == _GEN_102 ? _double_bytes_0_T_16 : _GEN_886; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_888 = 7'h25 == _GEN_102 ? _double_bytes_0_T_17 : _GEN_887; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_889 = 7'h26 == _GEN_102 ? _double_bytes_0_T_18 : _GEN_888; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_890 = 7'h27 == _GEN_102 ? _double_bytes_0_T_19 : _GEN_889; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_891 = 7'h28 == _GEN_102 ? _double_bytes_0_T_20 : _GEN_890; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_892 = 7'h29 == _GEN_102 ? _double_bytes_0_T_21 : _GEN_891; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_893 = 7'h2a == _GEN_102 ? _double_bytes_0_T_22 : _GEN_892; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_894 = 7'h2b == _GEN_102 ? _double_bytes_0_T_23 : _GEN_893; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_895 = 7'h2c == _GEN_102 ? _double_bytes_0_T_24 : _GEN_894; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_896 = 7'h2d == _GEN_102 ? _double_bytes_0_T_25 : _GEN_895; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_897 = 7'h2e == _GEN_102 ? _double_bytes_0_T_26 : _GEN_896; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_898 = 7'h2f == _GEN_102 ? _double_bytes_0_T_27 : _GEN_897; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_899 = 7'h30 == _GEN_102 ? _double_bytes_0_T_28 : _GEN_898; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_900 = 7'h31 == _GEN_102 ? _double_bytes_0_T_29 : _GEN_899; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_4_0 = _GEN_78 ? _GEN_900 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_902 = 7'h14 == _GEN_103 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_903 = 7'h15 == _GEN_103 ? _double_bytes_0_T_1 : _GEN_902; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_904 = 7'h16 == _GEN_103 ? _double_bytes_0_T_2 : _GEN_903; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_905 = 7'h17 == _GEN_103 ? _double_bytes_0_T_3 : _GEN_904; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_906 = 7'h18 == _GEN_103 ? _double_bytes_0_T_4 : _GEN_905; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_907 = 7'h19 == _GEN_103 ? _double_bytes_0_T_5 : _GEN_906; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_908 = 7'h1a == _GEN_103 ? _double_bytes_0_T_6 : _GEN_907; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_909 = 7'h1b == _GEN_103 ? _double_bytes_0_T_7 : _GEN_908; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_910 = 7'h1c == _GEN_103 ? _double_bytes_0_T_8 : _GEN_909; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_911 = 7'h1d == _GEN_103 ? _double_bytes_0_T_9 : _GEN_910; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_912 = 7'h1e == _GEN_103 ? _double_bytes_0_T_10 : _GEN_911; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_913 = 7'h1f == _GEN_103 ? _double_bytes_0_T_11 : _GEN_912; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_914 = 7'h20 == _GEN_103 ? _double_bytes_0_T_12 : _GEN_913; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_915 = 7'h21 == _GEN_103 ? _double_bytes_0_T_13 : _GEN_914; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_916 = 7'h22 == _GEN_103 ? _double_bytes_0_T_14 : _GEN_915; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_917 = 7'h23 == _GEN_103 ? _double_bytes_0_T_15 : _GEN_916; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_918 = 7'h24 == _GEN_103 ? _double_bytes_0_T_16 : _GEN_917; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_919 = 7'h25 == _GEN_103 ? _double_bytes_0_T_17 : _GEN_918; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_920 = 7'h26 == _GEN_103 ? _double_bytes_0_T_18 : _GEN_919; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_921 = 7'h27 == _GEN_103 ? _double_bytes_0_T_19 : _GEN_920; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_922 = 7'h28 == _GEN_103 ? _double_bytes_0_T_20 : _GEN_921; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_923 = 7'h29 == _GEN_103 ? _double_bytes_0_T_21 : _GEN_922; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_924 = 7'h2a == _GEN_103 ? _double_bytes_0_T_22 : _GEN_923; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_925 = 7'h2b == _GEN_103 ? _double_bytes_0_T_23 : _GEN_924; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_926 = 7'h2c == _GEN_103 ? _double_bytes_0_T_24 : _GEN_925; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_927 = 7'h2d == _GEN_103 ? _double_bytes_0_T_25 : _GEN_926; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_928 = 7'h2e == _GEN_103 ? _double_bytes_0_T_26 : _GEN_927; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_929 = 7'h2f == _GEN_103 ? _double_bytes_0_T_27 : _GEN_928; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_930 = 7'h30 == _GEN_103 ? _double_bytes_0_T_28 : _GEN_929; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_931 = 7'h31 == _GEN_103 ? _double_bytes_0_T_29 : _GEN_930; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_4_1 = _GEN_79 ? _GEN_931 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [31:0] _groups_4_T_1 = {double_bytes_4_0,double_bytes_4_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_933 = _GEN_60 == 2'h2 ? _groups_4_T_1 : _GEN_870; // @[matcher_pisa.scala 131:50 matcher_pisa.scala 145:31]
  wire [31:0] _GEN_934 = 7'h32 == _GEN_102 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39 matcher_pisa.scala 150:31]
  wire [31:0] _GEN_935 = 7'h33 == _GEN_102 ? _groups_0_T_3 : _GEN_934; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_936 = 7'h34 == _GEN_102 ? _groups_0_T_4 : _GEN_935; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_937 = 7'h35 == _GEN_102 ? _groups_0_T_5 : _GEN_936; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_938 = 7'h36 == _GEN_102 ? _groups_0_T_6 : _GEN_937; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_939 = 7'h37 == _GEN_102 ? _groups_0_T_7 : _GEN_938; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_940 = 7'h38 == _GEN_102 ? _groups_0_T_8 : _GEN_939; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_941 = 7'h39 == _GEN_102 ? _groups_0_T_9 : _GEN_940; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_942 = 7'h3a == _GEN_102 ? _groups_0_T_10 : _GEN_941; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_943 = 7'h3b == _GEN_102 ? _groups_0_T_11 : _GEN_942; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_944 = 7'h3c == _GEN_102 ? _groups_0_T_12 : _GEN_943; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_945 = 7'h3d == _GEN_102 ? _groups_0_T_13 : _GEN_944; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_946 = 7'h3e == _GEN_102 ? _groups_0_T_14 : _GEN_945; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_947 = 7'h3f == _GEN_102 ? _groups_0_T_15 : _GEN_946; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_948 = 7'h40 == _GEN_102 ? _groups_0_T_16 : _GEN_947; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_949 = 7'h41 == _GEN_102 ? _groups_0_T_17 : _GEN_948; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_950 = 7'h42 == _GEN_102 ? _groups_0_T_18 : _GEN_949; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_951 = 7'h43 == _GEN_102 ? _groups_0_T_19 : _GEN_950; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_952 = 7'h44 == _GEN_102 ? _groups_0_T_20 : _GEN_951; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_953 = 7'h45 == _GEN_102 ? _groups_0_T_21 : _GEN_952; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] groups_4 = _GEN_60 == 2'h3 ? _GEN_953 : _GEN_933; // @[matcher_pisa.scala 147:50]
  wire [7:0] _GEN_955 = 7'h0 == _GEN_106 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_956 = 7'h1 == _GEN_106 ? phv_data_1 : _GEN_955; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_957 = 7'h2 == _GEN_106 ? phv_data_2 : _GEN_956; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_958 = 7'h3 == _GEN_106 ? phv_data_3 : _GEN_957; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_959 = 7'h4 == _GEN_106 ? phv_data_4 : _GEN_958; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_960 = 7'h5 == _GEN_106 ? phv_data_5 : _GEN_959; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_961 = 7'h6 == _GEN_106 ? phv_data_6 : _GEN_960; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_962 = 7'h7 == _GEN_106 ? phv_data_7 : _GEN_961; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_963 = 7'h8 == _GEN_106 ? phv_data_8 : _GEN_962; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_964 = 7'h9 == _GEN_106 ? phv_data_9 : _GEN_963; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_965 = 7'ha == _GEN_106 ? phv_data_10 : _GEN_964; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_966 = 7'hb == _GEN_106 ? phv_data_11 : _GEN_965; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_967 = 7'hc == _GEN_106 ? phv_data_12 : _GEN_966; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_968 = 7'hd == _GEN_106 ? phv_data_13 : _GEN_967; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_969 = 7'he == _GEN_106 ? phv_data_14 : _GEN_968; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_970 = 7'hf == _GEN_106 ? phv_data_15 : _GEN_969; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_971 = 7'h10 == _GEN_106 ? phv_data_16 : _GEN_970; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_972 = 7'h11 == _GEN_106 ? phv_data_17 : _GEN_971; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_973 = 7'h12 == _GEN_106 ? phv_data_18 : _GEN_972; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_974 = 7'h13 == _GEN_106 ? phv_data_19 : _GEN_973; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_5_0 = _GEN_82 ? _GEN_974 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_976 = 7'h0 == _GEN_107 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_977 = 7'h1 == _GEN_107 ? phv_data_1 : _GEN_976; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_978 = 7'h2 == _GEN_107 ? phv_data_2 : _GEN_977; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_979 = 7'h3 == _GEN_107 ? phv_data_3 : _GEN_978; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_980 = 7'h4 == _GEN_107 ? phv_data_4 : _GEN_979; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_981 = 7'h5 == _GEN_107 ? phv_data_5 : _GEN_980; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_982 = 7'h6 == _GEN_107 ? phv_data_6 : _GEN_981; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_983 = 7'h7 == _GEN_107 ? phv_data_7 : _GEN_982; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_984 = 7'h8 == _GEN_107 ? phv_data_8 : _GEN_983; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_985 = 7'h9 == _GEN_107 ? phv_data_9 : _GEN_984; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_986 = 7'ha == _GEN_107 ? phv_data_10 : _GEN_985; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_987 = 7'hb == _GEN_107 ? phv_data_11 : _GEN_986; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_988 = 7'hc == _GEN_107 ? phv_data_12 : _GEN_987; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_989 = 7'hd == _GEN_107 ? phv_data_13 : _GEN_988; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_990 = 7'he == _GEN_107 ? phv_data_14 : _GEN_989; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_991 = 7'hf == _GEN_107 ? phv_data_15 : _GEN_990; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_992 = 7'h10 == _GEN_107 ? phv_data_16 : _GEN_991; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_993 = 7'h11 == _GEN_107 ? phv_data_17 : _GEN_992; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_994 = 7'h12 == _GEN_107 ? phv_data_18 : _GEN_993; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_995 = 7'h13 == _GEN_107 ? phv_data_19 : _GEN_994; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_5_1 = _GEN_83 ? _GEN_995 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_997 = 7'h0 == _GEN_108 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_998 = 7'h1 == _GEN_108 ? phv_data_1 : _GEN_997; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_999 = 7'h2 == _GEN_108 ? phv_data_2 : _GEN_998; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1000 = 7'h3 == _GEN_108 ? phv_data_3 : _GEN_999; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1001 = 7'h4 == _GEN_108 ? phv_data_4 : _GEN_1000; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1002 = 7'h5 == _GEN_108 ? phv_data_5 : _GEN_1001; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1003 = 7'h6 == _GEN_108 ? phv_data_6 : _GEN_1002; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1004 = 7'h7 == _GEN_108 ? phv_data_7 : _GEN_1003; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1005 = 7'h8 == _GEN_108 ? phv_data_8 : _GEN_1004; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1006 = 7'h9 == _GEN_108 ? phv_data_9 : _GEN_1005; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1007 = 7'ha == _GEN_108 ? phv_data_10 : _GEN_1006; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1008 = 7'hb == _GEN_108 ? phv_data_11 : _GEN_1007; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1009 = 7'hc == _GEN_108 ? phv_data_12 : _GEN_1008; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1010 = 7'hd == _GEN_108 ? phv_data_13 : _GEN_1009; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1011 = 7'he == _GEN_108 ? phv_data_14 : _GEN_1010; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1012 = 7'hf == _GEN_108 ? phv_data_15 : _GEN_1011; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1013 = 7'h10 == _GEN_108 ? phv_data_16 : _GEN_1012; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1014 = 7'h11 == _GEN_108 ? phv_data_17 : _GEN_1013; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1015 = 7'h12 == _GEN_108 ? phv_data_18 : _GEN_1014; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1016 = 7'h13 == _GEN_108 ? phv_data_19 : _GEN_1015; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_5_2 = _GEN_84 ? _GEN_1016 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_1018 = 7'h0 == _GEN_109 ? phv_data_0 : 8'h0; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46 matcher_pisa.scala 120:34]
  wire [7:0] _GEN_1019 = 7'h1 == _GEN_109 ? phv_data_1 : _GEN_1018; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1020 = 7'h2 == _GEN_109 ? phv_data_2 : _GEN_1019; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1021 = 7'h3 == _GEN_109 ? phv_data_3 : _GEN_1020; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1022 = 7'h4 == _GEN_109 ? phv_data_4 : _GEN_1021; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1023 = 7'h5 == _GEN_109 ? phv_data_5 : _GEN_1022; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1024 = 7'h6 == _GEN_109 ? phv_data_6 : _GEN_1023; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1025 = 7'h7 == _GEN_109 ? phv_data_7 : _GEN_1024; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1026 = 7'h8 == _GEN_109 ? phv_data_8 : _GEN_1025; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1027 = 7'h9 == _GEN_109 ? phv_data_9 : _GEN_1026; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1028 = 7'ha == _GEN_109 ? phv_data_10 : _GEN_1027; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1029 = 7'hb == _GEN_109 ? phv_data_11 : _GEN_1028; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1030 = 7'hc == _GEN_109 ? phv_data_12 : _GEN_1029; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1031 = 7'hd == _GEN_109 ? phv_data_13 : _GEN_1030; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1032 = 7'he == _GEN_109 ? phv_data_14 : _GEN_1031; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1033 = 7'hf == _GEN_109 ? phv_data_15 : _GEN_1032; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1034 = 7'h10 == _GEN_109 ? phv_data_16 : _GEN_1033; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1035 = 7'h11 == _GEN_109 ? phv_data_17 : _GEN_1034; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1036 = 7'h12 == _GEN_109 ? phv_data_18 : _GEN_1035; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] _GEN_1037 = 7'h13 == _GEN_109 ? phv_data_19 : _GEN_1036; // @[matcher_pisa.scala 123:62 matcher_pisa.scala 124:46]
  wire [7:0] bytes_5_3 = _GEN_85 ? _GEN_1037 : 8'h0; // @[matcher_pisa.scala 121:46 matcher_pisa.scala 120:34]
  wire [31:0] _groups_5_T = {bytes_5_0,bytes_5_1,bytes_5_2,bytes_5_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1039 = _GEN_61 == 2'h1 ? _groups_5_T : 32'h0; // @[matcher_pisa.scala 115:50 matcher_pisa.scala 129:31 matcher_pisa.scala 114:27]
  wire [15:0] _GEN_1040 = 7'h14 == _GEN_106 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_1041 = 7'h15 == _GEN_106 ? _double_bytes_0_T_1 : _GEN_1040; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1042 = 7'h16 == _GEN_106 ? _double_bytes_0_T_2 : _GEN_1041; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1043 = 7'h17 == _GEN_106 ? _double_bytes_0_T_3 : _GEN_1042; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1044 = 7'h18 == _GEN_106 ? _double_bytes_0_T_4 : _GEN_1043; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1045 = 7'h19 == _GEN_106 ? _double_bytes_0_T_5 : _GEN_1044; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1046 = 7'h1a == _GEN_106 ? _double_bytes_0_T_6 : _GEN_1045; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1047 = 7'h1b == _GEN_106 ? _double_bytes_0_T_7 : _GEN_1046; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1048 = 7'h1c == _GEN_106 ? _double_bytes_0_T_8 : _GEN_1047; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1049 = 7'h1d == _GEN_106 ? _double_bytes_0_T_9 : _GEN_1048; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1050 = 7'h1e == _GEN_106 ? _double_bytes_0_T_10 : _GEN_1049; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1051 = 7'h1f == _GEN_106 ? _double_bytes_0_T_11 : _GEN_1050; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1052 = 7'h20 == _GEN_106 ? _double_bytes_0_T_12 : _GEN_1051; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1053 = 7'h21 == _GEN_106 ? _double_bytes_0_T_13 : _GEN_1052; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1054 = 7'h22 == _GEN_106 ? _double_bytes_0_T_14 : _GEN_1053; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1055 = 7'h23 == _GEN_106 ? _double_bytes_0_T_15 : _GEN_1054; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1056 = 7'h24 == _GEN_106 ? _double_bytes_0_T_16 : _GEN_1055; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1057 = 7'h25 == _GEN_106 ? _double_bytes_0_T_17 : _GEN_1056; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1058 = 7'h26 == _GEN_106 ? _double_bytes_0_T_18 : _GEN_1057; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1059 = 7'h27 == _GEN_106 ? _double_bytes_0_T_19 : _GEN_1058; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1060 = 7'h28 == _GEN_106 ? _double_bytes_0_T_20 : _GEN_1059; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1061 = 7'h29 == _GEN_106 ? _double_bytes_0_T_21 : _GEN_1060; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1062 = 7'h2a == _GEN_106 ? _double_bytes_0_T_22 : _GEN_1061; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1063 = 7'h2b == _GEN_106 ? _double_bytes_0_T_23 : _GEN_1062; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1064 = 7'h2c == _GEN_106 ? _double_bytes_0_T_24 : _GEN_1063; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1065 = 7'h2d == _GEN_106 ? _double_bytes_0_T_25 : _GEN_1064; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1066 = 7'h2e == _GEN_106 ? _double_bytes_0_T_26 : _GEN_1065; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1067 = 7'h2f == _GEN_106 ? _double_bytes_0_T_27 : _GEN_1066; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1068 = 7'h30 == _GEN_106 ? _double_bytes_0_T_28 : _GEN_1067; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1069 = 7'h31 == _GEN_106 ? _double_bytes_0_T_29 : _GEN_1068; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_5_0 = _GEN_82 ? _GEN_1069 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_1071 = 7'h14 == _GEN_107 ? _double_bytes_0_T : 16'h0; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53 matcher_pisa.scala 136:41]
  wire [15:0] _GEN_1072 = 7'h15 == _GEN_107 ? _double_bytes_0_T_1 : _GEN_1071; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1073 = 7'h16 == _GEN_107 ? _double_bytes_0_T_2 : _GEN_1072; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1074 = 7'h17 == _GEN_107 ? _double_bytes_0_T_3 : _GEN_1073; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1075 = 7'h18 == _GEN_107 ? _double_bytes_0_T_4 : _GEN_1074; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1076 = 7'h19 == _GEN_107 ? _double_bytes_0_T_5 : _GEN_1075; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1077 = 7'h1a == _GEN_107 ? _double_bytes_0_T_6 : _GEN_1076; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1078 = 7'h1b == _GEN_107 ? _double_bytes_0_T_7 : _GEN_1077; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1079 = 7'h1c == _GEN_107 ? _double_bytes_0_T_8 : _GEN_1078; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1080 = 7'h1d == _GEN_107 ? _double_bytes_0_T_9 : _GEN_1079; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1081 = 7'h1e == _GEN_107 ? _double_bytes_0_T_10 : _GEN_1080; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1082 = 7'h1f == _GEN_107 ? _double_bytes_0_T_11 : _GEN_1081; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1083 = 7'h20 == _GEN_107 ? _double_bytes_0_T_12 : _GEN_1082; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1084 = 7'h21 == _GEN_107 ? _double_bytes_0_T_13 : _GEN_1083; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1085 = 7'h22 == _GEN_107 ? _double_bytes_0_T_14 : _GEN_1084; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1086 = 7'h23 == _GEN_107 ? _double_bytes_0_T_15 : _GEN_1085; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1087 = 7'h24 == _GEN_107 ? _double_bytes_0_T_16 : _GEN_1086; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1088 = 7'h25 == _GEN_107 ? _double_bytes_0_T_17 : _GEN_1087; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1089 = 7'h26 == _GEN_107 ? _double_bytes_0_T_18 : _GEN_1088; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1090 = 7'h27 == _GEN_107 ? _double_bytes_0_T_19 : _GEN_1089; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1091 = 7'h28 == _GEN_107 ? _double_bytes_0_T_20 : _GEN_1090; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1092 = 7'h29 == _GEN_107 ? _double_bytes_0_T_21 : _GEN_1091; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1093 = 7'h2a == _GEN_107 ? _double_bytes_0_T_22 : _GEN_1092; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1094 = 7'h2b == _GEN_107 ? _double_bytes_0_T_23 : _GEN_1093; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1095 = 7'h2c == _GEN_107 ? _double_bytes_0_T_24 : _GEN_1094; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1096 = 7'h2d == _GEN_107 ? _double_bytes_0_T_25 : _GEN_1095; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1097 = 7'h2e == _GEN_107 ? _double_bytes_0_T_26 : _GEN_1096; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1098 = 7'h2f == _GEN_107 ? _double_bytes_0_T_27 : _GEN_1097; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1099 = 7'h30 == _GEN_107 ? _double_bytes_0_T_28 : _GEN_1098; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] _GEN_1100 = 7'h31 == _GEN_107 ? _double_bytes_0_T_29 : _GEN_1099; // @[matcher_pisa.scala 139:62 matcher_pisa.scala 140:53]
  wire [15:0] double_bytes_5_1 = _GEN_83 ? _GEN_1100 : 16'h0; // @[matcher_pisa.scala 137:46 matcher_pisa.scala 136:41]
  wire [31:0] _groups_5_T_1 = {double_bytes_5_0,double_bytes_5_1}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1102 = _GEN_61 == 2'h2 ? _groups_5_T_1 : _GEN_1039; // @[matcher_pisa.scala 131:50 matcher_pisa.scala 145:31]
  wire [31:0] _GEN_1103 = 7'h32 == _GEN_106 ? _groups_0_T_2 : 32'h0; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39 matcher_pisa.scala 150:31]
  wire [31:0] _GEN_1104 = 7'h33 == _GEN_106 ? _groups_0_T_3 : _GEN_1103; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1105 = 7'h34 == _GEN_106 ? _groups_0_T_4 : _GEN_1104; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1106 = 7'h35 == _GEN_106 ? _groups_0_T_5 : _GEN_1105; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1107 = 7'h36 == _GEN_106 ? _groups_0_T_6 : _GEN_1106; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1108 = 7'h37 == _GEN_106 ? _groups_0_T_7 : _GEN_1107; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1109 = 7'h38 == _GEN_106 ? _groups_0_T_8 : _GEN_1108; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1110 = 7'h39 == _GEN_106 ? _groups_0_T_9 : _GEN_1109; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1111 = 7'h3a == _GEN_106 ? _groups_0_T_10 : _GEN_1110; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1112 = 7'h3b == _GEN_106 ? _groups_0_T_11 : _GEN_1111; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1113 = 7'h3c == _GEN_106 ? _groups_0_T_12 : _GEN_1112; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1114 = 7'h3d == _GEN_106 ? _groups_0_T_13 : _GEN_1113; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1115 = 7'h3e == _GEN_106 ? _groups_0_T_14 : _GEN_1114; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1116 = 7'h3f == _GEN_106 ? _groups_0_T_15 : _GEN_1115; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1117 = 7'h40 == _GEN_106 ? _groups_0_T_16 : _GEN_1116; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1118 = 7'h41 == _GEN_106 ? _groups_0_T_17 : _GEN_1117; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1119 = 7'h42 == _GEN_106 ? _groups_0_T_18 : _GEN_1118; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1120 = 7'h43 == _GEN_106 ? _groups_0_T_19 : _GEN_1119; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1121 = 7'h44 == _GEN_106 ? _groups_0_T_20 : _GEN_1120; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] _GEN_1122 = 7'h45 == _GEN_106 ? _groups_0_T_21 : _GEN_1121; // @[matcher_pisa.scala 152:54 matcher_pisa.scala 153:39]
  wire [31:0] groups_5 = _GEN_61 == 2'h3 ? _GEN_1122 : _GEN_1102; // @[matcher_pisa.scala 147:50]
  wire [191:0] _io_match_key_T = {groups_0,groups_1,groups_2,groups_3,groups_4,groups_5}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[matcher_pisa.scala 104:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[matcher_pisa.scala 104:25]
  assign io_match_key = phv_is_valid_processor ? _io_match_key_T : 192'h0; // @[matcher_pisa.scala 108:39 matcher_pisa.scala 158:26 matcher_pisa.scala 160:26]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[matcher_pisa.scala 103:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[matcher_pisa.scala 103:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[matcher_pisa.scala 103:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[matcher_pisa.scala 103:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[matcher_pisa.scala 103:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[matcher_pisa.scala 103:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[matcher_pisa.scala 103:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[matcher_pisa.scala 103:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[matcher_pisa.scala 103:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[matcher_pisa.scala 103:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[matcher_pisa.scala 103:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[matcher_pisa.scala 103:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[matcher_pisa.scala 103:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[matcher_pisa.scala 103:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[matcher_pisa.scala 103:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[matcher_pisa.scala 103:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[matcher_pisa.scala 103:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[matcher_pisa.scala 103:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[matcher_pisa.scala 103:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[matcher_pisa.scala 103:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[matcher_pisa.scala 103:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[matcher_pisa.scala 103:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[matcher_pisa.scala 103:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[matcher_pisa.scala 103:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[matcher_pisa.scala 103:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[matcher_pisa.scala 103:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[matcher_pisa.scala 103:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[matcher_pisa.scala 103:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[matcher_pisa.scala 103:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[matcher_pisa.scala 103:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[matcher_pisa.scala 103:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[matcher_pisa.scala 103:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[matcher_pisa.scala 103:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[matcher_pisa.scala 103:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[matcher_pisa.scala 103:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[matcher_pisa.scala 103:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[matcher_pisa.scala 103:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[matcher_pisa.scala 103:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[matcher_pisa.scala 103:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[matcher_pisa.scala 103:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[matcher_pisa.scala 103:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[matcher_pisa.scala 103:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[matcher_pisa.scala 103:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[matcher_pisa.scala 103:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[matcher_pisa.scala 103:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[matcher_pisa.scala 103:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[matcher_pisa.scala 103:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[matcher_pisa.scala 103:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[matcher_pisa.scala 103:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[matcher_pisa.scala 103:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[matcher_pisa.scala 103:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[matcher_pisa.scala 103:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[matcher_pisa.scala 103:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[matcher_pisa.scala 103:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[matcher_pisa.scala 103:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[matcher_pisa.scala 103:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[matcher_pisa.scala 103:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[matcher_pisa.scala 103:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[matcher_pisa.scala 103:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[matcher_pisa.scala 103:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[matcher_pisa.scala 103:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[matcher_pisa.scala 103:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[matcher_pisa.scala 103:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[matcher_pisa.scala 103:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[matcher_pisa.scala 103:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[matcher_pisa.scala 103:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[matcher_pisa.scala 103:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[matcher_pisa.scala 103:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[matcher_pisa.scala 103:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[matcher_pisa.scala 103:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[matcher_pisa.scala 103:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[matcher_pisa.scala 103:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[matcher_pisa.scala 103:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[matcher_pisa.scala 103:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[matcher_pisa.scala 103:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[matcher_pisa.scala 103:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[matcher_pisa.scala 103:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[matcher_pisa.scala 103:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[matcher_pisa.scala 103:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[matcher_pisa.scala 103:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[matcher_pisa.scala 103:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[matcher_pisa.scala 103:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[matcher_pisa.scala 103:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[matcher_pisa.scala 103:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[matcher_pisa.scala 103:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[matcher_pisa.scala 103:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[matcher_pisa.scala 103:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[matcher_pisa.scala 103:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[matcher_pisa.scala 103:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[matcher_pisa.scala 103:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[matcher_pisa.scala 103:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[matcher_pisa.scala 103:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[matcher_pisa.scala 103:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[matcher_pisa.scala 103:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[matcher_pisa.scala 103:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[matcher_pisa.scala 103:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[matcher_pisa.scala 103:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[matcher_pisa.scala 103:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[matcher_pisa.scala 103:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[matcher_pisa.scala 103:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[matcher_pisa.scala 103:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[matcher_pisa.scala 103:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[matcher_pisa.scala 103:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[matcher_pisa.scala 103:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[matcher_pisa.scala 103:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[matcher_pisa.scala 103:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[matcher_pisa.scala 103:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[matcher_pisa.scala 103:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[matcher_pisa.scala 103:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[matcher_pisa.scala 103:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[matcher_pisa.scala 103:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[matcher_pisa.scala 103:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[matcher_pisa.scala 103:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[matcher_pisa.scala 103:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[matcher_pisa.scala 103:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[matcher_pisa.scala 103:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[matcher_pisa.scala 103:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[matcher_pisa.scala 103:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[matcher_pisa.scala 103:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[matcher_pisa.scala 103:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[matcher_pisa.scala 103:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[matcher_pisa.scala 103:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[matcher_pisa.scala 103:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[matcher_pisa.scala 103:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[matcher_pisa.scala 103:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[matcher_pisa.scala 103:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[matcher_pisa.scala 103:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[matcher_pisa.scala 103:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[matcher_pisa.scala 103:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[matcher_pisa.scala 103:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[matcher_pisa.scala 103:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[matcher_pisa.scala 103:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[matcher_pisa.scala 103:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[matcher_pisa.scala 103:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[matcher_pisa.scala 103:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[matcher_pisa.scala 103:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[matcher_pisa.scala 103:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[matcher_pisa.scala 103:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[matcher_pisa.scala 103:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[matcher_pisa.scala 103:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[matcher_pisa.scala 103:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[matcher_pisa.scala 103:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[matcher_pisa.scala 103:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[matcher_pisa.scala 103:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[matcher_pisa.scala 103:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[matcher_pisa.scala 103:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[matcher_pisa.scala 103:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[matcher_pisa.scala 103:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[matcher_pisa.scala 103:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[matcher_pisa.scala 103:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[matcher_pisa.scala 103:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[matcher_pisa.scala 103:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[matcher_pisa.scala 103:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[matcher_pisa.scala 103:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[matcher_pisa.scala 103:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[matcher_pisa.scala 103:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[matcher_pisa.scala 103:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[matcher_pisa.scala 103:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[matcher_pisa.scala 103:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[matcher_pisa.scala 103:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[matcher_pisa.scala 103:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[matcher_pisa.scala 103:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_next_config_id = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_161[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
