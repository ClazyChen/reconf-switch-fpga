module Hash(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [1:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [1:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  output        io_pipe_phv_out_is_valid_processor,
  input         io_mod_hash_depth_mod,
  input         io_mod_config_id,
  input  [2:0]  io_mod_hash_depth,
  input  [63:0] io_key_in,
  output [63:0] io_key_out,
  output [7:0]  io_hash_val,
  output [2:0]  io_hash_val_cs
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[hash.scala 101:23]
  wire [1:0] pipe1_io_pipe_phv_in_next_processor_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 101:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 101:23]
  wire [1:0] pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 101:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 101:23]
  wire [63:0] pipe1_io_key_in; // @[hash.scala 101:23]
  wire [63:0] pipe1_io_key_out; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_sum_in; // @[hash.scala 101:23]
  wire [15:0] pipe1_io_sum_out; // @[hash.scala 101:23]
  wire  pipe2_clock; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[hash.scala 102:23]
  wire [1:0] pipe2_io_pipe_phv_in_next_processor_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 102:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 102:23]
  wire [1:0] pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 102:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 102:23]
  wire [63:0] pipe2_io_key_in; // @[hash.scala 102:23]
  wire [63:0] pipe2_io_key_out; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_sum_in; // @[hash.scala 102:23]
  wire [15:0] pipe2_io_sum_out; // @[hash.scala 102:23]
  wire  pipe3_clock; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[hash.scala 103:23]
  wire [1:0] pipe3_io_pipe_phv_in_next_processor_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 103:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 103:23]
  wire [1:0] pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 103:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 103:23]
  wire [63:0] pipe3_io_key_in; // @[hash.scala 103:23]
  wire [63:0] pipe3_io_key_out; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_sum_in; // @[hash.scala 103:23]
  wire [15:0] pipe3_io_sum_out; // @[hash.scala 103:23]
  wire  pipe4_clock; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[hash.scala 104:23]
  wire [1:0] pipe4_io_pipe_phv_in_next_processor_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 104:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 104:23]
  wire [1:0] pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 104:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 104:23]
  wire [2:0] pipe4_io_hash_depth_0; // @[hash.scala 104:23]
  wire [2:0] pipe4_io_hash_depth_1; // @[hash.scala 104:23]
  wire [63:0] pipe4_io_key_in; // @[hash.scala 104:23]
  wire [63:0] pipe4_io_key_out; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_sum_in; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_sum_out; // @[hash.scala 104:23]
  wire [15:0] pipe4_io_val_out; // @[hash.scala 104:23]
  wire  pipe5_clock; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[hash.scala 105:23]
  wire [1:0] pipe5_io_pipe_phv_in_next_processor_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 105:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 105:23]
  wire [1:0] pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 105:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 105:23]
  wire [2:0] pipe5_io_hash_depth_0; // @[hash.scala 105:23]
  wire [2:0] pipe5_io_hash_depth_1; // @[hash.scala 105:23]
  wire [63:0] pipe5_io_key_in; // @[hash.scala 105:23]
  wire [63:0] pipe5_io_key_out; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_sum_in; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_sum_out; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_val_in; // @[hash.scala 105:23]
  wire [15:0] pipe5_io_val_out; // @[hash.scala 105:23]
  wire  pipe6_clock; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[hash.scala 106:23]
  wire [1:0] pipe6_io_pipe_phv_in_next_processor_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 106:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 106:23]
  wire [1:0] pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 106:23]
  wire  pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 106:23]
  wire [2:0] pipe6_io_hash_depth_0; // @[hash.scala 106:23]
  wire [2:0] pipe6_io_hash_depth_1; // @[hash.scala 106:23]
  wire [63:0] pipe6_io_key_in; // @[hash.scala 106:23]
  wire [63:0] pipe6_io_key_out; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_sum_in; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_sum_out; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_val_in; // @[hash.scala 106:23]
  wire [15:0] pipe6_io_val_out; // @[hash.scala 106:23]
  reg [2:0] hash_depth_0; // @[hash.scala 18:26]
  reg [2:0] hash_depth_1; // @[hash.scala 18:26]
  HashSumLevel pipe1 ( // @[hash.scala 101:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe1_io_key_in),
    .io_key_out(pipe1_io_key_out),
    .io_sum_in(pipe1_io_sum_in),
    .io_sum_out(pipe1_io_sum_out)
  );
  HashSumLevel_1 pipe2 ( // @[hash.scala 102:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe2_io_key_in),
    .io_key_out(pipe2_io_key_out),
    .io_sum_in(pipe2_io_sum_in),
    .io_sum_out(pipe2_io_sum_out)
  );
  HashSumLevel_2 pipe3 ( // @[hash.scala 103:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe3_io_key_in),
    .io_key_out(pipe3_io_key_out),
    .io_sum_in(pipe3_io_sum_in),
    .io_sum_out(pipe3_io_sum_out)
  );
  HashReshapeLevel pipe4 ( // @[hash.scala 104:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe4_io_hash_depth_0),
    .io_hash_depth_1(pipe4_io_hash_depth_1),
    .io_key_in(pipe4_io_key_in),
    .io_key_out(pipe4_io_key_out),
    .io_sum_in(pipe4_io_sum_in),
    .io_sum_out(pipe4_io_sum_out),
    .io_val_out(pipe4_io_val_out)
  );
  HashReshapeLevel_1 pipe5 ( // @[hash.scala 105:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe5_io_hash_depth_0),
    .io_hash_depth_1(pipe5_io_hash_depth_1),
    .io_key_in(pipe5_io_key_in),
    .io_key_out(pipe5_io_key_out),
    .io_sum_in(pipe5_io_sum_in),
    .io_sum_out(pipe5_io_sum_out),
    .io_val_in(pipe5_io_val_in),
    .io_val_out(pipe5_io_val_out)
  );
  HashReshapeLevel_2 pipe6 ( // @[hash.scala 106:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe6_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe6_io_hash_depth_0),
    .io_hash_depth_1(pipe6_io_hash_depth_1),
    .io_key_in(pipe6_io_key_in),
    .io_key_out(pipe6_io_key_out),
    .io_sum_in(pipe6_io_sum_in),
    .io_sum_out(pipe6_io_sum_out),
    .io_val_in(pipe6_io_val_in),
    .io_val_out(pipe6_io_val_out)
  );
  assign io_pipe_phv_out_data_0 = pipe6_io_pipe_phv_out_data_0; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_1 = pipe6_io_pipe_phv_out_data_1; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_2 = pipe6_io_pipe_phv_out_data_2; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_3 = pipe6_io_pipe_phv_out_data_3; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_4 = pipe6_io_pipe_phv_out_data_4; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_5 = pipe6_io_pipe_phv_out_data_5; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_6 = pipe6_io_pipe_phv_out_data_6; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_7 = pipe6_io_pipe_phv_out_data_7; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_8 = pipe6_io_pipe_phv_out_data_8; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_9 = pipe6_io_pipe_phv_out_data_9; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_10 = pipe6_io_pipe_phv_out_data_10; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_11 = pipe6_io_pipe_phv_out_data_11; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_12 = pipe6_io_pipe_phv_out_data_12; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_13 = pipe6_io_pipe_phv_out_data_13; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_14 = pipe6_io_pipe_phv_out_data_14; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_15 = pipe6_io_pipe_phv_out_data_15; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_16 = pipe6_io_pipe_phv_out_data_16; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_17 = pipe6_io_pipe_phv_out_data_17; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_18 = pipe6_io_pipe_phv_out_data_18; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_19 = pipe6_io_pipe_phv_out_data_19; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_20 = pipe6_io_pipe_phv_out_data_20; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_21 = pipe6_io_pipe_phv_out_data_21; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_22 = pipe6_io_pipe_phv_out_data_22; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_23 = pipe6_io_pipe_phv_out_data_23; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_24 = pipe6_io_pipe_phv_out_data_24; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_25 = pipe6_io_pipe_phv_out_data_25; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_26 = pipe6_io_pipe_phv_out_data_26; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_27 = pipe6_io_pipe_phv_out_data_27; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_28 = pipe6_io_pipe_phv_out_data_28; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_29 = pipe6_io_pipe_phv_out_data_29; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_30 = pipe6_io_pipe_phv_out_data_30; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_31 = pipe6_io_pipe_phv_out_data_31; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_32 = pipe6_io_pipe_phv_out_data_32; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_33 = pipe6_io_pipe_phv_out_data_33; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_34 = pipe6_io_pipe_phv_out_data_34; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_35 = pipe6_io_pipe_phv_out_data_35; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_36 = pipe6_io_pipe_phv_out_data_36; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_37 = pipe6_io_pipe_phv_out_data_37; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_38 = pipe6_io_pipe_phv_out_data_38; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_39 = pipe6_io_pipe_phv_out_data_39; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_40 = pipe6_io_pipe_phv_out_data_40; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_41 = pipe6_io_pipe_phv_out_data_41; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_42 = pipe6_io_pipe_phv_out_data_42; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_43 = pipe6_io_pipe_phv_out_data_43; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_44 = pipe6_io_pipe_phv_out_data_44; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_45 = pipe6_io_pipe_phv_out_data_45; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_46 = pipe6_io_pipe_phv_out_data_46; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_47 = pipe6_io_pipe_phv_out_data_47; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_48 = pipe6_io_pipe_phv_out_data_48; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_49 = pipe6_io_pipe_phv_out_data_49; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_50 = pipe6_io_pipe_phv_out_data_50; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_51 = pipe6_io_pipe_phv_out_data_51; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_52 = pipe6_io_pipe_phv_out_data_52; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_53 = pipe6_io_pipe_phv_out_data_53; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_54 = pipe6_io_pipe_phv_out_data_54; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_55 = pipe6_io_pipe_phv_out_data_55; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_56 = pipe6_io_pipe_phv_out_data_56; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_57 = pipe6_io_pipe_phv_out_data_57; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_58 = pipe6_io_pipe_phv_out_data_58; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_59 = pipe6_io_pipe_phv_out_data_59; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_60 = pipe6_io_pipe_phv_out_data_60; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_61 = pipe6_io_pipe_phv_out_data_61; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_62 = pipe6_io_pipe_phv_out_data_62; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_63 = pipe6_io_pipe_phv_out_data_63; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_64 = pipe6_io_pipe_phv_out_data_64; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_65 = pipe6_io_pipe_phv_out_data_65; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_66 = pipe6_io_pipe_phv_out_data_66; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_67 = pipe6_io_pipe_phv_out_data_67; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_68 = pipe6_io_pipe_phv_out_data_68; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_69 = pipe6_io_pipe_phv_out_data_69; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_70 = pipe6_io_pipe_phv_out_data_70; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_71 = pipe6_io_pipe_phv_out_data_71; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_72 = pipe6_io_pipe_phv_out_data_72; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_73 = pipe6_io_pipe_phv_out_data_73; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_74 = pipe6_io_pipe_phv_out_data_74; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_75 = pipe6_io_pipe_phv_out_data_75; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_76 = pipe6_io_pipe_phv_out_data_76; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_77 = pipe6_io_pipe_phv_out_data_77; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_78 = pipe6_io_pipe_phv_out_data_78; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_79 = pipe6_io_pipe_phv_out_data_79; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_80 = pipe6_io_pipe_phv_out_data_80; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_81 = pipe6_io_pipe_phv_out_data_81; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_82 = pipe6_io_pipe_phv_out_data_82; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_83 = pipe6_io_pipe_phv_out_data_83; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_84 = pipe6_io_pipe_phv_out_data_84; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_85 = pipe6_io_pipe_phv_out_data_85; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_86 = pipe6_io_pipe_phv_out_data_86; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_87 = pipe6_io_pipe_phv_out_data_87; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_88 = pipe6_io_pipe_phv_out_data_88; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_89 = pipe6_io_pipe_phv_out_data_89; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_90 = pipe6_io_pipe_phv_out_data_90; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_91 = pipe6_io_pipe_phv_out_data_91; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_92 = pipe6_io_pipe_phv_out_data_92; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_93 = pipe6_io_pipe_phv_out_data_93; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_94 = pipe6_io_pipe_phv_out_data_94; // @[hash.scala 138:27]
  assign io_pipe_phv_out_data_95 = pipe6_io_pipe_phv_out_data_95; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_0 = pipe6_io_pipe_phv_out_header_0; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_1 = pipe6_io_pipe_phv_out_header_1; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_2 = pipe6_io_pipe_phv_out_header_2; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_3 = pipe6_io_pipe_phv_out_header_3; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_4 = pipe6_io_pipe_phv_out_header_4; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_5 = pipe6_io_pipe_phv_out_header_5; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_6 = pipe6_io_pipe_phv_out_header_6; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_7 = pipe6_io_pipe_phv_out_header_7; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_8 = pipe6_io_pipe_phv_out_header_8; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_9 = pipe6_io_pipe_phv_out_header_9; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_10 = pipe6_io_pipe_phv_out_header_10; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_11 = pipe6_io_pipe_phv_out_header_11; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_12 = pipe6_io_pipe_phv_out_header_12; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_13 = pipe6_io_pipe_phv_out_header_13; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_14 = pipe6_io_pipe_phv_out_header_14; // @[hash.scala 138:27]
  assign io_pipe_phv_out_header_15 = pipe6_io_pipe_phv_out_header_15; // @[hash.scala 138:27]
  assign io_pipe_phv_out_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 138:27]
  assign io_pipe_phv_out_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 138:27]
  assign io_pipe_phv_out_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 138:27]
  assign io_pipe_phv_out_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 138:27]
  assign io_pipe_phv_out_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 138:27]
  assign io_pipe_phv_out_is_valid_processor = pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 138:27]
  assign io_key_out = pipe6_io_key_out; // @[hash.scala 139:27]
  assign io_hash_val = pipe6_io_sum_out[7:0]; // @[hash.scala 140:46]
  assign io_hash_val_cs = pipe6_io_val_out[7:5]; // @[hash.scala 141:46]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[hash.scala 108:27]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[hash.scala 108:27]
  assign pipe1_io_key_in = io_key_in; // @[hash.scala 109:27]
  assign pipe1_io_sum_in = io_key_in[15:0]; // @[hash.scala 110:39]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 112:27]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 112:27]
  assign pipe2_io_key_in = pipe1_io_key_out; // @[hash.scala 113:27]
  assign pipe2_io_sum_in = pipe1_io_sum_out; // @[hash.scala 114:27]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 116:27]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 116:27]
  assign pipe3_io_key_in = pipe2_io_key_out; // @[hash.scala 117:27]
  assign pipe3_io_sum_in = pipe2_io_sum_out; // @[hash.scala 118:27]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 120:27]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 120:27]
  assign pipe4_io_hash_depth_0 = hash_depth_0; // @[hash.scala 124:27]
  assign pipe4_io_hash_depth_1 = hash_depth_1; // @[hash.scala 124:27]
  assign pipe4_io_key_in = pipe3_io_key_out; // @[hash.scala 121:27]
  assign pipe4_io_sum_in = pipe3_io_sum_out; // @[hash.scala 122:27]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 126:27]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 126:27]
  assign pipe5_io_hash_depth_0 = hash_depth_0; // @[hash.scala 130:27]
  assign pipe5_io_hash_depth_1 = hash_depth_1; // @[hash.scala 130:27]
  assign pipe5_io_key_in = pipe4_io_key_out; // @[hash.scala 127:27]
  assign pipe5_io_sum_in = pipe4_io_sum_out; // @[hash.scala 128:27]
  assign pipe5_io_val_in = pipe4_io_val_out; // @[hash.scala 129:27]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 132:27]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 132:27]
  assign pipe6_io_hash_depth_0 = hash_depth_0; // @[hash.scala 136:27]
  assign pipe6_io_hash_depth_1 = hash_depth_1; // @[hash.scala 136:27]
  assign pipe6_io_key_in = pipe5_io_key_out; // @[hash.scala 133:27]
  assign pipe6_io_sum_in = pipe5_io_sum_out; // @[hash.scala 134:27]
  assign pipe6_io_val_in = pipe5_io_val_out; // @[hash.scala 135:27]
  always @(posedge clock) begin
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (~io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_0 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_1 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hash_depth_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  hash_depth_1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
