module HashSumLevel(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [191:0] io_sum_in,
  output [191:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [191:0] _RAND_183;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 41:22]
  reg [7:0] phv_data_1; // @[hash.scala 41:22]
  reg [7:0] phv_data_2; // @[hash.scala 41:22]
  reg [7:0] phv_data_3; // @[hash.scala 41:22]
  reg [7:0] phv_data_4; // @[hash.scala 41:22]
  reg [7:0] phv_data_5; // @[hash.scala 41:22]
  reg [7:0] phv_data_6; // @[hash.scala 41:22]
  reg [7:0] phv_data_7; // @[hash.scala 41:22]
  reg [7:0] phv_data_8; // @[hash.scala 41:22]
  reg [7:0] phv_data_9; // @[hash.scala 41:22]
  reg [7:0] phv_data_10; // @[hash.scala 41:22]
  reg [7:0] phv_data_11; // @[hash.scala 41:22]
  reg [7:0] phv_data_12; // @[hash.scala 41:22]
  reg [7:0] phv_data_13; // @[hash.scala 41:22]
  reg [7:0] phv_data_14; // @[hash.scala 41:22]
  reg [7:0] phv_data_15; // @[hash.scala 41:22]
  reg [7:0] phv_data_16; // @[hash.scala 41:22]
  reg [7:0] phv_data_17; // @[hash.scala 41:22]
  reg [7:0] phv_data_18; // @[hash.scala 41:22]
  reg [7:0] phv_data_19; // @[hash.scala 41:22]
  reg [7:0] phv_data_20; // @[hash.scala 41:22]
  reg [7:0] phv_data_21; // @[hash.scala 41:22]
  reg [7:0] phv_data_22; // @[hash.scala 41:22]
  reg [7:0] phv_data_23; // @[hash.scala 41:22]
  reg [7:0] phv_data_24; // @[hash.scala 41:22]
  reg [7:0] phv_data_25; // @[hash.scala 41:22]
  reg [7:0] phv_data_26; // @[hash.scala 41:22]
  reg [7:0] phv_data_27; // @[hash.scala 41:22]
  reg [7:0] phv_data_28; // @[hash.scala 41:22]
  reg [7:0] phv_data_29; // @[hash.scala 41:22]
  reg [7:0] phv_data_30; // @[hash.scala 41:22]
  reg [7:0] phv_data_31; // @[hash.scala 41:22]
  reg [7:0] phv_data_32; // @[hash.scala 41:22]
  reg [7:0] phv_data_33; // @[hash.scala 41:22]
  reg [7:0] phv_data_34; // @[hash.scala 41:22]
  reg [7:0] phv_data_35; // @[hash.scala 41:22]
  reg [7:0] phv_data_36; // @[hash.scala 41:22]
  reg [7:0] phv_data_37; // @[hash.scala 41:22]
  reg [7:0] phv_data_38; // @[hash.scala 41:22]
  reg [7:0] phv_data_39; // @[hash.scala 41:22]
  reg [7:0] phv_data_40; // @[hash.scala 41:22]
  reg [7:0] phv_data_41; // @[hash.scala 41:22]
  reg [7:0] phv_data_42; // @[hash.scala 41:22]
  reg [7:0] phv_data_43; // @[hash.scala 41:22]
  reg [7:0] phv_data_44; // @[hash.scala 41:22]
  reg [7:0] phv_data_45; // @[hash.scala 41:22]
  reg [7:0] phv_data_46; // @[hash.scala 41:22]
  reg [7:0] phv_data_47; // @[hash.scala 41:22]
  reg [7:0] phv_data_48; // @[hash.scala 41:22]
  reg [7:0] phv_data_49; // @[hash.scala 41:22]
  reg [7:0] phv_data_50; // @[hash.scala 41:22]
  reg [7:0] phv_data_51; // @[hash.scala 41:22]
  reg [7:0] phv_data_52; // @[hash.scala 41:22]
  reg [7:0] phv_data_53; // @[hash.scala 41:22]
  reg [7:0] phv_data_54; // @[hash.scala 41:22]
  reg [7:0] phv_data_55; // @[hash.scala 41:22]
  reg [7:0] phv_data_56; // @[hash.scala 41:22]
  reg [7:0] phv_data_57; // @[hash.scala 41:22]
  reg [7:0] phv_data_58; // @[hash.scala 41:22]
  reg [7:0] phv_data_59; // @[hash.scala 41:22]
  reg [7:0] phv_data_60; // @[hash.scala 41:22]
  reg [7:0] phv_data_61; // @[hash.scala 41:22]
  reg [7:0] phv_data_62; // @[hash.scala 41:22]
  reg [7:0] phv_data_63; // @[hash.scala 41:22]
  reg [7:0] phv_data_64; // @[hash.scala 41:22]
  reg [7:0] phv_data_65; // @[hash.scala 41:22]
  reg [7:0] phv_data_66; // @[hash.scala 41:22]
  reg [7:0] phv_data_67; // @[hash.scala 41:22]
  reg [7:0] phv_data_68; // @[hash.scala 41:22]
  reg [7:0] phv_data_69; // @[hash.scala 41:22]
  reg [7:0] phv_data_70; // @[hash.scala 41:22]
  reg [7:0] phv_data_71; // @[hash.scala 41:22]
  reg [7:0] phv_data_72; // @[hash.scala 41:22]
  reg [7:0] phv_data_73; // @[hash.scala 41:22]
  reg [7:0] phv_data_74; // @[hash.scala 41:22]
  reg [7:0] phv_data_75; // @[hash.scala 41:22]
  reg [7:0] phv_data_76; // @[hash.scala 41:22]
  reg [7:0] phv_data_77; // @[hash.scala 41:22]
  reg [7:0] phv_data_78; // @[hash.scala 41:22]
  reg [7:0] phv_data_79; // @[hash.scala 41:22]
  reg [7:0] phv_data_80; // @[hash.scala 41:22]
  reg [7:0] phv_data_81; // @[hash.scala 41:22]
  reg [7:0] phv_data_82; // @[hash.scala 41:22]
  reg [7:0] phv_data_83; // @[hash.scala 41:22]
  reg [7:0] phv_data_84; // @[hash.scala 41:22]
  reg [7:0] phv_data_85; // @[hash.scala 41:22]
  reg [7:0] phv_data_86; // @[hash.scala 41:22]
  reg [7:0] phv_data_87; // @[hash.scala 41:22]
  reg [7:0] phv_data_88; // @[hash.scala 41:22]
  reg [7:0] phv_data_89; // @[hash.scala 41:22]
  reg [7:0] phv_data_90; // @[hash.scala 41:22]
  reg [7:0] phv_data_91; // @[hash.scala 41:22]
  reg [7:0] phv_data_92; // @[hash.scala 41:22]
  reg [7:0] phv_data_93; // @[hash.scala 41:22]
  reg [7:0] phv_data_94; // @[hash.scala 41:22]
  reg [7:0] phv_data_95; // @[hash.scala 41:22]
  reg [7:0] phv_data_96; // @[hash.scala 41:22]
  reg [7:0] phv_data_97; // @[hash.scala 41:22]
  reg [7:0] phv_data_98; // @[hash.scala 41:22]
  reg [7:0] phv_data_99; // @[hash.scala 41:22]
  reg [7:0] phv_data_100; // @[hash.scala 41:22]
  reg [7:0] phv_data_101; // @[hash.scala 41:22]
  reg [7:0] phv_data_102; // @[hash.scala 41:22]
  reg [7:0] phv_data_103; // @[hash.scala 41:22]
  reg [7:0] phv_data_104; // @[hash.scala 41:22]
  reg [7:0] phv_data_105; // @[hash.scala 41:22]
  reg [7:0] phv_data_106; // @[hash.scala 41:22]
  reg [7:0] phv_data_107; // @[hash.scala 41:22]
  reg [7:0] phv_data_108; // @[hash.scala 41:22]
  reg [7:0] phv_data_109; // @[hash.scala 41:22]
  reg [7:0] phv_data_110; // @[hash.scala 41:22]
  reg [7:0] phv_data_111; // @[hash.scala 41:22]
  reg [7:0] phv_data_112; // @[hash.scala 41:22]
  reg [7:0] phv_data_113; // @[hash.scala 41:22]
  reg [7:0] phv_data_114; // @[hash.scala 41:22]
  reg [7:0] phv_data_115; // @[hash.scala 41:22]
  reg [7:0] phv_data_116; // @[hash.scala 41:22]
  reg [7:0] phv_data_117; // @[hash.scala 41:22]
  reg [7:0] phv_data_118; // @[hash.scala 41:22]
  reg [7:0] phv_data_119; // @[hash.scala 41:22]
  reg [7:0] phv_data_120; // @[hash.scala 41:22]
  reg [7:0] phv_data_121; // @[hash.scala 41:22]
  reg [7:0] phv_data_122; // @[hash.scala 41:22]
  reg [7:0] phv_data_123; // @[hash.scala 41:22]
  reg [7:0] phv_data_124; // @[hash.scala 41:22]
  reg [7:0] phv_data_125; // @[hash.scala 41:22]
  reg [7:0] phv_data_126; // @[hash.scala 41:22]
  reg [7:0] phv_data_127; // @[hash.scala 41:22]
  reg [7:0] phv_data_128; // @[hash.scala 41:22]
  reg [7:0] phv_data_129; // @[hash.scala 41:22]
  reg [7:0] phv_data_130; // @[hash.scala 41:22]
  reg [7:0] phv_data_131; // @[hash.scala 41:22]
  reg [7:0] phv_data_132; // @[hash.scala 41:22]
  reg [7:0] phv_data_133; // @[hash.scala 41:22]
  reg [7:0] phv_data_134; // @[hash.scala 41:22]
  reg [7:0] phv_data_135; // @[hash.scala 41:22]
  reg [7:0] phv_data_136; // @[hash.scala 41:22]
  reg [7:0] phv_data_137; // @[hash.scala 41:22]
  reg [7:0] phv_data_138; // @[hash.scala 41:22]
  reg [7:0] phv_data_139; // @[hash.scala 41:22]
  reg [7:0] phv_data_140; // @[hash.scala 41:22]
  reg [7:0] phv_data_141; // @[hash.scala 41:22]
  reg [7:0] phv_data_142; // @[hash.scala 41:22]
  reg [7:0] phv_data_143; // @[hash.scala 41:22]
  reg [7:0] phv_data_144; // @[hash.scala 41:22]
  reg [7:0] phv_data_145; // @[hash.scala 41:22]
  reg [7:0] phv_data_146; // @[hash.scala 41:22]
  reg [7:0] phv_data_147; // @[hash.scala 41:22]
  reg [7:0] phv_data_148; // @[hash.scala 41:22]
  reg [7:0] phv_data_149; // @[hash.scala 41:22]
  reg [7:0] phv_data_150; // @[hash.scala 41:22]
  reg [7:0] phv_data_151; // @[hash.scala 41:22]
  reg [7:0] phv_data_152; // @[hash.scala 41:22]
  reg [7:0] phv_data_153; // @[hash.scala 41:22]
  reg [7:0] phv_data_154; // @[hash.scala 41:22]
  reg [7:0] phv_data_155; // @[hash.scala 41:22]
  reg [7:0] phv_data_156; // @[hash.scala 41:22]
  reg [7:0] phv_data_157; // @[hash.scala 41:22]
  reg [7:0] phv_data_158; // @[hash.scala 41:22]
  reg [7:0] phv_data_159; // @[hash.scala 41:22]
  reg [15:0] phv_header_0; // @[hash.scala 41:22]
  reg [15:0] phv_header_1; // @[hash.scala 41:22]
  reg [15:0] phv_header_2; // @[hash.scala 41:22]
  reg [15:0] phv_header_3; // @[hash.scala 41:22]
  reg [15:0] phv_header_4; // @[hash.scala 41:22]
  reg [15:0] phv_header_5; // @[hash.scala 41:22]
  reg [15:0] phv_header_6; // @[hash.scala 41:22]
  reg [15:0] phv_header_7; // @[hash.scala 41:22]
  reg [15:0] phv_header_8; // @[hash.scala 41:22]
  reg [15:0] phv_header_9; // @[hash.scala 41:22]
  reg [15:0] phv_header_10; // @[hash.scala 41:22]
  reg [15:0] phv_header_11; // @[hash.scala 41:22]
  reg [15:0] phv_header_12; // @[hash.scala 41:22]
  reg [15:0] phv_header_13; // @[hash.scala 41:22]
  reg [15:0] phv_header_14; // @[hash.scala 41:22]
  reg [15:0] phv_header_15; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 41:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 41:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 41:22]
  reg  phv_next_config_id; // @[hash.scala 41:22]
  reg  phv_is_valid_processor; // @[hash.scala 41:22]
  reg [191:0] key; // @[hash.scala 45:22]
  reg [191:0] sum; // @[hash.scala 49:22]
  wire [15:0] sum_temp_0 = sum[191:176]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_1 = sum[175:160]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_2 = sum[159:144]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_3 = sum[143:128]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_4 = sum[127:112]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_5 = sum[111:96]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_6 = sum[95:80]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_7 = sum[79:64]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_8 = sum[63:48]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_9 = sum[47:32]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_10 = sum[31:16]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_11 = sum[15:0]; // @[hash.scala 64:35]
  wire [15:0] out_temp_0 = sum_temp_0 + sum_temp_1; // @[hash.scala 70:51]
  wire [15:0] out_temp_1 = sum_temp_2 + sum_temp_3; // @[hash.scala 70:51]
  wire [15:0] out_temp_2 = sum_temp_4 + sum_temp_5; // @[hash.scala 70:51]
  wire [15:0] out_temp_3 = sum_temp_6 + sum_temp_7; // @[hash.scala 70:51]
  wire [15:0] out_temp_4 = sum_temp_8 + sum_temp_9; // @[hash.scala 70:51]
  wire [15:0] out_temp_5 = sum_temp_10 + sum_temp_11; // @[hash.scala 70:51]
  wire [95:0] _io_sum_out_T = {out_temp_0,out_temp_1,out_temp_2,out_temp_3,out_temp_4,out_temp_5}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 43:25]
  assign io_key_out = key; // @[hash.scala 47:20]
  assign io_sum_out = phv_is_valid_processor ? {{96'd0}, _io_sum_out_T} : sum; // @[hash.scala 52:39 hash.scala 75:24 hash.scala 77:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 42:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 42:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 42:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 42:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 42:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 42:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 42:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 42:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 42:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 42:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 42:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 42:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 42:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 42:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 42:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 42:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 42:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 42:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 42:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 42:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 42:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 42:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 42:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 42:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 42:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 42:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 42:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 42:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 42:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 42:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 42:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 42:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 42:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 42:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 42:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 42:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 42:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 42:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 42:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 42:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 42:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 42:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 42:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 42:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 42:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 42:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 42:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 42:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 42:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 42:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 42:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 42:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 42:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 42:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 42:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 42:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 42:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 42:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 42:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 42:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 42:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 42:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 42:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 42:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 42:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 42:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 42:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 42:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 42:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 42:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 42:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 42:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 42:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 42:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 42:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 42:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 42:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 42:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 42:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 42:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 42:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 42:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 42:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 42:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 42:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 42:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 42:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 42:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 42:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 42:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 42:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 42:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 42:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 42:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 42:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 42:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 42:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 42:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 42:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 42:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 42:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 42:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 42:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 42:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 42:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 42:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 42:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 42:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 42:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 42:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 42:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 42:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 42:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 42:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 42:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 42:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 42:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 42:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 42:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 42:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 42:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 42:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 42:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 42:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 42:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 42:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 42:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 42:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 42:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 42:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 42:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 42:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 42:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 42:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 42:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 42:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 42:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 42:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 42:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 42:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 42:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 42:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 42:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 42:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 42:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 42:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 42:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 42:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 42:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 42:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 42:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 42:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 42:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 42:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 42:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 42:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 42:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 42:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 42:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 42:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 42:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 42:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 42:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 42:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 42:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 42:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 42:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 42:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 42:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 42:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 42:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 42:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 42:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 42:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 42:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 42:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 42:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 42:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 42:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 42:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 42:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 42:13]
    key <= io_key_in; // @[hash.scala 46:13]
    sum <= io_sum_in; // @[hash.scala 50:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {6{`RANDOM}};
  sum = _RAND_183[191:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashSumLevel_1(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [191:0] io_sum_in,
  output [191:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [191:0] _RAND_183;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 41:22]
  reg [7:0] phv_data_1; // @[hash.scala 41:22]
  reg [7:0] phv_data_2; // @[hash.scala 41:22]
  reg [7:0] phv_data_3; // @[hash.scala 41:22]
  reg [7:0] phv_data_4; // @[hash.scala 41:22]
  reg [7:0] phv_data_5; // @[hash.scala 41:22]
  reg [7:0] phv_data_6; // @[hash.scala 41:22]
  reg [7:0] phv_data_7; // @[hash.scala 41:22]
  reg [7:0] phv_data_8; // @[hash.scala 41:22]
  reg [7:0] phv_data_9; // @[hash.scala 41:22]
  reg [7:0] phv_data_10; // @[hash.scala 41:22]
  reg [7:0] phv_data_11; // @[hash.scala 41:22]
  reg [7:0] phv_data_12; // @[hash.scala 41:22]
  reg [7:0] phv_data_13; // @[hash.scala 41:22]
  reg [7:0] phv_data_14; // @[hash.scala 41:22]
  reg [7:0] phv_data_15; // @[hash.scala 41:22]
  reg [7:0] phv_data_16; // @[hash.scala 41:22]
  reg [7:0] phv_data_17; // @[hash.scala 41:22]
  reg [7:0] phv_data_18; // @[hash.scala 41:22]
  reg [7:0] phv_data_19; // @[hash.scala 41:22]
  reg [7:0] phv_data_20; // @[hash.scala 41:22]
  reg [7:0] phv_data_21; // @[hash.scala 41:22]
  reg [7:0] phv_data_22; // @[hash.scala 41:22]
  reg [7:0] phv_data_23; // @[hash.scala 41:22]
  reg [7:0] phv_data_24; // @[hash.scala 41:22]
  reg [7:0] phv_data_25; // @[hash.scala 41:22]
  reg [7:0] phv_data_26; // @[hash.scala 41:22]
  reg [7:0] phv_data_27; // @[hash.scala 41:22]
  reg [7:0] phv_data_28; // @[hash.scala 41:22]
  reg [7:0] phv_data_29; // @[hash.scala 41:22]
  reg [7:0] phv_data_30; // @[hash.scala 41:22]
  reg [7:0] phv_data_31; // @[hash.scala 41:22]
  reg [7:0] phv_data_32; // @[hash.scala 41:22]
  reg [7:0] phv_data_33; // @[hash.scala 41:22]
  reg [7:0] phv_data_34; // @[hash.scala 41:22]
  reg [7:0] phv_data_35; // @[hash.scala 41:22]
  reg [7:0] phv_data_36; // @[hash.scala 41:22]
  reg [7:0] phv_data_37; // @[hash.scala 41:22]
  reg [7:0] phv_data_38; // @[hash.scala 41:22]
  reg [7:0] phv_data_39; // @[hash.scala 41:22]
  reg [7:0] phv_data_40; // @[hash.scala 41:22]
  reg [7:0] phv_data_41; // @[hash.scala 41:22]
  reg [7:0] phv_data_42; // @[hash.scala 41:22]
  reg [7:0] phv_data_43; // @[hash.scala 41:22]
  reg [7:0] phv_data_44; // @[hash.scala 41:22]
  reg [7:0] phv_data_45; // @[hash.scala 41:22]
  reg [7:0] phv_data_46; // @[hash.scala 41:22]
  reg [7:0] phv_data_47; // @[hash.scala 41:22]
  reg [7:0] phv_data_48; // @[hash.scala 41:22]
  reg [7:0] phv_data_49; // @[hash.scala 41:22]
  reg [7:0] phv_data_50; // @[hash.scala 41:22]
  reg [7:0] phv_data_51; // @[hash.scala 41:22]
  reg [7:0] phv_data_52; // @[hash.scala 41:22]
  reg [7:0] phv_data_53; // @[hash.scala 41:22]
  reg [7:0] phv_data_54; // @[hash.scala 41:22]
  reg [7:0] phv_data_55; // @[hash.scala 41:22]
  reg [7:0] phv_data_56; // @[hash.scala 41:22]
  reg [7:0] phv_data_57; // @[hash.scala 41:22]
  reg [7:0] phv_data_58; // @[hash.scala 41:22]
  reg [7:0] phv_data_59; // @[hash.scala 41:22]
  reg [7:0] phv_data_60; // @[hash.scala 41:22]
  reg [7:0] phv_data_61; // @[hash.scala 41:22]
  reg [7:0] phv_data_62; // @[hash.scala 41:22]
  reg [7:0] phv_data_63; // @[hash.scala 41:22]
  reg [7:0] phv_data_64; // @[hash.scala 41:22]
  reg [7:0] phv_data_65; // @[hash.scala 41:22]
  reg [7:0] phv_data_66; // @[hash.scala 41:22]
  reg [7:0] phv_data_67; // @[hash.scala 41:22]
  reg [7:0] phv_data_68; // @[hash.scala 41:22]
  reg [7:0] phv_data_69; // @[hash.scala 41:22]
  reg [7:0] phv_data_70; // @[hash.scala 41:22]
  reg [7:0] phv_data_71; // @[hash.scala 41:22]
  reg [7:0] phv_data_72; // @[hash.scala 41:22]
  reg [7:0] phv_data_73; // @[hash.scala 41:22]
  reg [7:0] phv_data_74; // @[hash.scala 41:22]
  reg [7:0] phv_data_75; // @[hash.scala 41:22]
  reg [7:0] phv_data_76; // @[hash.scala 41:22]
  reg [7:0] phv_data_77; // @[hash.scala 41:22]
  reg [7:0] phv_data_78; // @[hash.scala 41:22]
  reg [7:0] phv_data_79; // @[hash.scala 41:22]
  reg [7:0] phv_data_80; // @[hash.scala 41:22]
  reg [7:0] phv_data_81; // @[hash.scala 41:22]
  reg [7:0] phv_data_82; // @[hash.scala 41:22]
  reg [7:0] phv_data_83; // @[hash.scala 41:22]
  reg [7:0] phv_data_84; // @[hash.scala 41:22]
  reg [7:0] phv_data_85; // @[hash.scala 41:22]
  reg [7:0] phv_data_86; // @[hash.scala 41:22]
  reg [7:0] phv_data_87; // @[hash.scala 41:22]
  reg [7:0] phv_data_88; // @[hash.scala 41:22]
  reg [7:0] phv_data_89; // @[hash.scala 41:22]
  reg [7:0] phv_data_90; // @[hash.scala 41:22]
  reg [7:0] phv_data_91; // @[hash.scala 41:22]
  reg [7:0] phv_data_92; // @[hash.scala 41:22]
  reg [7:0] phv_data_93; // @[hash.scala 41:22]
  reg [7:0] phv_data_94; // @[hash.scala 41:22]
  reg [7:0] phv_data_95; // @[hash.scala 41:22]
  reg [7:0] phv_data_96; // @[hash.scala 41:22]
  reg [7:0] phv_data_97; // @[hash.scala 41:22]
  reg [7:0] phv_data_98; // @[hash.scala 41:22]
  reg [7:0] phv_data_99; // @[hash.scala 41:22]
  reg [7:0] phv_data_100; // @[hash.scala 41:22]
  reg [7:0] phv_data_101; // @[hash.scala 41:22]
  reg [7:0] phv_data_102; // @[hash.scala 41:22]
  reg [7:0] phv_data_103; // @[hash.scala 41:22]
  reg [7:0] phv_data_104; // @[hash.scala 41:22]
  reg [7:0] phv_data_105; // @[hash.scala 41:22]
  reg [7:0] phv_data_106; // @[hash.scala 41:22]
  reg [7:0] phv_data_107; // @[hash.scala 41:22]
  reg [7:0] phv_data_108; // @[hash.scala 41:22]
  reg [7:0] phv_data_109; // @[hash.scala 41:22]
  reg [7:0] phv_data_110; // @[hash.scala 41:22]
  reg [7:0] phv_data_111; // @[hash.scala 41:22]
  reg [7:0] phv_data_112; // @[hash.scala 41:22]
  reg [7:0] phv_data_113; // @[hash.scala 41:22]
  reg [7:0] phv_data_114; // @[hash.scala 41:22]
  reg [7:0] phv_data_115; // @[hash.scala 41:22]
  reg [7:0] phv_data_116; // @[hash.scala 41:22]
  reg [7:0] phv_data_117; // @[hash.scala 41:22]
  reg [7:0] phv_data_118; // @[hash.scala 41:22]
  reg [7:0] phv_data_119; // @[hash.scala 41:22]
  reg [7:0] phv_data_120; // @[hash.scala 41:22]
  reg [7:0] phv_data_121; // @[hash.scala 41:22]
  reg [7:0] phv_data_122; // @[hash.scala 41:22]
  reg [7:0] phv_data_123; // @[hash.scala 41:22]
  reg [7:0] phv_data_124; // @[hash.scala 41:22]
  reg [7:0] phv_data_125; // @[hash.scala 41:22]
  reg [7:0] phv_data_126; // @[hash.scala 41:22]
  reg [7:0] phv_data_127; // @[hash.scala 41:22]
  reg [7:0] phv_data_128; // @[hash.scala 41:22]
  reg [7:0] phv_data_129; // @[hash.scala 41:22]
  reg [7:0] phv_data_130; // @[hash.scala 41:22]
  reg [7:0] phv_data_131; // @[hash.scala 41:22]
  reg [7:0] phv_data_132; // @[hash.scala 41:22]
  reg [7:0] phv_data_133; // @[hash.scala 41:22]
  reg [7:0] phv_data_134; // @[hash.scala 41:22]
  reg [7:0] phv_data_135; // @[hash.scala 41:22]
  reg [7:0] phv_data_136; // @[hash.scala 41:22]
  reg [7:0] phv_data_137; // @[hash.scala 41:22]
  reg [7:0] phv_data_138; // @[hash.scala 41:22]
  reg [7:0] phv_data_139; // @[hash.scala 41:22]
  reg [7:0] phv_data_140; // @[hash.scala 41:22]
  reg [7:0] phv_data_141; // @[hash.scala 41:22]
  reg [7:0] phv_data_142; // @[hash.scala 41:22]
  reg [7:0] phv_data_143; // @[hash.scala 41:22]
  reg [7:0] phv_data_144; // @[hash.scala 41:22]
  reg [7:0] phv_data_145; // @[hash.scala 41:22]
  reg [7:0] phv_data_146; // @[hash.scala 41:22]
  reg [7:0] phv_data_147; // @[hash.scala 41:22]
  reg [7:0] phv_data_148; // @[hash.scala 41:22]
  reg [7:0] phv_data_149; // @[hash.scala 41:22]
  reg [7:0] phv_data_150; // @[hash.scala 41:22]
  reg [7:0] phv_data_151; // @[hash.scala 41:22]
  reg [7:0] phv_data_152; // @[hash.scala 41:22]
  reg [7:0] phv_data_153; // @[hash.scala 41:22]
  reg [7:0] phv_data_154; // @[hash.scala 41:22]
  reg [7:0] phv_data_155; // @[hash.scala 41:22]
  reg [7:0] phv_data_156; // @[hash.scala 41:22]
  reg [7:0] phv_data_157; // @[hash.scala 41:22]
  reg [7:0] phv_data_158; // @[hash.scala 41:22]
  reg [7:0] phv_data_159; // @[hash.scala 41:22]
  reg [15:0] phv_header_0; // @[hash.scala 41:22]
  reg [15:0] phv_header_1; // @[hash.scala 41:22]
  reg [15:0] phv_header_2; // @[hash.scala 41:22]
  reg [15:0] phv_header_3; // @[hash.scala 41:22]
  reg [15:0] phv_header_4; // @[hash.scala 41:22]
  reg [15:0] phv_header_5; // @[hash.scala 41:22]
  reg [15:0] phv_header_6; // @[hash.scala 41:22]
  reg [15:0] phv_header_7; // @[hash.scala 41:22]
  reg [15:0] phv_header_8; // @[hash.scala 41:22]
  reg [15:0] phv_header_9; // @[hash.scala 41:22]
  reg [15:0] phv_header_10; // @[hash.scala 41:22]
  reg [15:0] phv_header_11; // @[hash.scala 41:22]
  reg [15:0] phv_header_12; // @[hash.scala 41:22]
  reg [15:0] phv_header_13; // @[hash.scala 41:22]
  reg [15:0] phv_header_14; // @[hash.scala 41:22]
  reg [15:0] phv_header_15; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 41:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 41:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 41:22]
  reg  phv_next_config_id; // @[hash.scala 41:22]
  reg  phv_is_valid_processor; // @[hash.scala 41:22]
  reg [191:0] key; // @[hash.scala 45:22]
  reg [191:0] sum; // @[hash.scala 49:22]
  wire [15:0] sum_temp_0 = sum[191:176]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_1 = sum[175:160]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_2 = sum[159:144]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_3 = sum[143:128]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_4 = sum[127:112]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_5 = sum[111:96]; // @[hash.scala 64:35]
  wire [15:0] out_temp_0 = sum_temp_0 + sum_temp_1; // @[hash.scala 70:51]
  wire [15:0] out_temp_1 = sum_temp_2 + sum_temp_3; // @[hash.scala 70:51]
  wire [15:0] out_temp_2 = sum_temp_4 + sum_temp_5; // @[hash.scala 70:51]
  wire [47:0] _io_sum_out_T = {out_temp_0,out_temp_1,out_temp_2}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 43:25]
  assign io_key_out = key; // @[hash.scala 47:20]
  assign io_sum_out = phv_is_valid_processor ? {{144'd0}, _io_sum_out_T} : sum; // @[hash.scala 52:39 hash.scala 75:24 hash.scala 77:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 42:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 42:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 42:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 42:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 42:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 42:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 42:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 42:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 42:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 42:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 42:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 42:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 42:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 42:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 42:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 42:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 42:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 42:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 42:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 42:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 42:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 42:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 42:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 42:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 42:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 42:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 42:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 42:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 42:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 42:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 42:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 42:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 42:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 42:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 42:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 42:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 42:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 42:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 42:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 42:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 42:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 42:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 42:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 42:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 42:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 42:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 42:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 42:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 42:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 42:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 42:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 42:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 42:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 42:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 42:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 42:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 42:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 42:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 42:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 42:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 42:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 42:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 42:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 42:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 42:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 42:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 42:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 42:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 42:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 42:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 42:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 42:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 42:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 42:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 42:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 42:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 42:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 42:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 42:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 42:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 42:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 42:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 42:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 42:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 42:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 42:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 42:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 42:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 42:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 42:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 42:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 42:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 42:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 42:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 42:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 42:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 42:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 42:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 42:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 42:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 42:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 42:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 42:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 42:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 42:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 42:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 42:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 42:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 42:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 42:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 42:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 42:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 42:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 42:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 42:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 42:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 42:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 42:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 42:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 42:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 42:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 42:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 42:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 42:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 42:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 42:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 42:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 42:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 42:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 42:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 42:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 42:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 42:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 42:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 42:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 42:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 42:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 42:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 42:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 42:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 42:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 42:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 42:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 42:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 42:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 42:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 42:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 42:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 42:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 42:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 42:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 42:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 42:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 42:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 42:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 42:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 42:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 42:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 42:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 42:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 42:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 42:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 42:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 42:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 42:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 42:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 42:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 42:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 42:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 42:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 42:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 42:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 42:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 42:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 42:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 42:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 42:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 42:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 42:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 42:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 42:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 42:13]
    key <= io_key_in; // @[hash.scala 46:13]
    sum <= io_sum_in; // @[hash.scala 50:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {6{`RANDOM}};
  sum = _RAND_183[191:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashSumLevel_2(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [191:0] io_sum_in,
  output [191:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [191:0] _RAND_183;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 41:22]
  reg [7:0] phv_data_1; // @[hash.scala 41:22]
  reg [7:0] phv_data_2; // @[hash.scala 41:22]
  reg [7:0] phv_data_3; // @[hash.scala 41:22]
  reg [7:0] phv_data_4; // @[hash.scala 41:22]
  reg [7:0] phv_data_5; // @[hash.scala 41:22]
  reg [7:0] phv_data_6; // @[hash.scala 41:22]
  reg [7:0] phv_data_7; // @[hash.scala 41:22]
  reg [7:0] phv_data_8; // @[hash.scala 41:22]
  reg [7:0] phv_data_9; // @[hash.scala 41:22]
  reg [7:0] phv_data_10; // @[hash.scala 41:22]
  reg [7:0] phv_data_11; // @[hash.scala 41:22]
  reg [7:0] phv_data_12; // @[hash.scala 41:22]
  reg [7:0] phv_data_13; // @[hash.scala 41:22]
  reg [7:0] phv_data_14; // @[hash.scala 41:22]
  reg [7:0] phv_data_15; // @[hash.scala 41:22]
  reg [7:0] phv_data_16; // @[hash.scala 41:22]
  reg [7:0] phv_data_17; // @[hash.scala 41:22]
  reg [7:0] phv_data_18; // @[hash.scala 41:22]
  reg [7:0] phv_data_19; // @[hash.scala 41:22]
  reg [7:0] phv_data_20; // @[hash.scala 41:22]
  reg [7:0] phv_data_21; // @[hash.scala 41:22]
  reg [7:0] phv_data_22; // @[hash.scala 41:22]
  reg [7:0] phv_data_23; // @[hash.scala 41:22]
  reg [7:0] phv_data_24; // @[hash.scala 41:22]
  reg [7:0] phv_data_25; // @[hash.scala 41:22]
  reg [7:0] phv_data_26; // @[hash.scala 41:22]
  reg [7:0] phv_data_27; // @[hash.scala 41:22]
  reg [7:0] phv_data_28; // @[hash.scala 41:22]
  reg [7:0] phv_data_29; // @[hash.scala 41:22]
  reg [7:0] phv_data_30; // @[hash.scala 41:22]
  reg [7:0] phv_data_31; // @[hash.scala 41:22]
  reg [7:0] phv_data_32; // @[hash.scala 41:22]
  reg [7:0] phv_data_33; // @[hash.scala 41:22]
  reg [7:0] phv_data_34; // @[hash.scala 41:22]
  reg [7:0] phv_data_35; // @[hash.scala 41:22]
  reg [7:0] phv_data_36; // @[hash.scala 41:22]
  reg [7:0] phv_data_37; // @[hash.scala 41:22]
  reg [7:0] phv_data_38; // @[hash.scala 41:22]
  reg [7:0] phv_data_39; // @[hash.scala 41:22]
  reg [7:0] phv_data_40; // @[hash.scala 41:22]
  reg [7:0] phv_data_41; // @[hash.scala 41:22]
  reg [7:0] phv_data_42; // @[hash.scala 41:22]
  reg [7:0] phv_data_43; // @[hash.scala 41:22]
  reg [7:0] phv_data_44; // @[hash.scala 41:22]
  reg [7:0] phv_data_45; // @[hash.scala 41:22]
  reg [7:0] phv_data_46; // @[hash.scala 41:22]
  reg [7:0] phv_data_47; // @[hash.scala 41:22]
  reg [7:0] phv_data_48; // @[hash.scala 41:22]
  reg [7:0] phv_data_49; // @[hash.scala 41:22]
  reg [7:0] phv_data_50; // @[hash.scala 41:22]
  reg [7:0] phv_data_51; // @[hash.scala 41:22]
  reg [7:0] phv_data_52; // @[hash.scala 41:22]
  reg [7:0] phv_data_53; // @[hash.scala 41:22]
  reg [7:0] phv_data_54; // @[hash.scala 41:22]
  reg [7:0] phv_data_55; // @[hash.scala 41:22]
  reg [7:0] phv_data_56; // @[hash.scala 41:22]
  reg [7:0] phv_data_57; // @[hash.scala 41:22]
  reg [7:0] phv_data_58; // @[hash.scala 41:22]
  reg [7:0] phv_data_59; // @[hash.scala 41:22]
  reg [7:0] phv_data_60; // @[hash.scala 41:22]
  reg [7:0] phv_data_61; // @[hash.scala 41:22]
  reg [7:0] phv_data_62; // @[hash.scala 41:22]
  reg [7:0] phv_data_63; // @[hash.scala 41:22]
  reg [7:0] phv_data_64; // @[hash.scala 41:22]
  reg [7:0] phv_data_65; // @[hash.scala 41:22]
  reg [7:0] phv_data_66; // @[hash.scala 41:22]
  reg [7:0] phv_data_67; // @[hash.scala 41:22]
  reg [7:0] phv_data_68; // @[hash.scala 41:22]
  reg [7:0] phv_data_69; // @[hash.scala 41:22]
  reg [7:0] phv_data_70; // @[hash.scala 41:22]
  reg [7:0] phv_data_71; // @[hash.scala 41:22]
  reg [7:0] phv_data_72; // @[hash.scala 41:22]
  reg [7:0] phv_data_73; // @[hash.scala 41:22]
  reg [7:0] phv_data_74; // @[hash.scala 41:22]
  reg [7:0] phv_data_75; // @[hash.scala 41:22]
  reg [7:0] phv_data_76; // @[hash.scala 41:22]
  reg [7:0] phv_data_77; // @[hash.scala 41:22]
  reg [7:0] phv_data_78; // @[hash.scala 41:22]
  reg [7:0] phv_data_79; // @[hash.scala 41:22]
  reg [7:0] phv_data_80; // @[hash.scala 41:22]
  reg [7:0] phv_data_81; // @[hash.scala 41:22]
  reg [7:0] phv_data_82; // @[hash.scala 41:22]
  reg [7:0] phv_data_83; // @[hash.scala 41:22]
  reg [7:0] phv_data_84; // @[hash.scala 41:22]
  reg [7:0] phv_data_85; // @[hash.scala 41:22]
  reg [7:0] phv_data_86; // @[hash.scala 41:22]
  reg [7:0] phv_data_87; // @[hash.scala 41:22]
  reg [7:0] phv_data_88; // @[hash.scala 41:22]
  reg [7:0] phv_data_89; // @[hash.scala 41:22]
  reg [7:0] phv_data_90; // @[hash.scala 41:22]
  reg [7:0] phv_data_91; // @[hash.scala 41:22]
  reg [7:0] phv_data_92; // @[hash.scala 41:22]
  reg [7:0] phv_data_93; // @[hash.scala 41:22]
  reg [7:0] phv_data_94; // @[hash.scala 41:22]
  reg [7:0] phv_data_95; // @[hash.scala 41:22]
  reg [7:0] phv_data_96; // @[hash.scala 41:22]
  reg [7:0] phv_data_97; // @[hash.scala 41:22]
  reg [7:0] phv_data_98; // @[hash.scala 41:22]
  reg [7:0] phv_data_99; // @[hash.scala 41:22]
  reg [7:0] phv_data_100; // @[hash.scala 41:22]
  reg [7:0] phv_data_101; // @[hash.scala 41:22]
  reg [7:0] phv_data_102; // @[hash.scala 41:22]
  reg [7:0] phv_data_103; // @[hash.scala 41:22]
  reg [7:0] phv_data_104; // @[hash.scala 41:22]
  reg [7:0] phv_data_105; // @[hash.scala 41:22]
  reg [7:0] phv_data_106; // @[hash.scala 41:22]
  reg [7:0] phv_data_107; // @[hash.scala 41:22]
  reg [7:0] phv_data_108; // @[hash.scala 41:22]
  reg [7:0] phv_data_109; // @[hash.scala 41:22]
  reg [7:0] phv_data_110; // @[hash.scala 41:22]
  reg [7:0] phv_data_111; // @[hash.scala 41:22]
  reg [7:0] phv_data_112; // @[hash.scala 41:22]
  reg [7:0] phv_data_113; // @[hash.scala 41:22]
  reg [7:0] phv_data_114; // @[hash.scala 41:22]
  reg [7:0] phv_data_115; // @[hash.scala 41:22]
  reg [7:0] phv_data_116; // @[hash.scala 41:22]
  reg [7:0] phv_data_117; // @[hash.scala 41:22]
  reg [7:0] phv_data_118; // @[hash.scala 41:22]
  reg [7:0] phv_data_119; // @[hash.scala 41:22]
  reg [7:0] phv_data_120; // @[hash.scala 41:22]
  reg [7:0] phv_data_121; // @[hash.scala 41:22]
  reg [7:0] phv_data_122; // @[hash.scala 41:22]
  reg [7:0] phv_data_123; // @[hash.scala 41:22]
  reg [7:0] phv_data_124; // @[hash.scala 41:22]
  reg [7:0] phv_data_125; // @[hash.scala 41:22]
  reg [7:0] phv_data_126; // @[hash.scala 41:22]
  reg [7:0] phv_data_127; // @[hash.scala 41:22]
  reg [7:0] phv_data_128; // @[hash.scala 41:22]
  reg [7:0] phv_data_129; // @[hash.scala 41:22]
  reg [7:0] phv_data_130; // @[hash.scala 41:22]
  reg [7:0] phv_data_131; // @[hash.scala 41:22]
  reg [7:0] phv_data_132; // @[hash.scala 41:22]
  reg [7:0] phv_data_133; // @[hash.scala 41:22]
  reg [7:0] phv_data_134; // @[hash.scala 41:22]
  reg [7:0] phv_data_135; // @[hash.scala 41:22]
  reg [7:0] phv_data_136; // @[hash.scala 41:22]
  reg [7:0] phv_data_137; // @[hash.scala 41:22]
  reg [7:0] phv_data_138; // @[hash.scala 41:22]
  reg [7:0] phv_data_139; // @[hash.scala 41:22]
  reg [7:0] phv_data_140; // @[hash.scala 41:22]
  reg [7:0] phv_data_141; // @[hash.scala 41:22]
  reg [7:0] phv_data_142; // @[hash.scala 41:22]
  reg [7:0] phv_data_143; // @[hash.scala 41:22]
  reg [7:0] phv_data_144; // @[hash.scala 41:22]
  reg [7:0] phv_data_145; // @[hash.scala 41:22]
  reg [7:0] phv_data_146; // @[hash.scala 41:22]
  reg [7:0] phv_data_147; // @[hash.scala 41:22]
  reg [7:0] phv_data_148; // @[hash.scala 41:22]
  reg [7:0] phv_data_149; // @[hash.scala 41:22]
  reg [7:0] phv_data_150; // @[hash.scala 41:22]
  reg [7:0] phv_data_151; // @[hash.scala 41:22]
  reg [7:0] phv_data_152; // @[hash.scala 41:22]
  reg [7:0] phv_data_153; // @[hash.scala 41:22]
  reg [7:0] phv_data_154; // @[hash.scala 41:22]
  reg [7:0] phv_data_155; // @[hash.scala 41:22]
  reg [7:0] phv_data_156; // @[hash.scala 41:22]
  reg [7:0] phv_data_157; // @[hash.scala 41:22]
  reg [7:0] phv_data_158; // @[hash.scala 41:22]
  reg [7:0] phv_data_159; // @[hash.scala 41:22]
  reg [15:0] phv_header_0; // @[hash.scala 41:22]
  reg [15:0] phv_header_1; // @[hash.scala 41:22]
  reg [15:0] phv_header_2; // @[hash.scala 41:22]
  reg [15:0] phv_header_3; // @[hash.scala 41:22]
  reg [15:0] phv_header_4; // @[hash.scala 41:22]
  reg [15:0] phv_header_5; // @[hash.scala 41:22]
  reg [15:0] phv_header_6; // @[hash.scala 41:22]
  reg [15:0] phv_header_7; // @[hash.scala 41:22]
  reg [15:0] phv_header_8; // @[hash.scala 41:22]
  reg [15:0] phv_header_9; // @[hash.scala 41:22]
  reg [15:0] phv_header_10; // @[hash.scala 41:22]
  reg [15:0] phv_header_11; // @[hash.scala 41:22]
  reg [15:0] phv_header_12; // @[hash.scala 41:22]
  reg [15:0] phv_header_13; // @[hash.scala 41:22]
  reg [15:0] phv_header_14; // @[hash.scala 41:22]
  reg [15:0] phv_header_15; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 41:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 41:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 41:22]
  reg  phv_next_config_id; // @[hash.scala 41:22]
  reg  phv_is_valid_processor; // @[hash.scala 41:22]
  reg [191:0] key; // @[hash.scala 45:22]
  reg [191:0] sum; // @[hash.scala 49:22]
  wire [15:0] sum_temp_0 = sum[191:176]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_1 = sum[175:160]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_2 = sum[159:144]; // @[hash.scala 64:35]
  wire [15:0] out_temp_0 = sum_temp_0 + sum_temp_1; // @[hash.scala 70:51]
  wire [31:0] _io_sum_out_T = {out_temp_0,sum_temp_2}; // @[Cat.scala 30:58]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 43:25]
  assign io_key_out = key; // @[hash.scala 47:20]
  assign io_sum_out = phv_is_valid_processor ? {{160'd0}, _io_sum_out_T} : sum; // @[hash.scala 52:39 hash.scala 75:24 hash.scala 77:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 42:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 42:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 42:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 42:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 42:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 42:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 42:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 42:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 42:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 42:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 42:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 42:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 42:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 42:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 42:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 42:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 42:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 42:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 42:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 42:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 42:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 42:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 42:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 42:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 42:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 42:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 42:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 42:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 42:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 42:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 42:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 42:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 42:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 42:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 42:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 42:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 42:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 42:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 42:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 42:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 42:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 42:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 42:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 42:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 42:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 42:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 42:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 42:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 42:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 42:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 42:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 42:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 42:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 42:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 42:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 42:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 42:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 42:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 42:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 42:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 42:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 42:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 42:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 42:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 42:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 42:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 42:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 42:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 42:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 42:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 42:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 42:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 42:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 42:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 42:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 42:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 42:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 42:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 42:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 42:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 42:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 42:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 42:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 42:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 42:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 42:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 42:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 42:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 42:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 42:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 42:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 42:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 42:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 42:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 42:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 42:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 42:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 42:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 42:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 42:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 42:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 42:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 42:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 42:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 42:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 42:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 42:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 42:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 42:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 42:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 42:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 42:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 42:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 42:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 42:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 42:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 42:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 42:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 42:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 42:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 42:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 42:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 42:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 42:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 42:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 42:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 42:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 42:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 42:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 42:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 42:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 42:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 42:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 42:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 42:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 42:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 42:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 42:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 42:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 42:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 42:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 42:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 42:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 42:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 42:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 42:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 42:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 42:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 42:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 42:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 42:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 42:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 42:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 42:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 42:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 42:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 42:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 42:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 42:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 42:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 42:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 42:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 42:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 42:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 42:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 42:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 42:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 42:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 42:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 42:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 42:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 42:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 42:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 42:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 42:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 42:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 42:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 42:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 42:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 42:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 42:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 42:13]
    key <= io_key_in; // @[hash.scala 46:13]
    sum <= io_sum_in; // @[hash.scala 50:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {6{`RANDOM}};
  sum = _RAND_183[191:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashSumLevel_3(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [191:0] io_sum_in,
  output [191:0] io_sum_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [191:0] _RAND_183;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 41:22]
  reg [7:0] phv_data_1; // @[hash.scala 41:22]
  reg [7:0] phv_data_2; // @[hash.scala 41:22]
  reg [7:0] phv_data_3; // @[hash.scala 41:22]
  reg [7:0] phv_data_4; // @[hash.scala 41:22]
  reg [7:0] phv_data_5; // @[hash.scala 41:22]
  reg [7:0] phv_data_6; // @[hash.scala 41:22]
  reg [7:0] phv_data_7; // @[hash.scala 41:22]
  reg [7:0] phv_data_8; // @[hash.scala 41:22]
  reg [7:0] phv_data_9; // @[hash.scala 41:22]
  reg [7:0] phv_data_10; // @[hash.scala 41:22]
  reg [7:0] phv_data_11; // @[hash.scala 41:22]
  reg [7:0] phv_data_12; // @[hash.scala 41:22]
  reg [7:0] phv_data_13; // @[hash.scala 41:22]
  reg [7:0] phv_data_14; // @[hash.scala 41:22]
  reg [7:0] phv_data_15; // @[hash.scala 41:22]
  reg [7:0] phv_data_16; // @[hash.scala 41:22]
  reg [7:0] phv_data_17; // @[hash.scala 41:22]
  reg [7:0] phv_data_18; // @[hash.scala 41:22]
  reg [7:0] phv_data_19; // @[hash.scala 41:22]
  reg [7:0] phv_data_20; // @[hash.scala 41:22]
  reg [7:0] phv_data_21; // @[hash.scala 41:22]
  reg [7:0] phv_data_22; // @[hash.scala 41:22]
  reg [7:0] phv_data_23; // @[hash.scala 41:22]
  reg [7:0] phv_data_24; // @[hash.scala 41:22]
  reg [7:0] phv_data_25; // @[hash.scala 41:22]
  reg [7:0] phv_data_26; // @[hash.scala 41:22]
  reg [7:0] phv_data_27; // @[hash.scala 41:22]
  reg [7:0] phv_data_28; // @[hash.scala 41:22]
  reg [7:0] phv_data_29; // @[hash.scala 41:22]
  reg [7:0] phv_data_30; // @[hash.scala 41:22]
  reg [7:0] phv_data_31; // @[hash.scala 41:22]
  reg [7:0] phv_data_32; // @[hash.scala 41:22]
  reg [7:0] phv_data_33; // @[hash.scala 41:22]
  reg [7:0] phv_data_34; // @[hash.scala 41:22]
  reg [7:0] phv_data_35; // @[hash.scala 41:22]
  reg [7:0] phv_data_36; // @[hash.scala 41:22]
  reg [7:0] phv_data_37; // @[hash.scala 41:22]
  reg [7:0] phv_data_38; // @[hash.scala 41:22]
  reg [7:0] phv_data_39; // @[hash.scala 41:22]
  reg [7:0] phv_data_40; // @[hash.scala 41:22]
  reg [7:0] phv_data_41; // @[hash.scala 41:22]
  reg [7:0] phv_data_42; // @[hash.scala 41:22]
  reg [7:0] phv_data_43; // @[hash.scala 41:22]
  reg [7:0] phv_data_44; // @[hash.scala 41:22]
  reg [7:0] phv_data_45; // @[hash.scala 41:22]
  reg [7:0] phv_data_46; // @[hash.scala 41:22]
  reg [7:0] phv_data_47; // @[hash.scala 41:22]
  reg [7:0] phv_data_48; // @[hash.scala 41:22]
  reg [7:0] phv_data_49; // @[hash.scala 41:22]
  reg [7:0] phv_data_50; // @[hash.scala 41:22]
  reg [7:0] phv_data_51; // @[hash.scala 41:22]
  reg [7:0] phv_data_52; // @[hash.scala 41:22]
  reg [7:0] phv_data_53; // @[hash.scala 41:22]
  reg [7:0] phv_data_54; // @[hash.scala 41:22]
  reg [7:0] phv_data_55; // @[hash.scala 41:22]
  reg [7:0] phv_data_56; // @[hash.scala 41:22]
  reg [7:0] phv_data_57; // @[hash.scala 41:22]
  reg [7:0] phv_data_58; // @[hash.scala 41:22]
  reg [7:0] phv_data_59; // @[hash.scala 41:22]
  reg [7:0] phv_data_60; // @[hash.scala 41:22]
  reg [7:0] phv_data_61; // @[hash.scala 41:22]
  reg [7:0] phv_data_62; // @[hash.scala 41:22]
  reg [7:0] phv_data_63; // @[hash.scala 41:22]
  reg [7:0] phv_data_64; // @[hash.scala 41:22]
  reg [7:0] phv_data_65; // @[hash.scala 41:22]
  reg [7:0] phv_data_66; // @[hash.scala 41:22]
  reg [7:0] phv_data_67; // @[hash.scala 41:22]
  reg [7:0] phv_data_68; // @[hash.scala 41:22]
  reg [7:0] phv_data_69; // @[hash.scala 41:22]
  reg [7:0] phv_data_70; // @[hash.scala 41:22]
  reg [7:0] phv_data_71; // @[hash.scala 41:22]
  reg [7:0] phv_data_72; // @[hash.scala 41:22]
  reg [7:0] phv_data_73; // @[hash.scala 41:22]
  reg [7:0] phv_data_74; // @[hash.scala 41:22]
  reg [7:0] phv_data_75; // @[hash.scala 41:22]
  reg [7:0] phv_data_76; // @[hash.scala 41:22]
  reg [7:0] phv_data_77; // @[hash.scala 41:22]
  reg [7:0] phv_data_78; // @[hash.scala 41:22]
  reg [7:0] phv_data_79; // @[hash.scala 41:22]
  reg [7:0] phv_data_80; // @[hash.scala 41:22]
  reg [7:0] phv_data_81; // @[hash.scala 41:22]
  reg [7:0] phv_data_82; // @[hash.scala 41:22]
  reg [7:0] phv_data_83; // @[hash.scala 41:22]
  reg [7:0] phv_data_84; // @[hash.scala 41:22]
  reg [7:0] phv_data_85; // @[hash.scala 41:22]
  reg [7:0] phv_data_86; // @[hash.scala 41:22]
  reg [7:0] phv_data_87; // @[hash.scala 41:22]
  reg [7:0] phv_data_88; // @[hash.scala 41:22]
  reg [7:0] phv_data_89; // @[hash.scala 41:22]
  reg [7:0] phv_data_90; // @[hash.scala 41:22]
  reg [7:0] phv_data_91; // @[hash.scala 41:22]
  reg [7:0] phv_data_92; // @[hash.scala 41:22]
  reg [7:0] phv_data_93; // @[hash.scala 41:22]
  reg [7:0] phv_data_94; // @[hash.scala 41:22]
  reg [7:0] phv_data_95; // @[hash.scala 41:22]
  reg [7:0] phv_data_96; // @[hash.scala 41:22]
  reg [7:0] phv_data_97; // @[hash.scala 41:22]
  reg [7:0] phv_data_98; // @[hash.scala 41:22]
  reg [7:0] phv_data_99; // @[hash.scala 41:22]
  reg [7:0] phv_data_100; // @[hash.scala 41:22]
  reg [7:0] phv_data_101; // @[hash.scala 41:22]
  reg [7:0] phv_data_102; // @[hash.scala 41:22]
  reg [7:0] phv_data_103; // @[hash.scala 41:22]
  reg [7:0] phv_data_104; // @[hash.scala 41:22]
  reg [7:0] phv_data_105; // @[hash.scala 41:22]
  reg [7:0] phv_data_106; // @[hash.scala 41:22]
  reg [7:0] phv_data_107; // @[hash.scala 41:22]
  reg [7:0] phv_data_108; // @[hash.scala 41:22]
  reg [7:0] phv_data_109; // @[hash.scala 41:22]
  reg [7:0] phv_data_110; // @[hash.scala 41:22]
  reg [7:0] phv_data_111; // @[hash.scala 41:22]
  reg [7:0] phv_data_112; // @[hash.scala 41:22]
  reg [7:0] phv_data_113; // @[hash.scala 41:22]
  reg [7:0] phv_data_114; // @[hash.scala 41:22]
  reg [7:0] phv_data_115; // @[hash.scala 41:22]
  reg [7:0] phv_data_116; // @[hash.scala 41:22]
  reg [7:0] phv_data_117; // @[hash.scala 41:22]
  reg [7:0] phv_data_118; // @[hash.scala 41:22]
  reg [7:0] phv_data_119; // @[hash.scala 41:22]
  reg [7:0] phv_data_120; // @[hash.scala 41:22]
  reg [7:0] phv_data_121; // @[hash.scala 41:22]
  reg [7:0] phv_data_122; // @[hash.scala 41:22]
  reg [7:0] phv_data_123; // @[hash.scala 41:22]
  reg [7:0] phv_data_124; // @[hash.scala 41:22]
  reg [7:0] phv_data_125; // @[hash.scala 41:22]
  reg [7:0] phv_data_126; // @[hash.scala 41:22]
  reg [7:0] phv_data_127; // @[hash.scala 41:22]
  reg [7:0] phv_data_128; // @[hash.scala 41:22]
  reg [7:0] phv_data_129; // @[hash.scala 41:22]
  reg [7:0] phv_data_130; // @[hash.scala 41:22]
  reg [7:0] phv_data_131; // @[hash.scala 41:22]
  reg [7:0] phv_data_132; // @[hash.scala 41:22]
  reg [7:0] phv_data_133; // @[hash.scala 41:22]
  reg [7:0] phv_data_134; // @[hash.scala 41:22]
  reg [7:0] phv_data_135; // @[hash.scala 41:22]
  reg [7:0] phv_data_136; // @[hash.scala 41:22]
  reg [7:0] phv_data_137; // @[hash.scala 41:22]
  reg [7:0] phv_data_138; // @[hash.scala 41:22]
  reg [7:0] phv_data_139; // @[hash.scala 41:22]
  reg [7:0] phv_data_140; // @[hash.scala 41:22]
  reg [7:0] phv_data_141; // @[hash.scala 41:22]
  reg [7:0] phv_data_142; // @[hash.scala 41:22]
  reg [7:0] phv_data_143; // @[hash.scala 41:22]
  reg [7:0] phv_data_144; // @[hash.scala 41:22]
  reg [7:0] phv_data_145; // @[hash.scala 41:22]
  reg [7:0] phv_data_146; // @[hash.scala 41:22]
  reg [7:0] phv_data_147; // @[hash.scala 41:22]
  reg [7:0] phv_data_148; // @[hash.scala 41:22]
  reg [7:0] phv_data_149; // @[hash.scala 41:22]
  reg [7:0] phv_data_150; // @[hash.scala 41:22]
  reg [7:0] phv_data_151; // @[hash.scala 41:22]
  reg [7:0] phv_data_152; // @[hash.scala 41:22]
  reg [7:0] phv_data_153; // @[hash.scala 41:22]
  reg [7:0] phv_data_154; // @[hash.scala 41:22]
  reg [7:0] phv_data_155; // @[hash.scala 41:22]
  reg [7:0] phv_data_156; // @[hash.scala 41:22]
  reg [7:0] phv_data_157; // @[hash.scala 41:22]
  reg [7:0] phv_data_158; // @[hash.scala 41:22]
  reg [7:0] phv_data_159; // @[hash.scala 41:22]
  reg [15:0] phv_header_0; // @[hash.scala 41:22]
  reg [15:0] phv_header_1; // @[hash.scala 41:22]
  reg [15:0] phv_header_2; // @[hash.scala 41:22]
  reg [15:0] phv_header_3; // @[hash.scala 41:22]
  reg [15:0] phv_header_4; // @[hash.scala 41:22]
  reg [15:0] phv_header_5; // @[hash.scala 41:22]
  reg [15:0] phv_header_6; // @[hash.scala 41:22]
  reg [15:0] phv_header_7; // @[hash.scala 41:22]
  reg [15:0] phv_header_8; // @[hash.scala 41:22]
  reg [15:0] phv_header_9; // @[hash.scala 41:22]
  reg [15:0] phv_header_10; // @[hash.scala 41:22]
  reg [15:0] phv_header_11; // @[hash.scala 41:22]
  reg [15:0] phv_header_12; // @[hash.scala 41:22]
  reg [15:0] phv_header_13; // @[hash.scala 41:22]
  reg [15:0] phv_header_14; // @[hash.scala 41:22]
  reg [15:0] phv_header_15; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 41:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 41:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 41:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 41:22]
  reg  phv_next_config_id; // @[hash.scala 41:22]
  reg  phv_is_valid_processor; // @[hash.scala 41:22]
  reg [191:0] key; // @[hash.scala 45:22]
  reg [191:0] sum; // @[hash.scala 49:22]
  wire [15:0] sum_temp_0 = sum[191:176]; // @[hash.scala 64:35]
  wire [15:0] sum_temp_1 = sum[175:160]; // @[hash.scala 64:35]
  wire [15:0] out_temp_0 = sum_temp_0 + sum_temp_1; // @[hash.scala 70:51]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 43:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 43:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 43:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 43:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 43:25]
  assign io_key_out = key; // @[hash.scala 47:20]
  assign io_sum_out = phv_is_valid_processor ? {{176'd0}, out_temp_0} : sum; // @[hash.scala 52:39 hash.scala 75:24 hash.scala 77:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 42:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 42:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 42:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 42:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 42:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 42:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 42:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 42:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 42:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 42:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 42:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 42:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 42:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 42:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 42:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 42:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 42:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 42:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 42:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 42:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 42:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 42:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 42:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 42:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 42:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 42:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 42:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 42:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 42:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 42:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 42:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 42:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 42:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 42:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 42:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 42:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 42:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 42:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 42:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 42:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 42:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 42:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 42:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 42:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 42:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 42:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 42:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 42:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 42:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 42:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 42:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 42:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 42:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 42:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 42:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 42:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 42:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 42:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 42:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 42:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 42:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 42:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 42:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 42:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 42:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 42:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 42:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 42:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 42:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 42:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 42:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 42:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 42:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 42:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 42:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 42:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 42:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 42:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 42:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 42:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 42:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 42:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 42:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 42:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 42:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 42:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 42:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 42:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 42:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 42:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 42:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 42:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 42:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 42:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 42:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 42:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 42:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 42:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 42:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 42:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 42:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 42:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 42:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 42:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 42:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 42:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 42:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 42:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 42:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 42:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 42:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 42:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 42:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 42:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 42:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 42:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 42:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 42:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 42:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 42:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 42:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 42:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 42:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 42:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 42:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 42:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 42:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 42:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 42:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 42:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 42:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 42:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 42:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 42:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 42:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 42:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 42:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 42:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 42:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 42:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 42:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 42:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 42:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 42:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 42:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 42:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 42:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 42:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 42:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 42:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 42:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 42:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 42:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 42:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 42:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 42:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 42:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 42:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 42:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 42:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 42:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 42:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 42:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 42:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 42:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 42:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 42:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 42:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 42:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 42:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 42:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 42:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 42:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 42:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 42:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 42:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 42:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 42:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 42:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 42:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 42:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 42:13]
    key <= io_key_in; // @[hash.scala 46:13]
    sum <= io_sum_in; // @[hash.scala 50:13]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {6{`RANDOM}};
  sum = _RAND_183[191:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashReshapeLevel(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [3:0]   io_hash_depth_0,
  input  [3:0]   io_hash_depth_1,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [15:0]  io_sum_in,
  output [15:0]  io_sum_out,
  output [15:0]  io_val_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 94:22]
  reg [7:0] phv_data_1; // @[hash.scala 94:22]
  reg [7:0] phv_data_2; // @[hash.scala 94:22]
  reg [7:0] phv_data_3; // @[hash.scala 94:22]
  reg [7:0] phv_data_4; // @[hash.scala 94:22]
  reg [7:0] phv_data_5; // @[hash.scala 94:22]
  reg [7:0] phv_data_6; // @[hash.scala 94:22]
  reg [7:0] phv_data_7; // @[hash.scala 94:22]
  reg [7:0] phv_data_8; // @[hash.scala 94:22]
  reg [7:0] phv_data_9; // @[hash.scala 94:22]
  reg [7:0] phv_data_10; // @[hash.scala 94:22]
  reg [7:0] phv_data_11; // @[hash.scala 94:22]
  reg [7:0] phv_data_12; // @[hash.scala 94:22]
  reg [7:0] phv_data_13; // @[hash.scala 94:22]
  reg [7:0] phv_data_14; // @[hash.scala 94:22]
  reg [7:0] phv_data_15; // @[hash.scala 94:22]
  reg [7:0] phv_data_16; // @[hash.scala 94:22]
  reg [7:0] phv_data_17; // @[hash.scala 94:22]
  reg [7:0] phv_data_18; // @[hash.scala 94:22]
  reg [7:0] phv_data_19; // @[hash.scala 94:22]
  reg [7:0] phv_data_20; // @[hash.scala 94:22]
  reg [7:0] phv_data_21; // @[hash.scala 94:22]
  reg [7:0] phv_data_22; // @[hash.scala 94:22]
  reg [7:0] phv_data_23; // @[hash.scala 94:22]
  reg [7:0] phv_data_24; // @[hash.scala 94:22]
  reg [7:0] phv_data_25; // @[hash.scala 94:22]
  reg [7:0] phv_data_26; // @[hash.scala 94:22]
  reg [7:0] phv_data_27; // @[hash.scala 94:22]
  reg [7:0] phv_data_28; // @[hash.scala 94:22]
  reg [7:0] phv_data_29; // @[hash.scala 94:22]
  reg [7:0] phv_data_30; // @[hash.scala 94:22]
  reg [7:0] phv_data_31; // @[hash.scala 94:22]
  reg [7:0] phv_data_32; // @[hash.scala 94:22]
  reg [7:0] phv_data_33; // @[hash.scala 94:22]
  reg [7:0] phv_data_34; // @[hash.scala 94:22]
  reg [7:0] phv_data_35; // @[hash.scala 94:22]
  reg [7:0] phv_data_36; // @[hash.scala 94:22]
  reg [7:0] phv_data_37; // @[hash.scala 94:22]
  reg [7:0] phv_data_38; // @[hash.scala 94:22]
  reg [7:0] phv_data_39; // @[hash.scala 94:22]
  reg [7:0] phv_data_40; // @[hash.scala 94:22]
  reg [7:0] phv_data_41; // @[hash.scala 94:22]
  reg [7:0] phv_data_42; // @[hash.scala 94:22]
  reg [7:0] phv_data_43; // @[hash.scala 94:22]
  reg [7:0] phv_data_44; // @[hash.scala 94:22]
  reg [7:0] phv_data_45; // @[hash.scala 94:22]
  reg [7:0] phv_data_46; // @[hash.scala 94:22]
  reg [7:0] phv_data_47; // @[hash.scala 94:22]
  reg [7:0] phv_data_48; // @[hash.scala 94:22]
  reg [7:0] phv_data_49; // @[hash.scala 94:22]
  reg [7:0] phv_data_50; // @[hash.scala 94:22]
  reg [7:0] phv_data_51; // @[hash.scala 94:22]
  reg [7:0] phv_data_52; // @[hash.scala 94:22]
  reg [7:0] phv_data_53; // @[hash.scala 94:22]
  reg [7:0] phv_data_54; // @[hash.scala 94:22]
  reg [7:0] phv_data_55; // @[hash.scala 94:22]
  reg [7:0] phv_data_56; // @[hash.scala 94:22]
  reg [7:0] phv_data_57; // @[hash.scala 94:22]
  reg [7:0] phv_data_58; // @[hash.scala 94:22]
  reg [7:0] phv_data_59; // @[hash.scala 94:22]
  reg [7:0] phv_data_60; // @[hash.scala 94:22]
  reg [7:0] phv_data_61; // @[hash.scala 94:22]
  reg [7:0] phv_data_62; // @[hash.scala 94:22]
  reg [7:0] phv_data_63; // @[hash.scala 94:22]
  reg [7:0] phv_data_64; // @[hash.scala 94:22]
  reg [7:0] phv_data_65; // @[hash.scala 94:22]
  reg [7:0] phv_data_66; // @[hash.scala 94:22]
  reg [7:0] phv_data_67; // @[hash.scala 94:22]
  reg [7:0] phv_data_68; // @[hash.scala 94:22]
  reg [7:0] phv_data_69; // @[hash.scala 94:22]
  reg [7:0] phv_data_70; // @[hash.scala 94:22]
  reg [7:0] phv_data_71; // @[hash.scala 94:22]
  reg [7:0] phv_data_72; // @[hash.scala 94:22]
  reg [7:0] phv_data_73; // @[hash.scala 94:22]
  reg [7:0] phv_data_74; // @[hash.scala 94:22]
  reg [7:0] phv_data_75; // @[hash.scala 94:22]
  reg [7:0] phv_data_76; // @[hash.scala 94:22]
  reg [7:0] phv_data_77; // @[hash.scala 94:22]
  reg [7:0] phv_data_78; // @[hash.scala 94:22]
  reg [7:0] phv_data_79; // @[hash.scala 94:22]
  reg [7:0] phv_data_80; // @[hash.scala 94:22]
  reg [7:0] phv_data_81; // @[hash.scala 94:22]
  reg [7:0] phv_data_82; // @[hash.scala 94:22]
  reg [7:0] phv_data_83; // @[hash.scala 94:22]
  reg [7:0] phv_data_84; // @[hash.scala 94:22]
  reg [7:0] phv_data_85; // @[hash.scala 94:22]
  reg [7:0] phv_data_86; // @[hash.scala 94:22]
  reg [7:0] phv_data_87; // @[hash.scala 94:22]
  reg [7:0] phv_data_88; // @[hash.scala 94:22]
  reg [7:0] phv_data_89; // @[hash.scala 94:22]
  reg [7:0] phv_data_90; // @[hash.scala 94:22]
  reg [7:0] phv_data_91; // @[hash.scala 94:22]
  reg [7:0] phv_data_92; // @[hash.scala 94:22]
  reg [7:0] phv_data_93; // @[hash.scala 94:22]
  reg [7:0] phv_data_94; // @[hash.scala 94:22]
  reg [7:0] phv_data_95; // @[hash.scala 94:22]
  reg [7:0] phv_data_96; // @[hash.scala 94:22]
  reg [7:0] phv_data_97; // @[hash.scala 94:22]
  reg [7:0] phv_data_98; // @[hash.scala 94:22]
  reg [7:0] phv_data_99; // @[hash.scala 94:22]
  reg [7:0] phv_data_100; // @[hash.scala 94:22]
  reg [7:0] phv_data_101; // @[hash.scala 94:22]
  reg [7:0] phv_data_102; // @[hash.scala 94:22]
  reg [7:0] phv_data_103; // @[hash.scala 94:22]
  reg [7:0] phv_data_104; // @[hash.scala 94:22]
  reg [7:0] phv_data_105; // @[hash.scala 94:22]
  reg [7:0] phv_data_106; // @[hash.scala 94:22]
  reg [7:0] phv_data_107; // @[hash.scala 94:22]
  reg [7:0] phv_data_108; // @[hash.scala 94:22]
  reg [7:0] phv_data_109; // @[hash.scala 94:22]
  reg [7:0] phv_data_110; // @[hash.scala 94:22]
  reg [7:0] phv_data_111; // @[hash.scala 94:22]
  reg [7:0] phv_data_112; // @[hash.scala 94:22]
  reg [7:0] phv_data_113; // @[hash.scala 94:22]
  reg [7:0] phv_data_114; // @[hash.scala 94:22]
  reg [7:0] phv_data_115; // @[hash.scala 94:22]
  reg [7:0] phv_data_116; // @[hash.scala 94:22]
  reg [7:0] phv_data_117; // @[hash.scala 94:22]
  reg [7:0] phv_data_118; // @[hash.scala 94:22]
  reg [7:0] phv_data_119; // @[hash.scala 94:22]
  reg [7:0] phv_data_120; // @[hash.scala 94:22]
  reg [7:0] phv_data_121; // @[hash.scala 94:22]
  reg [7:0] phv_data_122; // @[hash.scala 94:22]
  reg [7:0] phv_data_123; // @[hash.scala 94:22]
  reg [7:0] phv_data_124; // @[hash.scala 94:22]
  reg [7:0] phv_data_125; // @[hash.scala 94:22]
  reg [7:0] phv_data_126; // @[hash.scala 94:22]
  reg [7:0] phv_data_127; // @[hash.scala 94:22]
  reg [7:0] phv_data_128; // @[hash.scala 94:22]
  reg [7:0] phv_data_129; // @[hash.scala 94:22]
  reg [7:0] phv_data_130; // @[hash.scala 94:22]
  reg [7:0] phv_data_131; // @[hash.scala 94:22]
  reg [7:0] phv_data_132; // @[hash.scala 94:22]
  reg [7:0] phv_data_133; // @[hash.scala 94:22]
  reg [7:0] phv_data_134; // @[hash.scala 94:22]
  reg [7:0] phv_data_135; // @[hash.scala 94:22]
  reg [7:0] phv_data_136; // @[hash.scala 94:22]
  reg [7:0] phv_data_137; // @[hash.scala 94:22]
  reg [7:0] phv_data_138; // @[hash.scala 94:22]
  reg [7:0] phv_data_139; // @[hash.scala 94:22]
  reg [7:0] phv_data_140; // @[hash.scala 94:22]
  reg [7:0] phv_data_141; // @[hash.scala 94:22]
  reg [7:0] phv_data_142; // @[hash.scala 94:22]
  reg [7:0] phv_data_143; // @[hash.scala 94:22]
  reg [7:0] phv_data_144; // @[hash.scala 94:22]
  reg [7:0] phv_data_145; // @[hash.scala 94:22]
  reg [7:0] phv_data_146; // @[hash.scala 94:22]
  reg [7:0] phv_data_147; // @[hash.scala 94:22]
  reg [7:0] phv_data_148; // @[hash.scala 94:22]
  reg [7:0] phv_data_149; // @[hash.scala 94:22]
  reg [7:0] phv_data_150; // @[hash.scala 94:22]
  reg [7:0] phv_data_151; // @[hash.scala 94:22]
  reg [7:0] phv_data_152; // @[hash.scala 94:22]
  reg [7:0] phv_data_153; // @[hash.scala 94:22]
  reg [7:0] phv_data_154; // @[hash.scala 94:22]
  reg [7:0] phv_data_155; // @[hash.scala 94:22]
  reg [7:0] phv_data_156; // @[hash.scala 94:22]
  reg [7:0] phv_data_157; // @[hash.scala 94:22]
  reg [7:0] phv_data_158; // @[hash.scala 94:22]
  reg [7:0] phv_data_159; // @[hash.scala 94:22]
  reg [15:0] phv_header_0; // @[hash.scala 94:22]
  reg [15:0] phv_header_1; // @[hash.scala 94:22]
  reg [15:0] phv_header_2; // @[hash.scala 94:22]
  reg [15:0] phv_header_3; // @[hash.scala 94:22]
  reg [15:0] phv_header_4; // @[hash.scala 94:22]
  reg [15:0] phv_header_5; // @[hash.scala 94:22]
  reg [15:0] phv_header_6; // @[hash.scala 94:22]
  reg [15:0] phv_header_7; // @[hash.scala 94:22]
  reg [15:0] phv_header_8; // @[hash.scala 94:22]
  reg [15:0] phv_header_9; // @[hash.scala 94:22]
  reg [15:0] phv_header_10; // @[hash.scala 94:22]
  reg [15:0] phv_header_11; // @[hash.scala 94:22]
  reg [15:0] phv_header_12; // @[hash.scala 94:22]
  reg [15:0] phv_header_13; // @[hash.scala 94:22]
  reg [15:0] phv_header_14; // @[hash.scala 94:22]
  reg [15:0] phv_header_15; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 94:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 94:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 94:22]
  reg  phv_next_config_id; // @[hash.scala 94:22]
  reg  phv_is_valid_processor; // @[hash.scala 94:22]
  reg [191:0] key; // @[hash.scala 98:22]
  reg [15:0] sum; // @[hash.scala 102:22]
  reg [3:0] hash_depth; // @[hash.scala 106:29]
  wire [16:0] _io_val_out_T_1 = {{1'd0}, sum}; // @[hash.scala 116:44]
  wire [15:0] _GEN_2 = hash_depth[0] ? _io_val_out_T_1[15:0] : 16'h0; // @[hash.scala 115:42 hash.scala 116:32 hash.scala 118:32]
  wire [15:0] _GEN_3 = hash_depth == 4'h0 ? sum : _GEN_2; // @[hash.scala 112:71 hash.scala 113:28]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 96:25]
  assign io_key_out = key; // @[hash.scala 100:20]
  assign io_sum_out = sum; // @[hash.scala 104:20]
  assign io_val_out = phv_is_valid_processor ? _GEN_3 : 16'h0; // @[hash.scala 111:39 hash.scala 122:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 95:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 95:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 95:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 95:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 95:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 95:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 95:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 95:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 95:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 95:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 95:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 95:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 95:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 95:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 95:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 95:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 95:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 95:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 95:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 95:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 95:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 95:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 95:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 95:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 95:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 95:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 95:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 95:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 95:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 95:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 95:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 95:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 95:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 95:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 95:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 95:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 95:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 95:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 95:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 95:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 95:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 95:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 95:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 95:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 95:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 95:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 95:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 95:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 95:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 95:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 95:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 95:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 95:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 95:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 95:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 95:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 95:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 95:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 95:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 95:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 95:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 95:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 95:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 95:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 95:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 95:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 95:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 95:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 95:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 95:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 95:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 95:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 95:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 95:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 95:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 95:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 95:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 95:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 95:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 95:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 95:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 95:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 95:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 95:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 95:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 95:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 95:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 95:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 95:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 95:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 95:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 95:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 95:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 95:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 95:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 95:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 95:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 95:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 95:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 95:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 95:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 95:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 95:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 95:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 95:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 95:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 95:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 95:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 95:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 95:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 95:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 95:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 95:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 95:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 95:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 95:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 95:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 95:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 95:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 95:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 95:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 95:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 95:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 95:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 95:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 95:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 95:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 95:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 95:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 95:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 95:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 95:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 95:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 95:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 95:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 95:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 95:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 95:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 95:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 95:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 95:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 95:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 95:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 95:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 95:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 95:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 95:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 95:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 95:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 95:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 95:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 95:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 95:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 95:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 95:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 95:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 95:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 95:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 95:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 95:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 95:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 95:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 95:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 95:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 95:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 95:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 95:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 95:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 95:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 95:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 95:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 95:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 95:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 95:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 95:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 95:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 95:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 95:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 95:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 95:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 95:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 95:13]
    key <= io_key_in; // @[hash.scala 99:13]
    sum <= io_sum_in; // @[hash.scala 103:13]
    if (io_pipe_phv_in_next_config_id) begin // @[hash.scala 107:20]
      hash_depth <= io_hash_depth_1; // @[hash.scala 107:20]
    end else begin
      hash_depth <= io_hash_depth_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {1{`RANDOM}};
  sum = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  hash_depth = _RAND_184[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashReshapeLevel_1(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [3:0]   io_hash_depth_0,
  input  [3:0]   io_hash_depth_1,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [15:0]  io_sum_in,
  output [15:0]  io_sum_out,
  input  [15:0]  io_val_in,
  output [15:0]  io_val_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 94:22]
  reg [7:0] phv_data_1; // @[hash.scala 94:22]
  reg [7:0] phv_data_2; // @[hash.scala 94:22]
  reg [7:0] phv_data_3; // @[hash.scala 94:22]
  reg [7:0] phv_data_4; // @[hash.scala 94:22]
  reg [7:0] phv_data_5; // @[hash.scala 94:22]
  reg [7:0] phv_data_6; // @[hash.scala 94:22]
  reg [7:0] phv_data_7; // @[hash.scala 94:22]
  reg [7:0] phv_data_8; // @[hash.scala 94:22]
  reg [7:0] phv_data_9; // @[hash.scala 94:22]
  reg [7:0] phv_data_10; // @[hash.scala 94:22]
  reg [7:0] phv_data_11; // @[hash.scala 94:22]
  reg [7:0] phv_data_12; // @[hash.scala 94:22]
  reg [7:0] phv_data_13; // @[hash.scala 94:22]
  reg [7:0] phv_data_14; // @[hash.scala 94:22]
  reg [7:0] phv_data_15; // @[hash.scala 94:22]
  reg [7:0] phv_data_16; // @[hash.scala 94:22]
  reg [7:0] phv_data_17; // @[hash.scala 94:22]
  reg [7:0] phv_data_18; // @[hash.scala 94:22]
  reg [7:0] phv_data_19; // @[hash.scala 94:22]
  reg [7:0] phv_data_20; // @[hash.scala 94:22]
  reg [7:0] phv_data_21; // @[hash.scala 94:22]
  reg [7:0] phv_data_22; // @[hash.scala 94:22]
  reg [7:0] phv_data_23; // @[hash.scala 94:22]
  reg [7:0] phv_data_24; // @[hash.scala 94:22]
  reg [7:0] phv_data_25; // @[hash.scala 94:22]
  reg [7:0] phv_data_26; // @[hash.scala 94:22]
  reg [7:0] phv_data_27; // @[hash.scala 94:22]
  reg [7:0] phv_data_28; // @[hash.scala 94:22]
  reg [7:0] phv_data_29; // @[hash.scala 94:22]
  reg [7:0] phv_data_30; // @[hash.scala 94:22]
  reg [7:0] phv_data_31; // @[hash.scala 94:22]
  reg [7:0] phv_data_32; // @[hash.scala 94:22]
  reg [7:0] phv_data_33; // @[hash.scala 94:22]
  reg [7:0] phv_data_34; // @[hash.scala 94:22]
  reg [7:0] phv_data_35; // @[hash.scala 94:22]
  reg [7:0] phv_data_36; // @[hash.scala 94:22]
  reg [7:0] phv_data_37; // @[hash.scala 94:22]
  reg [7:0] phv_data_38; // @[hash.scala 94:22]
  reg [7:0] phv_data_39; // @[hash.scala 94:22]
  reg [7:0] phv_data_40; // @[hash.scala 94:22]
  reg [7:0] phv_data_41; // @[hash.scala 94:22]
  reg [7:0] phv_data_42; // @[hash.scala 94:22]
  reg [7:0] phv_data_43; // @[hash.scala 94:22]
  reg [7:0] phv_data_44; // @[hash.scala 94:22]
  reg [7:0] phv_data_45; // @[hash.scala 94:22]
  reg [7:0] phv_data_46; // @[hash.scala 94:22]
  reg [7:0] phv_data_47; // @[hash.scala 94:22]
  reg [7:0] phv_data_48; // @[hash.scala 94:22]
  reg [7:0] phv_data_49; // @[hash.scala 94:22]
  reg [7:0] phv_data_50; // @[hash.scala 94:22]
  reg [7:0] phv_data_51; // @[hash.scala 94:22]
  reg [7:0] phv_data_52; // @[hash.scala 94:22]
  reg [7:0] phv_data_53; // @[hash.scala 94:22]
  reg [7:0] phv_data_54; // @[hash.scala 94:22]
  reg [7:0] phv_data_55; // @[hash.scala 94:22]
  reg [7:0] phv_data_56; // @[hash.scala 94:22]
  reg [7:0] phv_data_57; // @[hash.scala 94:22]
  reg [7:0] phv_data_58; // @[hash.scala 94:22]
  reg [7:0] phv_data_59; // @[hash.scala 94:22]
  reg [7:0] phv_data_60; // @[hash.scala 94:22]
  reg [7:0] phv_data_61; // @[hash.scala 94:22]
  reg [7:0] phv_data_62; // @[hash.scala 94:22]
  reg [7:0] phv_data_63; // @[hash.scala 94:22]
  reg [7:0] phv_data_64; // @[hash.scala 94:22]
  reg [7:0] phv_data_65; // @[hash.scala 94:22]
  reg [7:0] phv_data_66; // @[hash.scala 94:22]
  reg [7:0] phv_data_67; // @[hash.scala 94:22]
  reg [7:0] phv_data_68; // @[hash.scala 94:22]
  reg [7:0] phv_data_69; // @[hash.scala 94:22]
  reg [7:0] phv_data_70; // @[hash.scala 94:22]
  reg [7:0] phv_data_71; // @[hash.scala 94:22]
  reg [7:0] phv_data_72; // @[hash.scala 94:22]
  reg [7:0] phv_data_73; // @[hash.scala 94:22]
  reg [7:0] phv_data_74; // @[hash.scala 94:22]
  reg [7:0] phv_data_75; // @[hash.scala 94:22]
  reg [7:0] phv_data_76; // @[hash.scala 94:22]
  reg [7:0] phv_data_77; // @[hash.scala 94:22]
  reg [7:0] phv_data_78; // @[hash.scala 94:22]
  reg [7:0] phv_data_79; // @[hash.scala 94:22]
  reg [7:0] phv_data_80; // @[hash.scala 94:22]
  reg [7:0] phv_data_81; // @[hash.scala 94:22]
  reg [7:0] phv_data_82; // @[hash.scala 94:22]
  reg [7:0] phv_data_83; // @[hash.scala 94:22]
  reg [7:0] phv_data_84; // @[hash.scala 94:22]
  reg [7:0] phv_data_85; // @[hash.scala 94:22]
  reg [7:0] phv_data_86; // @[hash.scala 94:22]
  reg [7:0] phv_data_87; // @[hash.scala 94:22]
  reg [7:0] phv_data_88; // @[hash.scala 94:22]
  reg [7:0] phv_data_89; // @[hash.scala 94:22]
  reg [7:0] phv_data_90; // @[hash.scala 94:22]
  reg [7:0] phv_data_91; // @[hash.scala 94:22]
  reg [7:0] phv_data_92; // @[hash.scala 94:22]
  reg [7:0] phv_data_93; // @[hash.scala 94:22]
  reg [7:0] phv_data_94; // @[hash.scala 94:22]
  reg [7:0] phv_data_95; // @[hash.scala 94:22]
  reg [7:0] phv_data_96; // @[hash.scala 94:22]
  reg [7:0] phv_data_97; // @[hash.scala 94:22]
  reg [7:0] phv_data_98; // @[hash.scala 94:22]
  reg [7:0] phv_data_99; // @[hash.scala 94:22]
  reg [7:0] phv_data_100; // @[hash.scala 94:22]
  reg [7:0] phv_data_101; // @[hash.scala 94:22]
  reg [7:0] phv_data_102; // @[hash.scala 94:22]
  reg [7:0] phv_data_103; // @[hash.scala 94:22]
  reg [7:0] phv_data_104; // @[hash.scala 94:22]
  reg [7:0] phv_data_105; // @[hash.scala 94:22]
  reg [7:0] phv_data_106; // @[hash.scala 94:22]
  reg [7:0] phv_data_107; // @[hash.scala 94:22]
  reg [7:0] phv_data_108; // @[hash.scala 94:22]
  reg [7:0] phv_data_109; // @[hash.scala 94:22]
  reg [7:0] phv_data_110; // @[hash.scala 94:22]
  reg [7:0] phv_data_111; // @[hash.scala 94:22]
  reg [7:0] phv_data_112; // @[hash.scala 94:22]
  reg [7:0] phv_data_113; // @[hash.scala 94:22]
  reg [7:0] phv_data_114; // @[hash.scala 94:22]
  reg [7:0] phv_data_115; // @[hash.scala 94:22]
  reg [7:0] phv_data_116; // @[hash.scala 94:22]
  reg [7:0] phv_data_117; // @[hash.scala 94:22]
  reg [7:0] phv_data_118; // @[hash.scala 94:22]
  reg [7:0] phv_data_119; // @[hash.scala 94:22]
  reg [7:0] phv_data_120; // @[hash.scala 94:22]
  reg [7:0] phv_data_121; // @[hash.scala 94:22]
  reg [7:0] phv_data_122; // @[hash.scala 94:22]
  reg [7:0] phv_data_123; // @[hash.scala 94:22]
  reg [7:0] phv_data_124; // @[hash.scala 94:22]
  reg [7:0] phv_data_125; // @[hash.scala 94:22]
  reg [7:0] phv_data_126; // @[hash.scala 94:22]
  reg [7:0] phv_data_127; // @[hash.scala 94:22]
  reg [7:0] phv_data_128; // @[hash.scala 94:22]
  reg [7:0] phv_data_129; // @[hash.scala 94:22]
  reg [7:0] phv_data_130; // @[hash.scala 94:22]
  reg [7:0] phv_data_131; // @[hash.scala 94:22]
  reg [7:0] phv_data_132; // @[hash.scala 94:22]
  reg [7:0] phv_data_133; // @[hash.scala 94:22]
  reg [7:0] phv_data_134; // @[hash.scala 94:22]
  reg [7:0] phv_data_135; // @[hash.scala 94:22]
  reg [7:0] phv_data_136; // @[hash.scala 94:22]
  reg [7:0] phv_data_137; // @[hash.scala 94:22]
  reg [7:0] phv_data_138; // @[hash.scala 94:22]
  reg [7:0] phv_data_139; // @[hash.scala 94:22]
  reg [7:0] phv_data_140; // @[hash.scala 94:22]
  reg [7:0] phv_data_141; // @[hash.scala 94:22]
  reg [7:0] phv_data_142; // @[hash.scala 94:22]
  reg [7:0] phv_data_143; // @[hash.scala 94:22]
  reg [7:0] phv_data_144; // @[hash.scala 94:22]
  reg [7:0] phv_data_145; // @[hash.scala 94:22]
  reg [7:0] phv_data_146; // @[hash.scala 94:22]
  reg [7:0] phv_data_147; // @[hash.scala 94:22]
  reg [7:0] phv_data_148; // @[hash.scala 94:22]
  reg [7:0] phv_data_149; // @[hash.scala 94:22]
  reg [7:0] phv_data_150; // @[hash.scala 94:22]
  reg [7:0] phv_data_151; // @[hash.scala 94:22]
  reg [7:0] phv_data_152; // @[hash.scala 94:22]
  reg [7:0] phv_data_153; // @[hash.scala 94:22]
  reg [7:0] phv_data_154; // @[hash.scala 94:22]
  reg [7:0] phv_data_155; // @[hash.scala 94:22]
  reg [7:0] phv_data_156; // @[hash.scala 94:22]
  reg [7:0] phv_data_157; // @[hash.scala 94:22]
  reg [7:0] phv_data_158; // @[hash.scala 94:22]
  reg [7:0] phv_data_159; // @[hash.scala 94:22]
  reg [15:0] phv_header_0; // @[hash.scala 94:22]
  reg [15:0] phv_header_1; // @[hash.scala 94:22]
  reg [15:0] phv_header_2; // @[hash.scala 94:22]
  reg [15:0] phv_header_3; // @[hash.scala 94:22]
  reg [15:0] phv_header_4; // @[hash.scala 94:22]
  reg [15:0] phv_header_5; // @[hash.scala 94:22]
  reg [15:0] phv_header_6; // @[hash.scala 94:22]
  reg [15:0] phv_header_7; // @[hash.scala 94:22]
  reg [15:0] phv_header_8; // @[hash.scala 94:22]
  reg [15:0] phv_header_9; // @[hash.scala 94:22]
  reg [15:0] phv_header_10; // @[hash.scala 94:22]
  reg [15:0] phv_header_11; // @[hash.scala 94:22]
  reg [15:0] phv_header_12; // @[hash.scala 94:22]
  reg [15:0] phv_header_13; // @[hash.scala 94:22]
  reg [15:0] phv_header_14; // @[hash.scala 94:22]
  reg [15:0] phv_header_15; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 94:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 94:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 94:22]
  reg  phv_next_config_id; // @[hash.scala 94:22]
  reg  phv_is_valid_processor; // @[hash.scala 94:22]
  reg [191:0] key; // @[hash.scala 98:22]
  reg [15:0] sum; // @[hash.scala 102:22]
  reg [3:0] hash_depth; // @[hash.scala 106:29]
  reg [15:0] hash_val; // @[hash.scala 108:27]
  wire [15:0] _GEN_5 = {{1'd0}, sum[14:0]}; // @[hash.scala 116:44]
  wire [15:0] _io_val_out_T_2 = hash_val + _GEN_5; // @[hash.scala 116:44]
  wire [15:0] _GEN_2 = hash_depth[1] ? _io_val_out_T_2 : hash_val; // @[hash.scala 115:42 hash.scala 116:32 hash.scala 118:32]
  wire [15:0] _GEN_3 = hash_depth == 4'h0 ? sum : _GEN_2; // @[hash.scala 112:71 hash.scala 113:28]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 96:25]
  assign io_key_out = key; // @[hash.scala 100:20]
  assign io_sum_out = sum; // @[hash.scala 104:20]
  assign io_val_out = phv_is_valid_processor ? _GEN_3 : hash_val; // @[hash.scala 111:39 hash.scala 122:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 95:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 95:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 95:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 95:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 95:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 95:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 95:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 95:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 95:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 95:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 95:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 95:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 95:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 95:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 95:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 95:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 95:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 95:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 95:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 95:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 95:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 95:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 95:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 95:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 95:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 95:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 95:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 95:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 95:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 95:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 95:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 95:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 95:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 95:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 95:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 95:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 95:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 95:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 95:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 95:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 95:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 95:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 95:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 95:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 95:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 95:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 95:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 95:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 95:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 95:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 95:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 95:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 95:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 95:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 95:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 95:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 95:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 95:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 95:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 95:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 95:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 95:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 95:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 95:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 95:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 95:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 95:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 95:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 95:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 95:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 95:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 95:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 95:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 95:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 95:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 95:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 95:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 95:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 95:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 95:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 95:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 95:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 95:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 95:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 95:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 95:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 95:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 95:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 95:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 95:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 95:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 95:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 95:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 95:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 95:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 95:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 95:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 95:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 95:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 95:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 95:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 95:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 95:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 95:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 95:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 95:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 95:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 95:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 95:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 95:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 95:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 95:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 95:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 95:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 95:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 95:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 95:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 95:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 95:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 95:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 95:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 95:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 95:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 95:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 95:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 95:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 95:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 95:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 95:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 95:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 95:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 95:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 95:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 95:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 95:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 95:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 95:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 95:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 95:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 95:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 95:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 95:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 95:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 95:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 95:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 95:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 95:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 95:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 95:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 95:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 95:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 95:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 95:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 95:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 95:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 95:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 95:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 95:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 95:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 95:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 95:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 95:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 95:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 95:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 95:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 95:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 95:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 95:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 95:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 95:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 95:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 95:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 95:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 95:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 95:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 95:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 95:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 95:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 95:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 95:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 95:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 95:13]
    key <= io_key_in; // @[hash.scala 99:13]
    sum <= io_sum_in; // @[hash.scala 103:13]
    if (io_pipe_phv_in_next_config_id) begin // @[hash.scala 107:20]
      hash_depth <= io_hash_depth_1; // @[hash.scala 107:20]
    end else begin
      hash_depth <= io_hash_depth_0;
    end
    hash_val <= io_val_in; // @[hash.scala 109:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {1{`RANDOM}};
  sum = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  hash_depth = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  hash_val = _RAND_185[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashReshapeLevel_2(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [3:0]   io_hash_depth_0,
  input  [3:0]   io_hash_depth_1,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [15:0]  io_sum_in,
  output [15:0]  io_sum_out,
  input  [15:0]  io_val_in,
  output [15:0]  io_val_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 94:22]
  reg [7:0] phv_data_1; // @[hash.scala 94:22]
  reg [7:0] phv_data_2; // @[hash.scala 94:22]
  reg [7:0] phv_data_3; // @[hash.scala 94:22]
  reg [7:0] phv_data_4; // @[hash.scala 94:22]
  reg [7:0] phv_data_5; // @[hash.scala 94:22]
  reg [7:0] phv_data_6; // @[hash.scala 94:22]
  reg [7:0] phv_data_7; // @[hash.scala 94:22]
  reg [7:0] phv_data_8; // @[hash.scala 94:22]
  reg [7:0] phv_data_9; // @[hash.scala 94:22]
  reg [7:0] phv_data_10; // @[hash.scala 94:22]
  reg [7:0] phv_data_11; // @[hash.scala 94:22]
  reg [7:0] phv_data_12; // @[hash.scala 94:22]
  reg [7:0] phv_data_13; // @[hash.scala 94:22]
  reg [7:0] phv_data_14; // @[hash.scala 94:22]
  reg [7:0] phv_data_15; // @[hash.scala 94:22]
  reg [7:0] phv_data_16; // @[hash.scala 94:22]
  reg [7:0] phv_data_17; // @[hash.scala 94:22]
  reg [7:0] phv_data_18; // @[hash.scala 94:22]
  reg [7:0] phv_data_19; // @[hash.scala 94:22]
  reg [7:0] phv_data_20; // @[hash.scala 94:22]
  reg [7:0] phv_data_21; // @[hash.scala 94:22]
  reg [7:0] phv_data_22; // @[hash.scala 94:22]
  reg [7:0] phv_data_23; // @[hash.scala 94:22]
  reg [7:0] phv_data_24; // @[hash.scala 94:22]
  reg [7:0] phv_data_25; // @[hash.scala 94:22]
  reg [7:0] phv_data_26; // @[hash.scala 94:22]
  reg [7:0] phv_data_27; // @[hash.scala 94:22]
  reg [7:0] phv_data_28; // @[hash.scala 94:22]
  reg [7:0] phv_data_29; // @[hash.scala 94:22]
  reg [7:0] phv_data_30; // @[hash.scala 94:22]
  reg [7:0] phv_data_31; // @[hash.scala 94:22]
  reg [7:0] phv_data_32; // @[hash.scala 94:22]
  reg [7:0] phv_data_33; // @[hash.scala 94:22]
  reg [7:0] phv_data_34; // @[hash.scala 94:22]
  reg [7:0] phv_data_35; // @[hash.scala 94:22]
  reg [7:0] phv_data_36; // @[hash.scala 94:22]
  reg [7:0] phv_data_37; // @[hash.scala 94:22]
  reg [7:0] phv_data_38; // @[hash.scala 94:22]
  reg [7:0] phv_data_39; // @[hash.scala 94:22]
  reg [7:0] phv_data_40; // @[hash.scala 94:22]
  reg [7:0] phv_data_41; // @[hash.scala 94:22]
  reg [7:0] phv_data_42; // @[hash.scala 94:22]
  reg [7:0] phv_data_43; // @[hash.scala 94:22]
  reg [7:0] phv_data_44; // @[hash.scala 94:22]
  reg [7:0] phv_data_45; // @[hash.scala 94:22]
  reg [7:0] phv_data_46; // @[hash.scala 94:22]
  reg [7:0] phv_data_47; // @[hash.scala 94:22]
  reg [7:0] phv_data_48; // @[hash.scala 94:22]
  reg [7:0] phv_data_49; // @[hash.scala 94:22]
  reg [7:0] phv_data_50; // @[hash.scala 94:22]
  reg [7:0] phv_data_51; // @[hash.scala 94:22]
  reg [7:0] phv_data_52; // @[hash.scala 94:22]
  reg [7:0] phv_data_53; // @[hash.scala 94:22]
  reg [7:0] phv_data_54; // @[hash.scala 94:22]
  reg [7:0] phv_data_55; // @[hash.scala 94:22]
  reg [7:0] phv_data_56; // @[hash.scala 94:22]
  reg [7:0] phv_data_57; // @[hash.scala 94:22]
  reg [7:0] phv_data_58; // @[hash.scala 94:22]
  reg [7:0] phv_data_59; // @[hash.scala 94:22]
  reg [7:0] phv_data_60; // @[hash.scala 94:22]
  reg [7:0] phv_data_61; // @[hash.scala 94:22]
  reg [7:0] phv_data_62; // @[hash.scala 94:22]
  reg [7:0] phv_data_63; // @[hash.scala 94:22]
  reg [7:0] phv_data_64; // @[hash.scala 94:22]
  reg [7:0] phv_data_65; // @[hash.scala 94:22]
  reg [7:0] phv_data_66; // @[hash.scala 94:22]
  reg [7:0] phv_data_67; // @[hash.scala 94:22]
  reg [7:0] phv_data_68; // @[hash.scala 94:22]
  reg [7:0] phv_data_69; // @[hash.scala 94:22]
  reg [7:0] phv_data_70; // @[hash.scala 94:22]
  reg [7:0] phv_data_71; // @[hash.scala 94:22]
  reg [7:0] phv_data_72; // @[hash.scala 94:22]
  reg [7:0] phv_data_73; // @[hash.scala 94:22]
  reg [7:0] phv_data_74; // @[hash.scala 94:22]
  reg [7:0] phv_data_75; // @[hash.scala 94:22]
  reg [7:0] phv_data_76; // @[hash.scala 94:22]
  reg [7:0] phv_data_77; // @[hash.scala 94:22]
  reg [7:0] phv_data_78; // @[hash.scala 94:22]
  reg [7:0] phv_data_79; // @[hash.scala 94:22]
  reg [7:0] phv_data_80; // @[hash.scala 94:22]
  reg [7:0] phv_data_81; // @[hash.scala 94:22]
  reg [7:0] phv_data_82; // @[hash.scala 94:22]
  reg [7:0] phv_data_83; // @[hash.scala 94:22]
  reg [7:0] phv_data_84; // @[hash.scala 94:22]
  reg [7:0] phv_data_85; // @[hash.scala 94:22]
  reg [7:0] phv_data_86; // @[hash.scala 94:22]
  reg [7:0] phv_data_87; // @[hash.scala 94:22]
  reg [7:0] phv_data_88; // @[hash.scala 94:22]
  reg [7:0] phv_data_89; // @[hash.scala 94:22]
  reg [7:0] phv_data_90; // @[hash.scala 94:22]
  reg [7:0] phv_data_91; // @[hash.scala 94:22]
  reg [7:0] phv_data_92; // @[hash.scala 94:22]
  reg [7:0] phv_data_93; // @[hash.scala 94:22]
  reg [7:0] phv_data_94; // @[hash.scala 94:22]
  reg [7:0] phv_data_95; // @[hash.scala 94:22]
  reg [7:0] phv_data_96; // @[hash.scala 94:22]
  reg [7:0] phv_data_97; // @[hash.scala 94:22]
  reg [7:0] phv_data_98; // @[hash.scala 94:22]
  reg [7:0] phv_data_99; // @[hash.scala 94:22]
  reg [7:0] phv_data_100; // @[hash.scala 94:22]
  reg [7:0] phv_data_101; // @[hash.scala 94:22]
  reg [7:0] phv_data_102; // @[hash.scala 94:22]
  reg [7:0] phv_data_103; // @[hash.scala 94:22]
  reg [7:0] phv_data_104; // @[hash.scala 94:22]
  reg [7:0] phv_data_105; // @[hash.scala 94:22]
  reg [7:0] phv_data_106; // @[hash.scala 94:22]
  reg [7:0] phv_data_107; // @[hash.scala 94:22]
  reg [7:0] phv_data_108; // @[hash.scala 94:22]
  reg [7:0] phv_data_109; // @[hash.scala 94:22]
  reg [7:0] phv_data_110; // @[hash.scala 94:22]
  reg [7:0] phv_data_111; // @[hash.scala 94:22]
  reg [7:0] phv_data_112; // @[hash.scala 94:22]
  reg [7:0] phv_data_113; // @[hash.scala 94:22]
  reg [7:0] phv_data_114; // @[hash.scala 94:22]
  reg [7:0] phv_data_115; // @[hash.scala 94:22]
  reg [7:0] phv_data_116; // @[hash.scala 94:22]
  reg [7:0] phv_data_117; // @[hash.scala 94:22]
  reg [7:0] phv_data_118; // @[hash.scala 94:22]
  reg [7:0] phv_data_119; // @[hash.scala 94:22]
  reg [7:0] phv_data_120; // @[hash.scala 94:22]
  reg [7:0] phv_data_121; // @[hash.scala 94:22]
  reg [7:0] phv_data_122; // @[hash.scala 94:22]
  reg [7:0] phv_data_123; // @[hash.scala 94:22]
  reg [7:0] phv_data_124; // @[hash.scala 94:22]
  reg [7:0] phv_data_125; // @[hash.scala 94:22]
  reg [7:0] phv_data_126; // @[hash.scala 94:22]
  reg [7:0] phv_data_127; // @[hash.scala 94:22]
  reg [7:0] phv_data_128; // @[hash.scala 94:22]
  reg [7:0] phv_data_129; // @[hash.scala 94:22]
  reg [7:0] phv_data_130; // @[hash.scala 94:22]
  reg [7:0] phv_data_131; // @[hash.scala 94:22]
  reg [7:0] phv_data_132; // @[hash.scala 94:22]
  reg [7:0] phv_data_133; // @[hash.scala 94:22]
  reg [7:0] phv_data_134; // @[hash.scala 94:22]
  reg [7:0] phv_data_135; // @[hash.scala 94:22]
  reg [7:0] phv_data_136; // @[hash.scala 94:22]
  reg [7:0] phv_data_137; // @[hash.scala 94:22]
  reg [7:0] phv_data_138; // @[hash.scala 94:22]
  reg [7:0] phv_data_139; // @[hash.scala 94:22]
  reg [7:0] phv_data_140; // @[hash.scala 94:22]
  reg [7:0] phv_data_141; // @[hash.scala 94:22]
  reg [7:0] phv_data_142; // @[hash.scala 94:22]
  reg [7:0] phv_data_143; // @[hash.scala 94:22]
  reg [7:0] phv_data_144; // @[hash.scala 94:22]
  reg [7:0] phv_data_145; // @[hash.scala 94:22]
  reg [7:0] phv_data_146; // @[hash.scala 94:22]
  reg [7:0] phv_data_147; // @[hash.scala 94:22]
  reg [7:0] phv_data_148; // @[hash.scala 94:22]
  reg [7:0] phv_data_149; // @[hash.scala 94:22]
  reg [7:0] phv_data_150; // @[hash.scala 94:22]
  reg [7:0] phv_data_151; // @[hash.scala 94:22]
  reg [7:0] phv_data_152; // @[hash.scala 94:22]
  reg [7:0] phv_data_153; // @[hash.scala 94:22]
  reg [7:0] phv_data_154; // @[hash.scala 94:22]
  reg [7:0] phv_data_155; // @[hash.scala 94:22]
  reg [7:0] phv_data_156; // @[hash.scala 94:22]
  reg [7:0] phv_data_157; // @[hash.scala 94:22]
  reg [7:0] phv_data_158; // @[hash.scala 94:22]
  reg [7:0] phv_data_159; // @[hash.scala 94:22]
  reg [15:0] phv_header_0; // @[hash.scala 94:22]
  reg [15:0] phv_header_1; // @[hash.scala 94:22]
  reg [15:0] phv_header_2; // @[hash.scala 94:22]
  reg [15:0] phv_header_3; // @[hash.scala 94:22]
  reg [15:0] phv_header_4; // @[hash.scala 94:22]
  reg [15:0] phv_header_5; // @[hash.scala 94:22]
  reg [15:0] phv_header_6; // @[hash.scala 94:22]
  reg [15:0] phv_header_7; // @[hash.scala 94:22]
  reg [15:0] phv_header_8; // @[hash.scala 94:22]
  reg [15:0] phv_header_9; // @[hash.scala 94:22]
  reg [15:0] phv_header_10; // @[hash.scala 94:22]
  reg [15:0] phv_header_11; // @[hash.scala 94:22]
  reg [15:0] phv_header_12; // @[hash.scala 94:22]
  reg [15:0] phv_header_13; // @[hash.scala 94:22]
  reg [15:0] phv_header_14; // @[hash.scala 94:22]
  reg [15:0] phv_header_15; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 94:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 94:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 94:22]
  reg  phv_next_config_id; // @[hash.scala 94:22]
  reg  phv_is_valid_processor; // @[hash.scala 94:22]
  reg [191:0] key; // @[hash.scala 98:22]
  reg [15:0] sum; // @[hash.scala 102:22]
  reg [3:0] hash_depth; // @[hash.scala 106:29]
  reg [15:0] hash_val; // @[hash.scala 108:27]
  wire [15:0] _GEN_5 = {{2'd0}, sum[13:0]}; // @[hash.scala 116:44]
  wire [15:0] _io_val_out_T_2 = hash_val + _GEN_5; // @[hash.scala 116:44]
  wire [15:0] _GEN_2 = hash_depth[2] ? _io_val_out_T_2 : hash_val; // @[hash.scala 115:42 hash.scala 116:32 hash.scala 118:32]
  wire [15:0] _GEN_3 = hash_depth == 4'h0 ? sum : _GEN_2; // @[hash.scala 112:71 hash.scala 113:28]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 96:25]
  assign io_key_out = key; // @[hash.scala 100:20]
  assign io_sum_out = sum; // @[hash.scala 104:20]
  assign io_val_out = phv_is_valid_processor ? _GEN_3 : hash_val; // @[hash.scala 111:39 hash.scala 122:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 95:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 95:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 95:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 95:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 95:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 95:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 95:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 95:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 95:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 95:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 95:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 95:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 95:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 95:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 95:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 95:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 95:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 95:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 95:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 95:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 95:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 95:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 95:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 95:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 95:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 95:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 95:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 95:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 95:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 95:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 95:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 95:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 95:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 95:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 95:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 95:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 95:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 95:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 95:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 95:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 95:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 95:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 95:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 95:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 95:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 95:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 95:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 95:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 95:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 95:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 95:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 95:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 95:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 95:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 95:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 95:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 95:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 95:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 95:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 95:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 95:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 95:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 95:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 95:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 95:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 95:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 95:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 95:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 95:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 95:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 95:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 95:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 95:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 95:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 95:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 95:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 95:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 95:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 95:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 95:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 95:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 95:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 95:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 95:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 95:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 95:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 95:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 95:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 95:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 95:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 95:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 95:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 95:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 95:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 95:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 95:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 95:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 95:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 95:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 95:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 95:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 95:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 95:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 95:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 95:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 95:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 95:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 95:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 95:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 95:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 95:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 95:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 95:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 95:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 95:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 95:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 95:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 95:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 95:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 95:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 95:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 95:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 95:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 95:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 95:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 95:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 95:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 95:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 95:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 95:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 95:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 95:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 95:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 95:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 95:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 95:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 95:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 95:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 95:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 95:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 95:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 95:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 95:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 95:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 95:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 95:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 95:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 95:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 95:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 95:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 95:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 95:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 95:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 95:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 95:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 95:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 95:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 95:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 95:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 95:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 95:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 95:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 95:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 95:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 95:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 95:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 95:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 95:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 95:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 95:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 95:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 95:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 95:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 95:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 95:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 95:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 95:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 95:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 95:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 95:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 95:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 95:13]
    key <= io_key_in; // @[hash.scala 99:13]
    sum <= io_sum_in; // @[hash.scala 103:13]
    if (io_pipe_phv_in_next_config_id) begin // @[hash.scala 107:20]
      hash_depth <= io_hash_depth_1; // @[hash.scala 107:20]
    end else begin
      hash_depth <= io_hash_depth_0;
    end
    hash_val <= io_val_in; // @[hash.scala 109:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {1{`RANDOM}};
  sum = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  hash_depth = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  hash_val = _RAND_185[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module HashReshapeLevel_3(
  input          clock,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input  [3:0]   io_hash_depth_0,
  input  [3:0]   io_hash_depth_1,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  input  [15:0]  io_sum_in,
  output [15:0]  io_sum_out,
  input  [15:0]  io_val_in,
  output [15:0]  io_val_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] phv_data_0; // @[hash.scala 94:22]
  reg [7:0] phv_data_1; // @[hash.scala 94:22]
  reg [7:0] phv_data_2; // @[hash.scala 94:22]
  reg [7:0] phv_data_3; // @[hash.scala 94:22]
  reg [7:0] phv_data_4; // @[hash.scala 94:22]
  reg [7:0] phv_data_5; // @[hash.scala 94:22]
  reg [7:0] phv_data_6; // @[hash.scala 94:22]
  reg [7:0] phv_data_7; // @[hash.scala 94:22]
  reg [7:0] phv_data_8; // @[hash.scala 94:22]
  reg [7:0] phv_data_9; // @[hash.scala 94:22]
  reg [7:0] phv_data_10; // @[hash.scala 94:22]
  reg [7:0] phv_data_11; // @[hash.scala 94:22]
  reg [7:0] phv_data_12; // @[hash.scala 94:22]
  reg [7:0] phv_data_13; // @[hash.scala 94:22]
  reg [7:0] phv_data_14; // @[hash.scala 94:22]
  reg [7:0] phv_data_15; // @[hash.scala 94:22]
  reg [7:0] phv_data_16; // @[hash.scala 94:22]
  reg [7:0] phv_data_17; // @[hash.scala 94:22]
  reg [7:0] phv_data_18; // @[hash.scala 94:22]
  reg [7:0] phv_data_19; // @[hash.scala 94:22]
  reg [7:0] phv_data_20; // @[hash.scala 94:22]
  reg [7:0] phv_data_21; // @[hash.scala 94:22]
  reg [7:0] phv_data_22; // @[hash.scala 94:22]
  reg [7:0] phv_data_23; // @[hash.scala 94:22]
  reg [7:0] phv_data_24; // @[hash.scala 94:22]
  reg [7:0] phv_data_25; // @[hash.scala 94:22]
  reg [7:0] phv_data_26; // @[hash.scala 94:22]
  reg [7:0] phv_data_27; // @[hash.scala 94:22]
  reg [7:0] phv_data_28; // @[hash.scala 94:22]
  reg [7:0] phv_data_29; // @[hash.scala 94:22]
  reg [7:0] phv_data_30; // @[hash.scala 94:22]
  reg [7:0] phv_data_31; // @[hash.scala 94:22]
  reg [7:0] phv_data_32; // @[hash.scala 94:22]
  reg [7:0] phv_data_33; // @[hash.scala 94:22]
  reg [7:0] phv_data_34; // @[hash.scala 94:22]
  reg [7:0] phv_data_35; // @[hash.scala 94:22]
  reg [7:0] phv_data_36; // @[hash.scala 94:22]
  reg [7:0] phv_data_37; // @[hash.scala 94:22]
  reg [7:0] phv_data_38; // @[hash.scala 94:22]
  reg [7:0] phv_data_39; // @[hash.scala 94:22]
  reg [7:0] phv_data_40; // @[hash.scala 94:22]
  reg [7:0] phv_data_41; // @[hash.scala 94:22]
  reg [7:0] phv_data_42; // @[hash.scala 94:22]
  reg [7:0] phv_data_43; // @[hash.scala 94:22]
  reg [7:0] phv_data_44; // @[hash.scala 94:22]
  reg [7:0] phv_data_45; // @[hash.scala 94:22]
  reg [7:0] phv_data_46; // @[hash.scala 94:22]
  reg [7:0] phv_data_47; // @[hash.scala 94:22]
  reg [7:0] phv_data_48; // @[hash.scala 94:22]
  reg [7:0] phv_data_49; // @[hash.scala 94:22]
  reg [7:0] phv_data_50; // @[hash.scala 94:22]
  reg [7:0] phv_data_51; // @[hash.scala 94:22]
  reg [7:0] phv_data_52; // @[hash.scala 94:22]
  reg [7:0] phv_data_53; // @[hash.scala 94:22]
  reg [7:0] phv_data_54; // @[hash.scala 94:22]
  reg [7:0] phv_data_55; // @[hash.scala 94:22]
  reg [7:0] phv_data_56; // @[hash.scala 94:22]
  reg [7:0] phv_data_57; // @[hash.scala 94:22]
  reg [7:0] phv_data_58; // @[hash.scala 94:22]
  reg [7:0] phv_data_59; // @[hash.scala 94:22]
  reg [7:0] phv_data_60; // @[hash.scala 94:22]
  reg [7:0] phv_data_61; // @[hash.scala 94:22]
  reg [7:0] phv_data_62; // @[hash.scala 94:22]
  reg [7:0] phv_data_63; // @[hash.scala 94:22]
  reg [7:0] phv_data_64; // @[hash.scala 94:22]
  reg [7:0] phv_data_65; // @[hash.scala 94:22]
  reg [7:0] phv_data_66; // @[hash.scala 94:22]
  reg [7:0] phv_data_67; // @[hash.scala 94:22]
  reg [7:0] phv_data_68; // @[hash.scala 94:22]
  reg [7:0] phv_data_69; // @[hash.scala 94:22]
  reg [7:0] phv_data_70; // @[hash.scala 94:22]
  reg [7:0] phv_data_71; // @[hash.scala 94:22]
  reg [7:0] phv_data_72; // @[hash.scala 94:22]
  reg [7:0] phv_data_73; // @[hash.scala 94:22]
  reg [7:0] phv_data_74; // @[hash.scala 94:22]
  reg [7:0] phv_data_75; // @[hash.scala 94:22]
  reg [7:0] phv_data_76; // @[hash.scala 94:22]
  reg [7:0] phv_data_77; // @[hash.scala 94:22]
  reg [7:0] phv_data_78; // @[hash.scala 94:22]
  reg [7:0] phv_data_79; // @[hash.scala 94:22]
  reg [7:0] phv_data_80; // @[hash.scala 94:22]
  reg [7:0] phv_data_81; // @[hash.scala 94:22]
  reg [7:0] phv_data_82; // @[hash.scala 94:22]
  reg [7:0] phv_data_83; // @[hash.scala 94:22]
  reg [7:0] phv_data_84; // @[hash.scala 94:22]
  reg [7:0] phv_data_85; // @[hash.scala 94:22]
  reg [7:0] phv_data_86; // @[hash.scala 94:22]
  reg [7:0] phv_data_87; // @[hash.scala 94:22]
  reg [7:0] phv_data_88; // @[hash.scala 94:22]
  reg [7:0] phv_data_89; // @[hash.scala 94:22]
  reg [7:0] phv_data_90; // @[hash.scala 94:22]
  reg [7:0] phv_data_91; // @[hash.scala 94:22]
  reg [7:0] phv_data_92; // @[hash.scala 94:22]
  reg [7:0] phv_data_93; // @[hash.scala 94:22]
  reg [7:0] phv_data_94; // @[hash.scala 94:22]
  reg [7:0] phv_data_95; // @[hash.scala 94:22]
  reg [7:0] phv_data_96; // @[hash.scala 94:22]
  reg [7:0] phv_data_97; // @[hash.scala 94:22]
  reg [7:0] phv_data_98; // @[hash.scala 94:22]
  reg [7:0] phv_data_99; // @[hash.scala 94:22]
  reg [7:0] phv_data_100; // @[hash.scala 94:22]
  reg [7:0] phv_data_101; // @[hash.scala 94:22]
  reg [7:0] phv_data_102; // @[hash.scala 94:22]
  reg [7:0] phv_data_103; // @[hash.scala 94:22]
  reg [7:0] phv_data_104; // @[hash.scala 94:22]
  reg [7:0] phv_data_105; // @[hash.scala 94:22]
  reg [7:0] phv_data_106; // @[hash.scala 94:22]
  reg [7:0] phv_data_107; // @[hash.scala 94:22]
  reg [7:0] phv_data_108; // @[hash.scala 94:22]
  reg [7:0] phv_data_109; // @[hash.scala 94:22]
  reg [7:0] phv_data_110; // @[hash.scala 94:22]
  reg [7:0] phv_data_111; // @[hash.scala 94:22]
  reg [7:0] phv_data_112; // @[hash.scala 94:22]
  reg [7:0] phv_data_113; // @[hash.scala 94:22]
  reg [7:0] phv_data_114; // @[hash.scala 94:22]
  reg [7:0] phv_data_115; // @[hash.scala 94:22]
  reg [7:0] phv_data_116; // @[hash.scala 94:22]
  reg [7:0] phv_data_117; // @[hash.scala 94:22]
  reg [7:0] phv_data_118; // @[hash.scala 94:22]
  reg [7:0] phv_data_119; // @[hash.scala 94:22]
  reg [7:0] phv_data_120; // @[hash.scala 94:22]
  reg [7:0] phv_data_121; // @[hash.scala 94:22]
  reg [7:0] phv_data_122; // @[hash.scala 94:22]
  reg [7:0] phv_data_123; // @[hash.scala 94:22]
  reg [7:0] phv_data_124; // @[hash.scala 94:22]
  reg [7:0] phv_data_125; // @[hash.scala 94:22]
  reg [7:0] phv_data_126; // @[hash.scala 94:22]
  reg [7:0] phv_data_127; // @[hash.scala 94:22]
  reg [7:0] phv_data_128; // @[hash.scala 94:22]
  reg [7:0] phv_data_129; // @[hash.scala 94:22]
  reg [7:0] phv_data_130; // @[hash.scala 94:22]
  reg [7:0] phv_data_131; // @[hash.scala 94:22]
  reg [7:0] phv_data_132; // @[hash.scala 94:22]
  reg [7:0] phv_data_133; // @[hash.scala 94:22]
  reg [7:0] phv_data_134; // @[hash.scala 94:22]
  reg [7:0] phv_data_135; // @[hash.scala 94:22]
  reg [7:0] phv_data_136; // @[hash.scala 94:22]
  reg [7:0] phv_data_137; // @[hash.scala 94:22]
  reg [7:0] phv_data_138; // @[hash.scala 94:22]
  reg [7:0] phv_data_139; // @[hash.scala 94:22]
  reg [7:0] phv_data_140; // @[hash.scala 94:22]
  reg [7:0] phv_data_141; // @[hash.scala 94:22]
  reg [7:0] phv_data_142; // @[hash.scala 94:22]
  reg [7:0] phv_data_143; // @[hash.scala 94:22]
  reg [7:0] phv_data_144; // @[hash.scala 94:22]
  reg [7:0] phv_data_145; // @[hash.scala 94:22]
  reg [7:0] phv_data_146; // @[hash.scala 94:22]
  reg [7:0] phv_data_147; // @[hash.scala 94:22]
  reg [7:0] phv_data_148; // @[hash.scala 94:22]
  reg [7:0] phv_data_149; // @[hash.scala 94:22]
  reg [7:0] phv_data_150; // @[hash.scala 94:22]
  reg [7:0] phv_data_151; // @[hash.scala 94:22]
  reg [7:0] phv_data_152; // @[hash.scala 94:22]
  reg [7:0] phv_data_153; // @[hash.scala 94:22]
  reg [7:0] phv_data_154; // @[hash.scala 94:22]
  reg [7:0] phv_data_155; // @[hash.scala 94:22]
  reg [7:0] phv_data_156; // @[hash.scala 94:22]
  reg [7:0] phv_data_157; // @[hash.scala 94:22]
  reg [7:0] phv_data_158; // @[hash.scala 94:22]
  reg [7:0] phv_data_159; // @[hash.scala 94:22]
  reg [15:0] phv_header_0; // @[hash.scala 94:22]
  reg [15:0] phv_header_1; // @[hash.scala 94:22]
  reg [15:0] phv_header_2; // @[hash.scala 94:22]
  reg [15:0] phv_header_3; // @[hash.scala 94:22]
  reg [15:0] phv_header_4; // @[hash.scala 94:22]
  reg [15:0] phv_header_5; // @[hash.scala 94:22]
  reg [15:0] phv_header_6; // @[hash.scala 94:22]
  reg [15:0] phv_header_7; // @[hash.scala 94:22]
  reg [15:0] phv_header_8; // @[hash.scala 94:22]
  reg [15:0] phv_header_9; // @[hash.scala 94:22]
  reg [15:0] phv_header_10; // @[hash.scala 94:22]
  reg [15:0] phv_header_11; // @[hash.scala 94:22]
  reg [15:0] phv_header_12; // @[hash.scala 94:22]
  reg [15:0] phv_header_13; // @[hash.scala 94:22]
  reg [15:0] phv_header_14; // @[hash.scala 94:22]
  reg [15:0] phv_header_15; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_state; // @[hash.scala 94:22]
  reg [7:0] phv_parse_current_offset; // @[hash.scala 94:22]
  reg [15:0] phv_parse_transition_field; // @[hash.scala 94:22]
  reg [3:0] phv_next_processor_id; // @[hash.scala 94:22]
  reg  phv_next_config_id; // @[hash.scala 94:22]
  reg  phv_is_valid_processor; // @[hash.scala 94:22]
  reg [191:0] key; // @[hash.scala 98:22]
  reg [15:0] sum; // @[hash.scala 102:22]
  reg [3:0] hash_depth; // @[hash.scala 106:29]
  reg [15:0] hash_val; // @[hash.scala 108:27]
  wire [15:0] _GEN_5 = {{3'd0}, sum[12:0]}; // @[hash.scala 116:44]
  wire [15:0] _io_val_out_T_2 = hash_val + _GEN_5; // @[hash.scala 116:44]
  wire [15:0] _GEN_2 = hash_depth[3] ? _io_val_out_T_2 : hash_val; // @[hash.scala 115:42 hash.scala 116:32 hash.scala 118:32]
  wire [15:0] _GEN_3 = hash_depth == 4'h0 ? sum : _GEN_2; // @[hash.scala 112:71 hash.scala 113:28]
  assign io_pipe_phv_out_data_0 = phv_data_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_1 = phv_data_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_2 = phv_data_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_3 = phv_data_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_4 = phv_data_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_5 = phv_data_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_6 = phv_data_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_7 = phv_data_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_8 = phv_data_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_9 = phv_data_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_10 = phv_data_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_11 = phv_data_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_12 = phv_data_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_13 = phv_data_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_14 = phv_data_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_15 = phv_data_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_16 = phv_data_16; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_17 = phv_data_17; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_18 = phv_data_18; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_19 = phv_data_19; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_20 = phv_data_20; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_21 = phv_data_21; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_22 = phv_data_22; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_23 = phv_data_23; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_24 = phv_data_24; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_25 = phv_data_25; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_26 = phv_data_26; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_27 = phv_data_27; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_28 = phv_data_28; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_29 = phv_data_29; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_30 = phv_data_30; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_31 = phv_data_31; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_32 = phv_data_32; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_33 = phv_data_33; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_34 = phv_data_34; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_35 = phv_data_35; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_36 = phv_data_36; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_37 = phv_data_37; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_38 = phv_data_38; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_39 = phv_data_39; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_40 = phv_data_40; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_41 = phv_data_41; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_42 = phv_data_42; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_43 = phv_data_43; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_44 = phv_data_44; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_45 = phv_data_45; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_46 = phv_data_46; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_47 = phv_data_47; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_48 = phv_data_48; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_49 = phv_data_49; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_50 = phv_data_50; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_51 = phv_data_51; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_52 = phv_data_52; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_53 = phv_data_53; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_54 = phv_data_54; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_55 = phv_data_55; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_56 = phv_data_56; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_57 = phv_data_57; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_58 = phv_data_58; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_59 = phv_data_59; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_60 = phv_data_60; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_61 = phv_data_61; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_62 = phv_data_62; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_63 = phv_data_63; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_64 = phv_data_64; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_65 = phv_data_65; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_66 = phv_data_66; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_67 = phv_data_67; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_68 = phv_data_68; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_69 = phv_data_69; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_70 = phv_data_70; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_71 = phv_data_71; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_72 = phv_data_72; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_73 = phv_data_73; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_74 = phv_data_74; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_75 = phv_data_75; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_76 = phv_data_76; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_77 = phv_data_77; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_78 = phv_data_78; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_79 = phv_data_79; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_80 = phv_data_80; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_81 = phv_data_81; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_82 = phv_data_82; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_83 = phv_data_83; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_84 = phv_data_84; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_85 = phv_data_85; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_86 = phv_data_86; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_87 = phv_data_87; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_88 = phv_data_88; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_89 = phv_data_89; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_90 = phv_data_90; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_91 = phv_data_91; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_92 = phv_data_92; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_93 = phv_data_93; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_94 = phv_data_94; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_95 = phv_data_95; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_96 = phv_data_96; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_97 = phv_data_97; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_98 = phv_data_98; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_99 = phv_data_99; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_100 = phv_data_100; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_101 = phv_data_101; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_102 = phv_data_102; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_103 = phv_data_103; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_104 = phv_data_104; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_105 = phv_data_105; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_106 = phv_data_106; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_107 = phv_data_107; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_108 = phv_data_108; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_109 = phv_data_109; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_110 = phv_data_110; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_111 = phv_data_111; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_112 = phv_data_112; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_113 = phv_data_113; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_114 = phv_data_114; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_115 = phv_data_115; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_116 = phv_data_116; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_117 = phv_data_117; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_118 = phv_data_118; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_119 = phv_data_119; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_120 = phv_data_120; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_121 = phv_data_121; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_122 = phv_data_122; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_123 = phv_data_123; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_124 = phv_data_124; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_125 = phv_data_125; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_126 = phv_data_126; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_127 = phv_data_127; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_128 = phv_data_128; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_129 = phv_data_129; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_130 = phv_data_130; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_131 = phv_data_131; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_132 = phv_data_132; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_133 = phv_data_133; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_134 = phv_data_134; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_135 = phv_data_135; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_136 = phv_data_136; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_137 = phv_data_137; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_138 = phv_data_138; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_139 = phv_data_139; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_140 = phv_data_140; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_141 = phv_data_141; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_142 = phv_data_142; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_143 = phv_data_143; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_144 = phv_data_144; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_145 = phv_data_145; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_146 = phv_data_146; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_147 = phv_data_147; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_148 = phv_data_148; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_149 = phv_data_149; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_150 = phv_data_150; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_151 = phv_data_151; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_152 = phv_data_152; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_153 = phv_data_153; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_154 = phv_data_154; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_155 = phv_data_155; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_156 = phv_data_156; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_157 = phv_data_157; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_158 = phv_data_158; // @[hash.scala 96:25]
  assign io_pipe_phv_out_data_159 = phv_data_159; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_0 = phv_header_0; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_1 = phv_header_1; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_2 = phv_header_2; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_3 = phv_header_3; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_4 = phv_header_4; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_5 = phv_header_5; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_6 = phv_header_6; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_7 = phv_header_7; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_8 = phv_header_8; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_9 = phv_header_9; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_10 = phv_header_10; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_11 = phv_header_11; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_12 = phv_header_12; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_13 = phv_header_13; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_14 = phv_header_14; // @[hash.scala 96:25]
  assign io_pipe_phv_out_header_15 = phv_header_15; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_state = phv_parse_current_state; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_current_offset = phv_parse_current_offset; // @[hash.scala 96:25]
  assign io_pipe_phv_out_parse_transition_field = phv_parse_transition_field; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_processor_id = phv_next_processor_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_next_config_id = phv_next_config_id; // @[hash.scala 96:25]
  assign io_pipe_phv_out_is_valid_processor = phv_is_valid_processor; // @[hash.scala 96:25]
  assign io_key_out = key; // @[hash.scala 100:20]
  assign io_sum_out = sum; // @[hash.scala 104:20]
  assign io_val_out = phv_is_valid_processor ? _GEN_3 : hash_val; // @[hash.scala 111:39 hash.scala 122:24]
  always @(posedge clock) begin
    phv_data_0 <= io_pipe_phv_in_data_0; // @[hash.scala 95:13]
    phv_data_1 <= io_pipe_phv_in_data_1; // @[hash.scala 95:13]
    phv_data_2 <= io_pipe_phv_in_data_2; // @[hash.scala 95:13]
    phv_data_3 <= io_pipe_phv_in_data_3; // @[hash.scala 95:13]
    phv_data_4 <= io_pipe_phv_in_data_4; // @[hash.scala 95:13]
    phv_data_5 <= io_pipe_phv_in_data_5; // @[hash.scala 95:13]
    phv_data_6 <= io_pipe_phv_in_data_6; // @[hash.scala 95:13]
    phv_data_7 <= io_pipe_phv_in_data_7; // @[hash.scala 95:13]
    phv_data_8 <= io_pipe_phv_in_data_8; // @[hash.scala 95:13]
    phv_data_9 <= io_pipe_phv_in_data_9; // @[hash.scala 95:13]
    phv_data_10 <= io_pipe_phv_in_data_10; // @[hash.scala 95:13]
    phv_data_11 <= io_pipe_phv_in_data_11; // @[hash.scala 95:13]
    phv_data_12 <= io_pipe_phv_in_data_12; // @[hash.scala 95:13]
    phv_data_13 <= io_pipe_phv_in_data_13; // @[hash.scala 95:13]
    phv_data_14 <= io_pipe_phv_in_data_14; // @[hash.scala 95:13]
    phv_data_15 <= io_pipe_phv_in_data_15; // @[hash.scala 95:13]
    phv_data_16 <= io_pipe_phv_in_data_16; // @[hash.scala 95:13]
    phv_data_17 <= io_pipe_phv_in_data_17; // @[hash.scala 95:13]
    phv_data_18 <= io_pipe_phv_in_data_18; // @[hash.scala 95:13]
    phv_data_19 <= io_pipe_phv_in_data_19; // @[hash.scala 95:13]
    phv_data_20 <= io_pipe_phv_in_data_20; // @[hash.scala 95:13]
    phv_data_21 <= io_pipe_phv_in_data_21; // @[hash.scala 95:13]
    phv_data_22 <= io_pipe_phv_in_data_22; // @[hash.scala 95:13]
    phv_data_23 <= io_pipe_phv_in_data_23; // @[hash.scala 95:13]
    phv_data_24 <= io_pipe_phv_in_data_24; // @[hash.scala 95:13]
    phv_data_25 <= io_pipe_phv_in_data_25; // @[hash.scala 95:13]
    phv_data_26 <= io_pipe_phv_in_data_26; // @[hash.scala 95:13]
    phv_data_27 <= io_pipe_phv_in_data_27; // @[hash.scala 95:13]
    phv_data_28 <= io_pipe_phv_in_data_28; // @[hash.scala 95:13]
    phv_data_29 <= io_pipe_phv_in_data_29; // @[hash.scala 95:13]
    phv_data_30 <= io_pipe_phv_in_data_30; // @[hash.scala 95:13]
    phv_data_31 <= io_pipe_phv_in_data_31; // @[hash.scala 95:13]
    phv_data_32 <= io_pipe_phv_in_data_32; // @[hash.scala 95:13]
    phv_data_33 <= io_pipe_phv_in_data_33; // @[hash.scala 95:13]
    phv_data_34 <= io_pipe_phv_in_data_34; // @[hash.scala 95:13]
    phv_data_35 <= io_pipe_phv_in_data_35; // @[hash.scala 95:13]
    phv_data_36 <= io_pipe_phv_in_data_36; // @[hash.scala 95:13]
    phv_data_37 <= io_pipe_phv_in_data_37; // @[hash.scala 95:13]
    phv_data_38 <= io_pipe_phv_in_data_38; // @[hash.scala 95:13]
    phv_data_39 <= io_pipe_phv_in_data_39; // @[hash.scala 95:13]
    phv_data_40 <= io_pipe_phv_in_data_40; // @[hash.scala 95:13]
    phv_data_41 <= io_pipe_phv_in_data_41; // @[hash.scala 95:13]
    phv_data_42 <= io_pipe_phv_in_data_42; // @[hash.scala 95:13]
    phv_data_43 <= io_pipe_phv_in_data_43; // @[hash.scala 95:13]
    phv_data_44 <= io_pipe_phv_in_data_44; // @[hash.scala 95:13]
    phv_data_45 <= io_pipe_phv_in_data_45; // @[hash.scala 95:13]
    phv_data_46 <= io_pipe_phv_in_data_46; // @[hash.scala 95:13]
    phv_data_47 <= io_pipe_phv_in_data_47; // @[hash.scala 95:13]
    phv_data_48 <= io_pipe_phv_in_data_48; // @[hash.scala 95:13]
    phv_data_49 <= io_pipe_phv_in_data_49; // @[hash.scala 95:13]
    phv_data_50 <= io_pipe_phv_in_data_50; // @[hash.scala 95:13]
    phv_data_51 <= io_pipe_phv_in_data_51; // @[hash.scala 95:13]
    phv_data_52 <= io_pipe_phv_in_data_52; // @[hash.scala 95:13]
    phv_data_53 <= io_pipe_phv_in_data_53; // @[hash.scala 95:13]
    phv_data_54 <= io_pipe_phv_in_data_54; // @[hash.scala 95:13]
    phv_data_55 <= io_pipe_phv_in_data_55; // @[hash.scala 95:13]
    phv_data_56 <= io_pipe_phv_in_data_56; // @[hash.scala 95:13]
    phv_data_57 <= io_pipe_phv_in_data_57; // @[hash.scala 95:13]
    phv_data_58 <= io_pipe_phv_in_data_58; // @[hash.scala 95:13]
    phv_data_59 <= io_pipe_phv_in_data_59; // @[hash.scala 95:13]
    phv_data_60 <= io_pipe_phv_in_data_60; // @[hash.scala 95:13]
    phv_data_61 <= io_pipe_phv_in_data_61; // @[hash.scala 95:13]
    phv_data_62 <= io_pipe_phv_in_data_62; // @[hash.scala 95:13]
    phv_data_63 <= io_pipe_phv_in_data_63; // @[hash.scala 95:13]
    phv_data_64 <= io_pipe_phv_in_data_64; // @[hash.scala 95:13]
    phv_data_65 <= io_pipe_phv_in_data_65; // @[hash.scala 95:13]
    phv_data_66 <= io_pipe_phv_in_data_66; // @[hash.scala 95:13]
    phv_data_67 <= io_pipe_phv_in_data_67; // @[hash.scala 95:13]
    phv_data_68 <= io_pipe_phv_in_data_68; // @[hash.scala 95:13]
    phv_data_69 <= io_pipe_phv_in_data_69; // @[hash.scala 95:13]
    phv_data_70 <= io_pipe_phv_in_data_70; // @[hash.scala 95:13]
    phv_data_71 <= io_pipe_phv_in_data_71; // @[hash.scala 95:13]
    phv_data_72 <= io_pipe_phv_in_data_72; // @[hash.scala 95:13]
    phv_data_73 <= io_pipe_phv_in_data_73; // @[hash.scala 95:13]
    phv_data_74 <= io_pipe_phv_in_data_74; // @[hash.scala 95:13]
    phv_data_75 <= io_pipe_phv_in_data_75; // @[hash.scala 95:13]
    phv_data_76 <= io_pipe_phv_in_data_76; // @[hash.scala 95:13]
    phv_data_77 <= io_pipe_phv_in_data_77; // @[hash.scala 95:13]
    phv_data_78 <= io_pipe_phv_in_data_78; // @[hash.scala 95:13]
    phv_data_79 <= io_pipe_phv_in_data_79; // @[hash.scala 95:13]
    phv_data_80 <= io_pipe_phv_in_data_80; // @[hash.scala 95:13]
    phv_data_81 <= io_pipe_phv_in_data_81; // @[hash.scala 95:13]
    phv_data_82 <= io_pipe_phv_in_data_82; // @[hash.scala 95:13]
    phv_data_83 <= io_pipe_phv_in_data_83; // @[hash.scala 95:13]
    phv_data_84 <= io_pipe_phv_in_data_84; // @[hash.scala 95:13]
    phv_data_85 <= io_pipe_phv_in_data_85; // @[hash.scala 95:13]
    phv_data_86 <= io_pipe_phv_in_data_86; // @[hash.scala 95:13]
    phv_data_87 <= io_pipe_phv_in_data_87; // @[hash.scala 95:13]
    phv_data_88 <= io_pipe_phv_in_data_88; // @[hash.scala 95:13]
    phv_data_89 <= io_pipe_phv_in_data_89; // @[hash.scala 95:13]
    phv_data_90 <= io_pipe_phv_in_data_90; // @[hash.scala 95:13]
    phv_data_91 <= io_pipe_phv_in_data_91; // @[hash.scala 95:13]
    phv_data_92 <= io_pipe_phv_in_data_92; // @[hash.scala 95:13]
    phv_data_93 <= io_pipe_phv_in_data_93; // @[hash.scala 95:13]
    phv_data_94 <= io_pipe_phv_in_data_94; // @[hash.scala 95:13]
    phv_data_95 <= io_pipe_phv_in_data_95; // @[hash.scala 95:13]
    phv_data_96 <= io_pipe_phv_in_data_96; // @[hash.scala 95:13]
    phv_data_97 <= io_pipe_phv_in_data_97; // @[hash.scala 95:13]
    phv_data_98 <= io_pipe_phv_in_data_98; // @[hash.scala 95:13]
    phv_data_99 <= io_pipe_phv_in_data_99; // @[hash.scala 95:13]
    phv_data_100 <= io_pipe_phv_in_data_100; // @[hash.scala 95:13]
    phv_data_101 <= io_pipe_phv_in_data_101; // @[hash.scala 95:13]
    phv_data_102 <= io_pipe_phv_in_data_102; // @[hash.scala 95:13]
    phv_data_103 <= io_pipe_phv_in_data_103; // @[hash.scala 95:13]
    phv_data_104 <= io_pipe_phv_in_data_104; // @[hash.scala 95:13]
    phv_data_105 <= io_pipe_phv_in_data_105; // @[hash.scala 95:13]
    phv_data_106 <= io_pipe_phv_in_data_106; // @[hash.scala 95:13]
    phv_data_107 <= io_pipe_phv_in_data_107; // @[hash.scala 95:13]
    phv_data_108 <= io_pipe_phv_in_data_108; // @[hash.scala 95:13]
    phv_data_109 <= io_pipe_phv_in_data_109; // @[hash.scala 95:13]
    phv_data_110 <= io_pipe_phv_in_data_110; // @[hash.scala 95:13]
    phv_data_111 <= io_pipe_phv_in_data_111; // @[hash.scala 95:13]
    phv_data_112 <= io_pipe_phv_in_data_112; // @[hash.scala 95:13]
    phv_data_113 <= io_pipe_phv_in_data_113; // @[hash.scala 95:13]
    phv_data_114 <= io_pipe_phv_in_data_114; // @[hash.scala 95:13]
    phv_data_115 <= io_pipe_phv_in_data_115; // @[hash.scala 95:13]
    phv_data_116 <= io_pipe_phv_in_data_116; // @[hash.scala 95:13]
    phv_data_117 <= io_pipe_phv_in_data_117; // @[hash.scala 95:13]
    phv_data_118 <= io_pipe_phv_in_data_118; // @[hash.scala 95:13]
    phv_data_119 <= io_pipe_phv_in_data_119; // @[hash.scala 95:13]
    phv_data_120 <= io_pipe_phv_in_data_120; // @[hash.scala 95:13]
    phv_data_121 <= io_pipe_phv_in_data_121; // @[hash.scala 95:13]
    phv_data_122 <= io_pipe_phv_in_data_122; // @[hash.scala 95:13]
    phv_data_123 <= io_pipe_phv_in_data_123; // @[hash.scala 95:13]
    phv_data_124 <= io_pipe_phv_in_data_124; // @[hash.scala 95:13]
    phv_data_125 <= io_pipe_phv_in_data_125; // @[hash.scala 95:13]
    phv_data_126 <= io_pipe_phv_in_data_126; // @[hash.scala 95:13]
    phv_data_127 <= io_pipe_phv_in_data_127; // @[hash.scala 95:13]
    phv_data_128 <= io_pipe_phv_in_data_128; // @[hash.scala 95:13]
    phv_data_129 <= io_pipe_phv_in_data_129; // @[hash.scala 95:13]
    phv_data_130 <= io_pipe_phv_in_data_130; // @[hash.scala 95:13]
    phv_data_131 <= io_pipe_phv_in_data_131; // @[hash.scala 95:13]
    phv_data_132 <= io_pipe_phv_in_data_132; // @[hash.scala 95:13]
    phv_data_133 <= io_pipe_phv_in_data_133; // @[hash.scala 95:13]
    phv_data_134 <= io_pipe_phv_in_data_134; // @[hash.scala 95:13]
    phv_data_135 <= io_pipe_phv_in_data_135; // @[hash.scala 95:13]
    phv_data_136 <= io_pipe_phv_in_data_136; // @[hash.scala 95:13]
    phv_data_137 <= io_pipe_phv_in_data_137; // @[hash.scala 95:13]
    phv_data_138 <= io_pipe_phv_in_data_138; // @[hash.scala 95:13]
    phv_data_139 <= io_pipe_phv_in_data_139; // @[hash.scala 95:13]
    phv_data_140 <= io_pipe_phv_in_data_140; // @[hash.scala 95:13]
    phv_data_141 <= io_pipe_phv_in_data_141; // @[hash.scala 95:13]
    phv_data_142 <= io_pipe_phv_in_data_142; // @[hash.scala 95:13]
    phv_data_143 <= io_pipe_phv_in_data_143; // @[hash.scala 95:13]
    phv_data_144 <= io_pipe_phv_in_data_144; // @[hash.scala 95:13]
    phv_data_145 <= io_pipe_phv_in_data_145; // @[hash.scala 95:13]
    phv_data_146 <= io_pipe_phv_in_data_146; // @[hash.scala 95:13]
    phv_data_147 <= io_pipe_phv_in_data_147; // @[hash.scala 95:13]
    phv_data_148 <= io_pipe_phv_in_data_148; // @[hash.scala 95:13]
    phv_data_149 <= io_pipe_phv_in_data_149; // @[hash.scala 95:13]
    phv_data_150 <= io_pipe_phv_in_data_150; // @[hash.scala 95:13]
    phv_data_151 <= io_pipe_phv_in_data_151; // @[hash.scala 95:13]
    phv_data_152 <= io_pipe_phv_in_data_152; // @[hash.scala 95:13]
    phv_data_153 <= io_pipe_phv_in_data_153; // @[hash.scala 95:13]
    phv_data_154 <= io_pipe_phv_in_data_154; // @[hash.scala 95:13]
    phv_data_155 <= io_pipe_phv_in_data_155; // @[hash.scala 95:13]
    phv_data_156 <= io_pipe_phv_in_data_156; // @[hash.scala 95:13]
    phv_data_157 <= io_pipe_phv_in_data_157; // @[hash.scala 95:13]
    phv_data_158 <= io_pipe_phv_in_data_158; // @[hash.scala 95:13]
    phv_data_159 <= io_pipe_phv_in_data_159; // @[hash.scala 95:13]
    phv_header_0 <= io_pipe_phv_in_header_0; // @[hash.scala 95:13]
    phv_header_1 <= io_pipe_phv_in_header_1; // @[hash.scala 95:13]
    phv_header_2 <= io_pipe_phv_in_header_2; // @[hash.scala 95:13]
    phv_header_3 <= io_pipe_phv_in_header_3; // @[hash.scala 95:13]
    phv_header_4 <= io_pipe_phv_in_header_4; // @[hash.scala 95:13]
    phv_header_5 <= io_pipe_phv_in_header_5; // @[hash.scala 95:13]
    phv_header_6 <= io_pipe_phv_in_header_6; // @[hash.scala 95:13]
    phv_header_7 <= io_pipe_phv_in_header_7; // @[hash.scala 95:13]
    phv_header_8 <= io_pipe_phv_in_header_8; // @[hash.scala 95:13]
    phv_header_9 <= io_pipe_phv_in_header_9; // @[hash.scala 95:13]
    phv_header_10 <= io_pipe_phv_in_header_10; // @[hash.scala 95:13]
    phv_header_11 <= io_pipe_phv_in_header_11; // @[hash.scala 95:13]
    phv_header_12 <= io_pipe_phv_in_header_12; // @[hash.scala 95:13]
    phv_header_13 <= io_pipe_phv_in_header_13; // @[hash.scala 95:13]
    phv_header_14 <= io_pipe_phv_in_header_14; // @[hash.scala 95:13]
    phv_header_15 <= io_pipe_phv_in_header_15; // @[hash.scala 95:13]
    phv_parse_current_state <= io_pipe_phv_in_parse_current_state; // @[hash.scala 95:13]
    phv_parse_current_offset <= io_pipe_phv_in_parse_current_offset; // @[hash.scala 95:13]
    phv_parse_transition_field <= io_pipe_phv_in_parse_transition_field; // @[hash.scala 95:13]
    phv_next_processor_id <= io_pipe_phv_in_next_processor_id; // @[hash.scala 95:13]
    phv_next_config_id <= io_pipe_phv_in_next_config_id; // @[hash.scala 95:13]
    phv_is_valid_processor <= io_pipe_phv_in_is_valid_processor; // @[hash.scala 95:13]
    key <= io_key_in; // @[hash.scala 99:13]
    sum <= io_sum_in; // @[hash.scala 103:13]
    if (io_pipe_phv_in_next_config_id) begin // @[hash.scala 107:20]
      hash_depth <= io_hash_depth_1; // @[hash.scala 107:20]
    end else begin
      hash_depth <= io_hash_depth_0;
    end
    hash_val <= io_val_in; // @[hash.scala 109:18]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phv_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  phv_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  phv_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  phv_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  phv_data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  phv_data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  phv_data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  phv_data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  phv_data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  phv_data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  phv_data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  phv_data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  phv_data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  phv_data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  phv_data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  phv_data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  phv_data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  phv_data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  phv_data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  phv_data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  phv_data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  phv_data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  phv_data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  phv_data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  phv_data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  phv_data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  phv_data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  phv_data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  phv_data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  phv_data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  phv_data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  phv_data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  phv_data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  phv_data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  phv_data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  phv_data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  phv_data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  phv_data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  phv_data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  phv_data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  phv_data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  phv_data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  phv_data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  phv_data_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  phv_data_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  phv_data_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  phv_data_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  phv_data_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  phv_data_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  phv_data_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  phv_data_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  phv_data_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  phv_data_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  phv_data_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  phv_data_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  phv_data_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  phv_data_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  phv_data_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  phv_data_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  phv_data_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  phv_data_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  phv_data_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  phv_data_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  phv_data_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  phv_data_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  phv_data_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  phv_data_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  phv_data_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  phv_data_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  phv_data_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  phv_data_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  phv_data_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  phv_data_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  phv_data_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  phv_data_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  phv_data_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  phv_data_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  phv_data_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  phv_data_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  phv_data_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  phv_data_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  phv_data_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  phv_data_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  phv_data_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  phv_data_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  phv_data_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  phv_data_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  phv_data_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  phv_data_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  phv_data_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  phv_data_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  phv_data_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  phv_data_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  phv_data_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  phv_data_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  phv_data_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  phv_data_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  phv_data_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  phv_data_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  phv_data_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  phv_data_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  phv_data_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  phv_data_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  phv_data_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  phv_data_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  phv_data_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  phv_data_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  phv_data_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  phv_data_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  phv_data_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  phv_data_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  phv_data_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  phv_data_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  phv_data_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  phv_data_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  phv_data_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  phv_data_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  phv_data_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  phv_data_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  phv_data_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  phv_data_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  phv_data_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  phv_data_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  phv_data_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  phv_data_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  phv_data_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  phv_data_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  phv_data_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  phv_data_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  phv_data_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  phv_data_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  phv_data_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  phv_data_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  phv_data_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  phv_data_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  phv_data_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  phv_data_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  phv_data_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  phv_data_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  phv_data_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  phv_data_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  phv_data_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  phv_data_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  phv_data_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  phv_data_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  phv_data_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  phv_data_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  phv_data_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  phv_data_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  phv_data_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  phv_data_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  phv_data_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  phv_data_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  phv_data_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  phv_data_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  phv_data_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  phv_data_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  phv_data_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  phv_data_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  phv_data_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  phv_header_0 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  phv_header_1 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  phv_header_2 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  phv_header_3 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  phv_header_4 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  phv_header_5 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  phv_header_6 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  phv_header_7 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  phv_header_8 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  phv_header_9 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  phv_header_10 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  phv_header_11 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  phv_header_12 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  phv_header_13 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  phv_header_14 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  phv_header_15 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  phv_parse_current_state = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  phv_parse_current_offset = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  phv_parse_transition_field = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  phv_next_processor_id = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  phv_next_config_id = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  phv_is_valid_processor = _RAND_181[0:0];
  _RAND_182 = {6{`RANDOM}};
  key = _RAND_182[191:0];
  _RAND_183 = {1{`RANDOM}};
  sum = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  hash_depth = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  hash_val = _RAND_185[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Hash(
  input          clock,
  input          reset,
  input  [7:0]   io_pipe_phv_in_data_0,
  input  [7:0]   io_pipe_phv_in_data_1,
  input  [7:0]   io_pipe_phv_in_data_2,
  input  [7:0]   io_pipe_phv_in_data_3,
  input  [7:0]   io_pipe_phv_in_data_4,
  input  [7:0]   io_pipe_phv_in_data_5,
  input  [7:0]   io_pipe_phv_in_data_6,
  input  [7:0]   io_pipe_phv_in_data_7,
  input  [7:0]   io_pipe_phv_in_data_8,
  input  [7:0]   io_pipe_phv_in_data_9,
  input  [7:0]   io_pipe_phv_in_data_10,
  input  [7:0]   io_pipe_phv_in_data_11,
  input  [7:0]   io_pipe_phv_in_data_12,
  input  [7:0]   io_pipe_phv_in_data_13,
  input  [7:0]   io_pipe_phv_in_data_14,
  input  [7:0]   io_pipe_phv_in_data_15,
  input  [7:0]   io_pipe_phv_in_data_16,
  input  [7:0]   io_pipe_phv_in_data_17,
  input  [7:0]   io_pipe_phv_in_data_18,
  input  [7:0]   io_pipe_phv_in_data_19,
  input  [7:0]   io_pipe_phv_in_data_20,
  input  [7:0]   io_pipe_phv_in_data_21,
  input  [7:0]   io_pipe_phv_in_data_22,
  input  [7:0]   io_pipe_phv_in_data_23,
  input  [7:0]   io_pipe_phv_in_data_24,
  input  [7:0]   io_pipe_phv_in_data_25,
  input  [7:0]   io_pipe_phv_in_data_26,
  input  [7:0]   io_pipe_phv_in_data_27,
  input  [7:0]   io_pipe_phv_in_data_28,
  input  [7:0]   io_pipe_phv_in_data_29,
  input  [7:0]   io_pipe_phv_in_data_30,
  input  [7:0]   io_pipe_phv_in_data_31,
  input  [7:0]   io_pipe_phv_in_data_32,
  input  [7:0]   io_pipe_phv_in_data_33,
  input  [7:0]   io_pipe_phv_in_data_34,
  input  [7:0]   io_pipe_phv_in_data_35,
  input  [7:0]   io_pipe_phv_in_data_36,
  input  [7:0]   io_pipe_phv_in_data_37,
  input  [7:0]   io_pipe_phv_in_data_38,
  input  [7:0]   io_pipe_phv_in_data_39,
  input  [7:0]   io_pipe_phv_in_data_40,
  input  [7:0]   io_pipe_phv_in_data_41,
  input  [7:0]   io_pipe_phv_in_data_42,
  input  [7:0]   io_pipe_phv_in_data_43,
  input  [7:0]   io_pipe_phv_in_data_44,
  input  [7:0]   io_pipe_phv_in_data_45,
  input  [7:0]   io_pipe_phv_in_data_46,
  input  [7:0]   io_pipe_phv_in_data_47,
  input  [7:0]   io_pipe_phv_in_data_48,
  input  [7:0]   io_pipe_phv_in_data_49,
  input  [7:0]   io_pipe_phv_in_data_50,
  input  [7:0]   io_pipe_phv_in_data_51,
  input  [7:0]   io_pipe_phv_in_data_52,
  input  [7:0]   io_pipe_phv_in_data_53,
  input  [7:0]   io_pipe_phv_in_data_54,
  input  [7:0]   io_pipe_phv_in_data_55,
  input  [7:0]   io_pipe_phv_in_data_56,
  input  [7:0]   io_pipe_phv_in_data_57,
  input  [7:0]   io_pipe_phv_in_data_58,
  input  [7:0]   io_pipe_phv_in_data_59,
  input  [7:0]   io_pipe_phv_in_data_60,
  input  [7:0]   io_pipe_phv_in_data_61,
  input  [7:0]   io_pipe_phv_in_data_62,
  input  [7:0]   io_pipe_phv_in_data_63,
  input  [7:0]   io_pipe_phv_in_data_64,
  input  [7:0]   io_pipe_phv_in_data_65,
  input  [7:0]   io_pipe_phv_in_data_66,
  input  [7:0]   io_pipe_phv_in_data_67,
  input  [7:0]   io_pipe_phv_in_data_68,
  input  [7:0]   io_pipe_phv_in_data_69,
  input  [7:0]   io_pipe_phv_in_data_70,
  input  [7:0]   io_pipe_phv_in_data_71,
  input  [7:0]   io_pipe_phv_in_data_72,
  input  [7:0]   io_pipe_phv_in_data_73,
  input  [7:0]   io_pipe_phv_in_data_74,
  input  [7:0]   io_pipe_phv_in_data_75,
  input  [7:0]   io_pipe_phv_in_data_76,
  input  [7:0]   io_pipe_phv_in_data_77,
  input  [7:0]   io_pipe_phv_in_data_78,
  input  [7:0]   io_pipe_phv_in_data_79,
  input  [7:0]   io_pipe_phv_in_data_80,
  input  [7:0]   io_pipe_phv_in_data_81,
  input  [7:0]   io_pipe_phv_in_data_82,
  input  [7:0]   io_pipe_phv_in_data_83,
  input  [7:0]   io_pipe_phv_in_data_84,
  input  [7:0]   io_pipe_phv_in_data_85,
  input  [7:0]   io_pipe_phv_in_data_86,
  input  [7:0]   io_pipe_phv_in_data_87,
  input  [7:0]   io_pipe_phv_in_data_88,
  input  [7:0]   io_pipe_phv_in_data_89,
  input  [7:0]   io_pipe_phv_in_data_90,
  input  [7:0]   io_pipe_phv_in_data_91,
  input  [7:0]   io_pipe_phv_in_data_92,
  input  [7:0]   io_pipe_phv_in_data_93,
  input  [7:0]   io_pipe_phv_in_data_94,
  input  [7:0]   io_pipe_phv_in_data_95,
  input  [7:0]   io_pipe_phv_in_data_96,
  input  [7:0]   io_pipe_phv_in_data_97,
  input  [7:0]   io_pipe_phv_in_data_98,
  input  [7:0]   io_pipe_phv_in_data_99,
  input  [7:0]   io_pipe_phv_in_data_100,
  input  [7:0]   io_pipe_phv_in_data_101,
  input  [7:0]   io_pipe_phv_in_data_102,
  input  [7:0]   io_pipe_phv_in_data_103,
  input  [7:0]   io_pipe_phv_in_data_104,
  input  [7:0]   io_pipe_phv_in_data_105,
  input  [7:0]   io_pipe_phv_in_data_106,
  input  [7:0]   io_pipe_phv_in_data_107,
  input  [7:0]   io_pipe_phv_in_data_108,
  input  [7:0]   io_pipe_phv_in_data_109,
  input  [7:0]   io_pipe_phv_in_data_110,
  input  [7:0]   io_pipe_phv_in_data_111,
  input  [7:0]   io_pipe_phv_in_data_112,
  input  [7:0]   io_pipe_phv_in_data_113,
  input  [7:0]   io_pipe_phv_in_data_114,
  input  [7:0]   io_pipe_phv_in_data_115,
  input  [7:0]   io_pipe_phv_in_data_116,
  input  [7:0]   io_pipe_phv_in_data_117,
  input  [7:0]   io_pipe_phv_in_data_118,
  input  [7:0]   io_pipe_phv_in_data_119,
  input  [7:0]   io_pipe_phv_in_data_120,
  input  [7:0]   io_pipe_phv_in_data_121,
  input  [7:0]   io_pipe_phv_in_data_122,
  input  [7:0]   io_pipe_phv_in_data_123,
  input  [7:0]   io_pipe_phv_in_data_124,
  input  [7:0]   io_pipe_phv_in_data_125,
  input  [7:0]   io_pipe_phv_in_data_126,
  input  [7:0]   io_pipe_phv_in_data_127,
  input  [7:0]   io_pipe_phv_in_data_128,
  input  [7:0]   io_pipe_phv_in_data_129,
  input  [7:0]   io_pipe_phv_in_data_130,
  input  [7:0]   io_pipe_phv_in_data_131,
  input  [7:0]   io_pipe_phv_in_data_132,
  input  [7:0]   io_pipe_phv_in_data_133,
  input  [7:0]   io_pipe_phv_in_data_134,
  input  [7:0]   io_pipe_phv_in_data_135,
  input  [7:0]   io_pipe_phv_in_data_136,
  input  [7:0]   io_pipe_phv_in_data_137,
  input  [7:0]   io_pipe_phv_in_data_138,
  input  [7:0]   io_pipe_phv_in_data_139,
  input  [7:0]   io_pipe_phv_in_data_140,
  input  [7:0]   io_pipe_phv_in_data_141,
  input  [7:0]   io_pipe_phv_in_data_142,
  input  [7:0]   io_pipe_phv_in_data_143,
  input  [7:0]   io_pipe_phv_in_data_144,
  input  [7:0]   io_pipe_phv_in_data_145,
  input  [7:0]   io_pipe_phv_in_data_146,
  input  [7:0]   io_pipe_phv_in_data_147,
  input  [7:0]   io_pipe_phv_in_data_148,
  input  [7:0]   io_pipe_phv_in_data_149,
  input  [7:0]   io_pipe_phv_in_data_150,
  input  [7:0]   io_pipe_phv_in_data_151,
  input  [7:0]   io_pipe_phv_in_data_152,
  input  [7:0]   io_pipe_phv_in_data_153,
  input  [7:0]   io_pipe_phv_in_data_154,
  input  [7:0]   io_pipe_phv_in_data_155,
  input  [7:0]   io_pipe_phv_in_data_156,
  input  [7:0]   io_pipe_phv_in_data_157,
  input  [7:0]   io_pipe_phv_in_data_158,
  input  [7:0]   io_pipe_phv_in_data_159,
  input  [15:0]  io_pipe_phv_in_header_0,
  input  [15:0]  io_pipe_phv_in_header_1,
  input  [15:0]  io_pipe_phv_in_header_2,
  input  [15:0]  io_pipe_phv_in_header_3,
  input  [15:0]  io_pipe_phv_in_header_4,
  input  [15:0]  io_pipe_phv_in_header_5,
  input  [15:0]  io_pipe_phv_in_header_6,
  input  [15:0]  io_pipe_phv_in_header_7,
  input  [15:0]  io_pipe_phv_in_header_8,
  input  [15:0]  io_pipe_phv_in_header_9,
  input  [15:0]  io_pipe_phv_in_header_10,
  input  [15:0]  io_pipe_phv_in_header_11,
  input  [15:0]  io_pipe_phv_in_header_12,
  input  [15:0]  io_pipe_phv_in_header_13,
  input  [15:0]  io_pipe_phv_in_header_14,
  input  [15:0]  io_pipe_phv_in_header_15,
  input  [7:0]   io_pipe_phv_in_parse_current_state,
  input  [7:0]   io_pipe_phv_in_parse_current_offset,
  input  [15:0]  io_pipe_phv_in_parse_transition_field,
  input  [3:0]   io_pipe_phv_in_next_processor_id,
  input          io_pipe_phv_in_next_config_id,
  input          io_pipe_phv_in_is_valid_processor,
  output [7:0]   io_pipe_phv_out_data_0,
  output [7:0]   io_pipe_phv_out_data_1,
  output [7:0]   io_pipe_phv_out_data_2,
  output [7:0]   io_pipe_phv_out_data_3,
  output [7:0]   io_pipe_phv_out_data_4,
  output [7:0]   io_pipe_phv_out_data_5,
  output [7:0]   io_pipe_phv_out_data_6,
  output [7:0]   io_pipe_phv_out_data_7,
  output [7:0]   io_pipe_phv_out_data_8,
  output [7:0]   io_pipe_phv_out_data_9,
  output [7:0]   io_pipe_phv_out_data_10,
  output [7:0]   io_pipe_phv_out_data_11,
  output [7:0]   io_pipe_phv_out_data_12,
  output [7:0]   io_pipe_phv_out_data_13,
  output [7:0]   io_pipe_phv_out_data_14,
  output [7:0]   io_pipe_phv_out_data_15,
  output [7:0]   io_pipe_phv_out_data_16,
  output [7:0]   io_pipe_phv_out_data_17,
  output [7:0]   io_pipe_phv_out_data_18,
  output [7:0]   io_pipe_phv_out_data_19,
  output [7:0]   io_pipe_phv_out_data_20,
  output [7:0]   io_pipe_phv_out_data_21,
  output [7:0]   io_pipe_phv_out_data_22,
  output [7:0]   io_pipe_phv_out_data_23,
  output [7:0]   io_pipe_phv_out_data_24,
  output [7:0]   io_pipe_phv_out_data_25,
  output [7:0]   io_pipe_phv_out_data_26,
  output [7:0]   io_pipe_phv_out_data_27,
  output [7:0]   io_pipe_phv_out_data_28,
  output [7:0]   io_pipe_phv_out_data_29,
  output [7:0]   io_pipe_phv_out_data_30,
  output [7:0]   io_pipe_phv_out_data_31,
  output [7:0]   io_pipe_phv_out_data_32,
  output [7:0]   io_pipe_phv_out_data_33,
  output [7:0]   io_pipe_phv_out_data_34,
  output [7:0]   io_pipe_phv_out_data_35,
  output [7:0]   io_pipe_phv_out_data_36,
  output [7:0]   io_pipe_phv_out_data_37,
  output [7:0]   io_pipe_phv_out_data_38,
  output [7:0]   io_pipe_phv_out_data_39,
  output [7:0]   io_pipe_phv_out_data_40,
  output [7:0]   io_pipe_phv_out_data_41,
  output [7:0]   io_pipe_phv_out_data_42,
  output [7:0]   io_pipe_phv_out_data_43,
  output [7:0]   io_pipe_phv_out_data_44,
  output [7:0]   io_pipe_phv_out_data_45,
  output [7:0]   io_pipe_phv_out_data_46,
  output [7:0]   io_pipe_phv_out_data_47,
  output [7:0]   io_pipe_phv_out_data_48,
  output [7:0]   io_pipe_phv_out_data_49,
  output [7:0]   io_pipe_phv_out_data_50,
  output [7:0]   io_pipe_phv_out_data_51,
  output [7:0]   io_pipe_phv_out_data_52,
  output [7:0]   io_pipe_phv_out_data_53,
  output [7:0]   io_pipe_phv_out_data_54,
  output [7:0]   io_pipe_phv_out_data_55,
  output [7:0]   io_pipe_phv_out_data_56,
  output [7:0]   io_pipe_phv_out_data_57,
  output [7:0]   io_pipe_phv_out_data_58,
  output [7:0]   io_pipe_phv_out_data_59,
  output [7:0]   io_pipe_phv_out_data_60,
  output [7:0]   io_pipe_phv_out_data_61,
  output [7:0]   io_pipe_phv_out_data_62,
  output [7:0]   io_pipe_phv_out_data_63,
  output [7:0]   io_pipe_phv_out_data_64,
  output [7:0]   io_pipe_phv_out_data_65,
  output [7:0]   io_pipe_phv_out_data_66,
  output [7:0]   io_pipe_phv_out_data_67,
  output [7:0]   io_pipe_phv_out_data_68,
  output [7:0]   io_pipe_phv_out_data_69,
  output [7:0]   io_pipe_phv_out_data_70,
  output [7:0]   io_pipe_phv_out_data_71,
  output [7:0]   io_pipe_phv_out_data_72,
  output [7:0]   io_pipe_phv_out_data_73,
  output [7:0]   io_pipe_phv_out_data_74,
  output [7:0]   io_pipe_phv_out_data_75,
  output [7:0]   io_pipe_phv_out_data_76,
  output [7:0]   io_pipe_phv_out_data_77,
  output [7:0]   io_pipe_phv_out_data_78,
  output [7:0]   io_pipe_phv_out_data_79,
  output [7:0]   io_pipe_phv_out_data_80,
  output [7:0]   io_pipe_phv_out_data_81,
  output [7:0]   io_pipe_phv_out_data_82,
  output [7:0]   io_pipe_phv_out_data_83,
  output [7:0]   io_pipe_phv_out_data_84,
  output [7:0]   io_pipe_phv_out_data_85,
  output [7:0]   io_pipe_phv_out_data_86,
  output [7:0]   io_pipe_phv_out_data_87,
  output [7:0]   io_pipe_phv_out_data_88,
  output [7:0]   io_pipe_phv_out_data_89,
  output [7:0]   io_pipe_phv_out_data_90,
  output [7:0]   io_pipe_phv_out_data_91,
  output [7:0]   io_pipe_phv_out_data_92,
  output [7:0]   io_pipe_phv_out_data_93,
  output [7:0]   io_pipe_phv_out_data_94,
  output [7:0]   io_pipe_phv_out_data_95,
  output [7:0]   io_pipe_phv_out_data_96,
  output [7:0]   io_pipe_phv_out_data_97,
  output [7:0]   io_pipe_phv_out_data_98,
  output [7:0]   io_pipe_phv_out_data_99,
  output [7:0]   io_pipe_phv_out_data_100,
  output [7:0]   io_pipe_phv_out_data_101,
  output [7:0]   io_pipe_phv_out_data_102,
  output [7:0]   io_pipe_phv_out_data_103,
  output [7:0]   io_pipe_phv_out_data_104,
  output [7:0]   io_pipe_phv_out_data_105,
  output [7:0]   io_pipe_phv_out_data_106,
  output [7:0]   io_pipe_phv_out_data_107,
  output [7:0]   io_pipe_phv_out_data_108,
  output [7:0]   io_pipe_phv_out_data_109,
  output [7:0]   io_pipe_phv_out_data_110,
  output [7:0]   io_pipe_phv_out_data_111,
  output [7:0]   io_pipe_phv_out_data_112,
  output [7:0]   io_pipe_phv_out_data_113,
  output [7:0]   io_pipe_phv_out_data_114,
  output [7:0]   io_pipe_phv_out_data_115,
  output [7:0]   io_pipe_phv_out_data_116,
  output [7:0]   io_pipe_phv_out_data_117,
  output [7:0]   io_pipe_phv_out_data_118,
  output [7:0]   io_pipe_phv_out_data_119,
  output [7:0]   io_pipe_phv_out_data_120,
  output [7:0]   io_pipe_phv_out_data_121,
  output [7:0]   io_pipe_phv_out_data_122,
  output [7:0]   io_pipe_phv_out_data_123,
  output [7:0]   io_pipe_phv_out_data_124,
  output [7:0]   io_pipe_phv_out_data_125,
  output [7:0]   io_pipe_phv_out_data_126,
  output [7:0]   io_pipe_phv_out_data_127,
  output [7:0]   io_pipe_phv_out_data_128,
  output [7:0]   io_pipe_phv_out_data_129,
  output [7:0]   io_pipe_phv_out_data_130,
  output [7:0]   io_pipe_phv_out_data_131,
  output [7:0]   io_pipe_phv_out_data_132,
  output [7:0]   io_pipe_phv_out_data_133,
  output [7:0]   io_pipe_phv_out_data_134,
  output [7:0]   io_pipe_phv_out_data_135,
  output [7:0]   io_pipe_phv_out_data_136,
  output [7:0]   io_pipe_phv_out_data_137,
  output [7:0]   io_pipe_phv_out_data_138,
  output [7:0]   io_pipe_phv_out_data_139,
  output [7:0]   io_pipe_phv_out_data_140,
  output [7:0]   io_pipe_phv_out_data_141,
  output [7:0]   io_pipe_phv_out_data_142,
  output [7:0]   io_pipe_phv_out_data_143,
  output [7:0]   io_pipe_phv_out_data_144,
  output [7:0]   io_pipe_phv_out_data_145,
  output [7:0]   io_pipe_phv_out_data_146,
  output [7:0]   io_pipe_phv_out_data_147,
  output [7:0]   io_pipe_phv_out_data_148,
  output [7:0]   io_pipe_phv_out_data_149,
  output [7:0]   io_pipe_phv_out_data_150,
  output [7:0]   io_pipe_phv_out_data_151,
  output [7:0]   io_pipe_phv_out_data_152,
  output [7:0]   io_pipe_phv_out_data_153,
  output [7:0]   io_pipe_phv_out_data_154,
  output [7:0]   io_pipe_phv_out_data_155,
  output [7:0]   io_pipe_phv_out_data_156,
  output [7:0]   io_pipe_phv_out_data_157,
  output [7:0]   io_pipe_phv_out_data_158,
  output [7:0]   io_pipe_phv_out_data_159,
  output [15:0]  io_pipe_phv_out_header_0,
  output [15:0]  io_pipe_phv_out_header_1,
  output [15:0]  io_pipe_phv_out_header_2,
  output [15:0]  io_pipe_phv_out_header_3,
  output [15:0]  io_pipe_phv_out_header_4,
  output [15:0]  io_pipe_phv_out_header_5,
  output [15:0]  io_pipe_phv_out_header_6,
  output [15:0]  io_pipe_phv_out_header_7,
  output [15:0]  io_pipe_phv_out_header_8,
  output [15:0]  io_pipe_phv_out_header_9,
  output [15:0]  io_pipe_phv_out_header_10,
  output [15:0]  io_pipe_phv_out_header_11,
  output [15:0]  io_pipe_phv_out_header_12,
  output [15:0]  io_pipe_phv_out_header_13,
  output [15:0]  io_pipe_phv_out_header_14,
  output [15:0]  io_pipe_phv_out_header_15,
  output [7:0]   io_pipe_phv_out_parse_current_state,
  output [7:0]   io_pipe_phv_out_parse_current_offset,
  output [15:0]  io_pipe_phv_out_parse_transition_field,
  output [3:0]   io_pipe_phv_out_next_processor_id,
  output         io_pipe_phv_out_next_config_id,
  output         io_pipe_phv_out_is_valid_processor,
  input          io_mod_hash_depth_mod,
  input          io_mod_config_id,
  input  [3:0]   io_mod_hash_depth,
  input  [191:0] io_key_in,
  output [191:0] io_key_out,
  output [7:0]   io_hash_val,
  output [3:0]   io_hash_val_cs
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pipe1_clock; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[hash.scala 127:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 127:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 127:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 127:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 127:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_key_in; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_key_out; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_sum_in; // @[hash.scala 127:23]
  wire [191:0] pipe1_io_sum_out; // @[hash.scala 127:23]
  wire  pipe2_clock; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[hash.scala 128:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 128:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 128:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 128:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 128:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_key_in; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_key_out; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_sum_in; // @[hash.scala 128:23]
  wire [191:0] pipe2_io_sum_out; // @[hash.scala 128:23]
  wire  pipe3_clock; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[hash.scala 129:23]
  wire [3:0] pipe3_io_pipe_phv_in_next_processor_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 129:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 129:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 129:23]
  wire [3:0] pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 129:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_key_in; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_key_out; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_sum_in; // @[hash.scala 129:23]
  wire [191:0] pipe3_io_sum_out; // @[hash.scala 129:23]
  wire  pipe4_clock; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[hash.scala 130:23]
  wire [3:0] pipe4_io_pipe_phv_in_next_processor_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 130:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 130:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 130:23]
  wire [3:0] pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 130:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_key_in; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_key_out; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_sum_in; // @[hash.scala 130:23]
  wire [191:0] pipe4_io_sum_out; // @[hash.scala 130:23]
  wire  pipe5_clock; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_96; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_97; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_98; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_99; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_100; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_101; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_102; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_103; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_104; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_105; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_106; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_107; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_108; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_109; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_110; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_111; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_112; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_113; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_114; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_115; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_116; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_117; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_118; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_119; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_120; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_121; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_122; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_123; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_124; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_125; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_126; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_127; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_128; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_129; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_130; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_131; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_132; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_133; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_134; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_135; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_136; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_137; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_138; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_139; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_140; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_141; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_142; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_143; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_144; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_145; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_146; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_147; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_148; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_149; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_150; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_151; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_152; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_153; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_154; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_155; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_156; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_157; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_158; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_159; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_pipe_phv_in_next_processor_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_96; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_97; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_98; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_99; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_100; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_101; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_102; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_103; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_104; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_105; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_106; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_107; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_108; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_109; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_110; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_111; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_112; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_113; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_114; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_115; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_116; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_117; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_118; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_119; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_120; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_121; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_122; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_123; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_124; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_125; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_126; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_127; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_128; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_129; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_130; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_131; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_132; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_133; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_134; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_135; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_136; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_137; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_138; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_139; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_140; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_141; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_142; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_143; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_144; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_145; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_146; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_147; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_148; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_149; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_150; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_151; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_152; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_153; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_154; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_155; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_156; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_157; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_158; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_159; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 131:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 131:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_hash_depth_0; // @[hash.scala 131:23]
  wire [3:0] pipe5_io_hash_depth_1; // @[hash.scala 131:23]
  wire [191:0] pipe5_io_key_in; // @[hash.scala 131:23]
  wire [191:0] pipe5_io_key_out; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_sum_in; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_sum_out; // @[hash.scala 131:23]
  wire [15:0] pipe5_io_val_out; // @[hash.scala 131:23]
  wire  pipe6_clock; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_96; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_97; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_98; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_99; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_100; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_101; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_102; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_103; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_104; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_105; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_106; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_107; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_108; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_109; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_110; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_111; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_112; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_113; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_114; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_115; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_116; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_117; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_118; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_119; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_120; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_121; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_122; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_123; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_124; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_125; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_126; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_127; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_128; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_129; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_130; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_131; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_132; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_133; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_134; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_135; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_136; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_137; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_138; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_139; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_140; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_141; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_142; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_143; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_144; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_145; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_146; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_147; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_148; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_149; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_150; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_151; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_152; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_153; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_154; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_155; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_156; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_157; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_158; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_159; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_pipe_phv_in_next_processor_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_96; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_97; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_98; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_99; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_100; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_101; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_102; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_103; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_104; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_105; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_106; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_107; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_108; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_109; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_110; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_111; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_112; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_113; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_114; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_115; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_116; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_117; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_118; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_119; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_120; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_121; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_122; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_123; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_124; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_125; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_126; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_127; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_128; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_129; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_130; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_131; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_132; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_133; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_134; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_135; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_136; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_137; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_138; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_139; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_140; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_141; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_142; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_143; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_144; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_145; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_146; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_147; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_148; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_149; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_150; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_151; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_152; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_153; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_154; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_155; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_156; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_157; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_158; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_159; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 132:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 132:23]
  wire  pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_hash_depth_0; // @[hash.scala 132:23]
  wire [3:0] pipe6_io_hash_depth_1; // @[hash.scala 132:23]
  wire [191:0] pipe6_io_key_in; // @[hash.scala 132:23]
  wire [191:0] pipe6_io_key_out; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_sum_in; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_sum_out; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_val_in; // @[hash.scala 132:23]
  wire [15:0] pipe6_io_val_out; // @[hash.scala 132:23]
  wire  pipe7_clock; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_0; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_1; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_2; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_3; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_4; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_5; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_6; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_7; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_8; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_9; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_10; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_11; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_12; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_13; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_14; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_16; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_17; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_18; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_19; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_20; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_21; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_22; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_23; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_24; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_25; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_26; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_27; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_28; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_29; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_30; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_31; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_32; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_33; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_34; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_35; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_36; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_37; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_38; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_39; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_40; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_41; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_42; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_43; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_44; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_45; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_46; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_47; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_48; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_49; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_50; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_51; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_52; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_53; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_54; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_55; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_56; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_57; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_58; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_59; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_60; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_61; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_62; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_63; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_64; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_65; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_66; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_67; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_68; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_69; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_70; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_71; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_72; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_73; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_74; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_75; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_76; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_77; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_78; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_79; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_80; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_81; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_82; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_83; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_84; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_85; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_86; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_87; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_88; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_89; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_90; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_91; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_92; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_93; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_94; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_95; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_96; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_97; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_98; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_99; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_100; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_101; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_102; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_103; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_104; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_105; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_106; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_107; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_108; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_109; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_110; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_111; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_112; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_113; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_114; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_115; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_116; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_117; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_118; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_119; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_120; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_121; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_122; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_123; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_124; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_125; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_126; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_127; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_128; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_129; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_130; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_131; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_132; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_133; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_134; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_135; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_136; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_137; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_138; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_139; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_140; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_141; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_142; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_143; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_144; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_145; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_146; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_147; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_148; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_149; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_150; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_151; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_152; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_153; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_154; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_155; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_156; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_157; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_158; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_data_159; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_0; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_1; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_2; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_3; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_4; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_5; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_6; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_7; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_8; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_9; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_10; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_11; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_12; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_13; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_14; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_header_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_parse_current_state; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_in_parse_current_offset; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_in_parse_transition_field; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_pipe_phv_in_next_processor_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_in_next_config_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_in_is_valid_processor; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_0; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_1; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_2; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_3; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_4; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_5; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_6; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_7; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_8; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_9; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_10; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_11; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_12; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_13; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_14; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_16; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_17; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_18; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_19; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_20; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_21; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_22; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_23; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_24; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_25; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_26; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_27; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_28; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_29; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_30; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_31; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_32; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_33; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_34; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_35; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_36; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_37; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_38; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_39; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_40; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_41; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_42; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_43; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_44; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_45; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_46; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_47; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_48; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_49; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_50; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_51; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_52; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_53; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_54; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_55; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_56; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_57; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_58; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_59; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_60; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_61; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_62; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_63; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_64; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_65; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_66; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_67; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_68; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_69; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_70; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_71; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_72; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_73; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_74; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_75; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_76; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_77; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_78; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_79; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_80; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_81; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_82; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_83; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_84; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_85; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_86; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_87; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_88; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_89; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_90; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_91; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_92; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_93; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_94; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_95; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_96; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_97; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_98; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_99; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_100; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_101; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_102; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_103; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_104; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_105; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_106; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_107; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_108; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_109; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_110; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_111; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_112; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_113; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_114; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_115; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_116; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_117; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_118; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_119; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_120; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_121; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_122; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_123; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_124; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_125; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_126; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_127; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_128; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_129; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_130; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_131; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_132; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_133; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_134; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_135; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_136; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_137; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_138; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_139; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_140; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_141; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_142; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_143; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_144; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_145; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_146; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_147; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_148; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_149; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_150; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_151; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_152; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_153; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_154; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_155; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_156; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_157; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_158; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_data_159; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_0; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_1; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_2; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_3; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_4; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_5; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_6; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_7; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_8; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_9; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_10; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_11; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_12; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_13; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_14; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_header_15; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_parse_current_state; // @[hash.scala 133:23]
  wire [7:0] pipe7_io_pipe_phv_out_parse_current_offset; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_pipe_phv_out_parse_transition_field; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_pipe_phv_out_next_processor_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_out_next_config_id; // @[hash.scala 133:23]
  wire  pipe7_io_pipe_phv_out_is_valid_processor; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_hash_depth_0; // @[hash.scala 133:23]
  wire [3:0] pipe7_io_hash_depth_1; // @[hash.scala 133:23]
  wire [191:0] pipe7_io_key_in; // @[hash.scala 133:23]
  wire [191:0] pipe7_io_key_out; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_sum_in; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_sum_out; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_val_in; // @[hash.scala 133:23]
  wire [15:0] pipe7_io_val_out; // @[hash.scala 133:23]
  wire  pipe8_clock; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_0; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_1; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_2; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_3; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_4; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_5; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_6; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_7; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_8; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_9; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_10; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_11; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_12; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_13; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_14; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_16; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_17; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_18; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_19; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_20; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_21; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_22; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_23; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_24; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_25; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_26; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_27; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_28; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_29; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_30; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_31; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_32; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_33; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_34; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_35; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_36; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_37; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_38; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_39; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_40; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_41; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_42; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_43; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_44; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_45; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_46; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_47; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_48; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_49; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_50; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_51; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_52; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_53; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_54; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_55; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_56; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_57; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_58; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_59; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_60; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_61; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_62; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_63; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_64; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_65; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_66; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_67; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_68; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_69; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_70; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_71; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_72; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_73; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_74; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_75; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_76; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_77; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_78; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_79; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_80; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_81; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_82; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_83; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_84; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_85; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_86; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_87; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_88; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_89; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_90; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_91; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_92; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_93; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_94; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_95; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_96; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_97; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_98; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_99; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_100; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_101; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_102; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_103; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_104; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_105; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_106; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_107; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_108; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_109; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_110; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_111; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_112; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_113; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_114; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_115; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_116; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_117; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_118; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_119; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_120; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_121; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_122; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_123; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_124; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_125; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_126; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_127; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_128; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_129; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_130; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_131; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_132; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_133; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_134; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_135; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_136; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_137; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_138; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_139; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_140; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_141; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_142; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_143; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_144; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_145; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_146; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_147; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_148; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_149; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_150; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_151; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_152; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_153; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_154; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_155; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_156; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_157; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_158; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_data_159; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_0; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_1; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_2; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_3; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_4; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_5; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_6; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_7; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_8; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_9; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_10; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_11; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_12; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_13; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_14; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_header_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_parse_current_state; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_in_parse_current_offset; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_in_parse_transition_field; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_pipe_phv_in_next_processor_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_in_next_config_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_in_is_valid_processor; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_0; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_1; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_2; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_3; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_4; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_5; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_6; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_7; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_8; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_9; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_10; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_11; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_12; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_13; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_14; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_16; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_17; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_18; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_19; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_20; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_21; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_22; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_23; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_24; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_25; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_26; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_27; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_28; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_29; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_30; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_31; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_32; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_33; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_34; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_35; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_36; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_37; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_38; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_39; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_40; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_41; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_42; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_43; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_44; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_45; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_46; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_47; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_48; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_49; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_50; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_51; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_52; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_53; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_54; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_55; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_56; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_57; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_58; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_59; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_60; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_61; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_62; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_63; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_64; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_65; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_66; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_67; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_68; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_69; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_70; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_71; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_72; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_73; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_74; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_75; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_76; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_77; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_78; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_79; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_80; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_81; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_82; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_83; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_84; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_85; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_86; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_87; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_88; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_89; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_90; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_91; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_92; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_93; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_94; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_95; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_96; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_97; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_98; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_99; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_100; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_101; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_102; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_103; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_104; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_105; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_106; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_107; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_108; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_109; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_110; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_111; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_112; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_113; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_114; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_115; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_116; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_117; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_118; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_119; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_120; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_121; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_122; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_123; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_124; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_125; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_126; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_127; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_128; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_129; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_130; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_131; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_132; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_133; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_134; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_135; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_136; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_137; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_138; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_139; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_140; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_141; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_142; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_143; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_144; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_145; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_146; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_147; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_148; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_149; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_150; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_151; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_152; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_153; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_154; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_155; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_156; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_157; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_158; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_data_159; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_0; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_1; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_2; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_3; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_4; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_5; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_6; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_7; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_8; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_9; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_10; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_11; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_12; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_13; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_14; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_header_15; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_parse_current_state; // @[hash.scala 134:23]
  wire [7:0] pipe8_io_pipe_phv_out_parse_current_offset; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_pipe_phv_out_parse_transition_field; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_pipe_phv_out_next_processor_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_out_next_config_id; // @[hash.scala 134:23]
  wire  pipe8_io_pipe_phv_out_is_valid_processor; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_hash_depth_0; // @[hash.scala 134:23]
  wire [3:0] pipe8_io_hash_depth_1; // @[hash.scala 134:23]
  wire [191:0] pipe8_io_key_in; // @[hash.scala 134:23]
  wire [191:0] pipe8_io_key_out; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_sum_in; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_sum_out; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_val_in; // @[hash.scala 134:23]
  wire [15:0] pipe8_io_val_out; // @[hash.scala 134:23]
  reg [3:0] hash_depth_0; // @[hash.scala 18:26]
  reg [3:0] hash_depth_1; // @[hash.scala 18:26]
  HashSumLevel pipe1 ( // @[hash.scala 127:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe1_io_key_in),
    .io_key_out(pipe1_io_key_out),
    .io_sum_in(pipe1_io_sum_in),
    .io_sum_out(pipe1_io_sum_out)
  );
  HashSumLevel_1 pipe2 ( // @[hash.scala 128:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe2_io_key_in),
    .io_key_out(pipe2_io_key_out),
    .io_sum_in(pipe2_io_sum_in),
    .io_sum_out(pipe2_io_sum_out)
  );
  HashSumLevel_2 pipe3 ( // @[hash.scala 129:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe3_io_key_in),
    .io_key_out(pipe3_io_key_out),
    .io_sum_in(pipe3_io_sum_in),
    .io_sum_out(pipe3_io_sum_out)
  );
  HashSumLevel_3 pipe4 ( // @[hash.scala 130:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_key_in(pipe4_io_key_in),
    .io_key_out(pipe4_io_key_out),
    .io_sum_in(pipe4_io_sum_in),
    .io_sum_out(pipe4_io_sum_out)
  );
  HashReshapeLevel pipe5 ( // @[hash.scala 131:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe5_io_hash_depth_0),
    .io_hash_depth_1(pipe5_io_hash_depth_1),
    .io_key_in(pipe5_io_key_in),
    .io_key_out(pipe5_io_key_out),
    .io_sum_in(pipe5_io_sum_in),
    .io_sum_out(pipe5_io_sum_out),
    .io_val_out(pipe5_io_val_out)
  );
  HashReshapeLevel_1 pipe6 ( // @[hash.scala 132:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe6_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe6_io_hash_depth_0),
    .io_hash_depth_1(pipe6_io_hash_depth_1),
    .io_key_in(pipe6_io_key_in),
    .io_key_out(pipe6_io_key_out),
    .io_sum_in(pipe6_io_sum_in),
    .io_sum_out(pipe6_io_sum_out),
    .io_val_in(pipe6_io_val_in),
    .io_val_out(pipe6_io_val_out)
  );
  HashReshapeLevel_2 pipe7 ( // @[hash.scala 133:23]
    .clock(pipe7_clock),
    .io_pipe_phv_in_data_0(pipe7_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe7_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe7_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe7_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe7_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe7_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe7_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe7_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe7_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe7_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe7_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe7_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe7_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe7_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe7_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe7_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe7_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe7_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe7_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe7_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe7_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe7_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe7_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe7_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe7_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe7_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe7_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe7_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe7_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe7_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe7_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe7_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe7_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe7_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe7_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe7_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe7_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe7_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe7_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe7_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe7_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe7_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe7_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe7_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe7_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe7_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe7_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe7_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe7_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe7_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe7_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe7_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe7_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe7_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe7_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe7_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe7_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe7_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe7_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe7_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe7_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe7_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe7_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe7_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe7_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe7_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe7_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe7_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe7_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe7_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe7_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe7_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe7_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe7_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe7_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe7_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe7_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe7_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe7_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe7_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe7_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe7_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe7_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe7_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe7_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe7_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe7_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe7_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe7_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe7_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe7_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe7_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe7_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe7_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe7_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe7_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe7_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe7_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe7_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe7_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe7_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe7_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe7_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe7_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe7_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe7_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe7_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe7_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe7_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe7_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe7_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe7_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe7_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe7_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe7_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe7_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe7_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe7_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe7_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe7_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe7_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe7_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe7_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe7_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe7_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe7_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe7_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe7_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe7_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe7_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe7_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe7_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe7_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe7_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe7_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe7_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe7_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe7_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe7_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe7_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe7_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe7_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe7_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe7_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe7_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe7_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe7_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe7_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe7_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe7_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe7_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe7_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe7_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe7_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe7_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe7_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe7_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe7_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe7_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe7_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe7_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe7_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe7_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe7_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe7_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe7_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe7_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe7_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe7_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe7_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe7_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe7_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe7_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe7_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe7_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe7_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe7_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe7_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe7_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe7_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe7_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe7_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe7_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe7_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe7_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe7_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe7_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe7_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe7_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe7_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe7_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe7_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe7_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe7_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe7_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe7_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe7_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe7_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe7_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe7_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe7_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe7_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe7_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe7_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe7_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe7_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe7_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe7_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe7_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe7_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe7_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe7_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe7_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe7_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe7_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe7_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe7_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe7_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe7_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe7_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe7_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe7_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe7_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe7_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe7_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe7_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe7_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe7_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe7_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe7_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe7_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe7_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe7_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe7_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe7_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe7_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe7_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe7_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe7_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe7_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe7_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe7_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe7_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe7_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe7_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe7_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe7_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe7_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe7_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe7_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe7_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe7_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe7_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe7_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe7_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe7_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe7_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe7_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe7_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe7_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe7_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe7_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe7_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe7_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe7_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe7_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe7_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe7_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe7_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe7_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe7_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe7_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe7_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe7_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe7_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe7_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe7_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe7_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe7_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe7_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe7_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe7_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe7_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe7_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe7_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe7_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe7_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe7_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe7_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe7_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe7_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe7_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe7_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe7_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe7_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe7_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe7_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe7_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe7_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe7_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe7_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe7_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe7_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe7_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe7_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe7_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe7_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe7_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe7_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe7_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe7_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe7_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe7_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe7_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe7_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe7_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe7_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe7_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe7_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe7_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe7_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe7_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe7_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe7_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe7_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe7_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe7_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe7_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe7_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe7_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe7_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe7_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe7_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe7_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe7_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe7_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe7_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe7_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe7_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe7_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe7_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe7_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe7_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe7_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe7_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe7_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe7_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe7_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe7_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe7_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe7_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe7_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe7_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe7_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe7_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe7_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe7_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe7_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe7_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe7_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe7_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe7_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe7_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe7_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe7_io_hash_depth_0),
    .io_hash_depth_1(pipe7_io_hash_depth_1),
    .io_key_in(pipe7_io_key_in),
    .io_key_out(pipe7_io_key_out),
    .io_sum_in(pipe7_io_sum_in),
    .io_sum_out(pipe7_io_sum_out),
    .io_val_in(pipe7_io_val_in),
    .io_val_out(pipe7_io_val_out)
  );
  HashReshapeLevel_3 pipe8 ( // @[hash.scala 134:23]
    .clock(pipe8_clock),
    .io_pipe_phv_in_data_0(pipe8_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe8_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe8_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe8_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe8_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe8_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe8_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe8_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe8_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe8_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe8_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe8_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe8_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe8_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe8_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe8_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe8_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe8_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe8_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe8_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe8_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe8_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe8_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe8_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe8_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe8_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe8_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe8_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe8_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe8_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe8_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe8_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe8_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe8_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe8_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe8_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe8_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe8_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe8_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe8_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe8_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe8_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe8_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe8_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe8_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe8_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe8_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe8_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe8_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe8_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe8_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe8_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe8_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe8_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe8_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe8_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe8_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe8_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe8_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe8_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe8_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe8_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe8_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe8_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe8_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe8_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe8_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe8_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe8_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe8_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe8_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe8_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe8_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe8_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe8_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe8_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe8_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe8_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe8_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe8_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe8_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe8_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe8_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe8_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe8_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe8_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe8_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe8_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe8_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe8_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe8_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe8_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe8_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe8_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe8_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe8_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe8_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe8_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe8_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe8_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe8_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe8_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe8_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe8_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe8_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe8_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe8_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe8_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe8_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe8_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe8_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe8_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe8_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe8_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe8_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe8_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe8_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe8_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe8_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe8_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe8_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe8_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe8_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe8_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe8_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe8_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe8_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe8_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe8_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe8_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe8_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe8_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe8_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe8_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe8_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe8_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe8_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe8_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe8_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe8_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe8_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe8_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe8_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe8_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe8_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe8_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe8_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe8_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe8_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe8_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe8_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe8_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe8_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe8_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe8_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe8_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe8_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe8_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe8_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe8_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_header_0(pipe8_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe8_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe8_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe8_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe8_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe8_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe8_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe8_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe8_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe8_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe8_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe8_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe8_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe8_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe8_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe8_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe8_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe8_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe8_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe8_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe8_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe8_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe8_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe8_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe8_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe8_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe8_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe8_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe8_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe8_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe8_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe8_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe8_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe8_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe8_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe8_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe8_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe8_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe8_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe8_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe8_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe8_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe8_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe8_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe8_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe8_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe8_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe8_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe8_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe8_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe8_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe8_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe8_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe8_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe8_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe8_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe8_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe8_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe8_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe8_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe8_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe8_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe8_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe8_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe8_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe8_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe8_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe8_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe8_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe8_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe8_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe8_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe8_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe8_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe8_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe8_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe8_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe8_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe8_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe8_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe8_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe8_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe8_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe8_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe8_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe8_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe8_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe8_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe8_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe8_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe8_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe8_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe8_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe8_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe8_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe8_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe8_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe8_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe8_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe8_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe8_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe8_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe8_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe8_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe8_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe8_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe8_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe8_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe8_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe8_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe8_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe8_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe8_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe8_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe8_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe8_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe8_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe8_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe8_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe8_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe8_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe8_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe8_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe8_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe8_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe8_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe8_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe8_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe8_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe8_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe8_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe8_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe8_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe8_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe8_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe8_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe8_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe8_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe8_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe8_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe8_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe8_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe8_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe8_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe8_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe8_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe8_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe8_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe8_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe8_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe8_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe8_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe8_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe8_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe8_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe8_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe8_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe8_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe8_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe8_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe8_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe8_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe8_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe8_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe8_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe8_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe8_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe8_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe8_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe8_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe8_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe8_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe8_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe8_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe8_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe8_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe8_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe8_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe8_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe8_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe8_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe8_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_header_0(pipe8_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe8_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe8_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe8_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe8_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe8_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe8_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe8_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe8_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe8_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe8_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe8_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe8_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe8_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe8_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe8_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe8_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe8_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe8_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe8_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe8_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe8_io_pipe_phv_out_is_valid_processor),
    .io_hash_depth_0(pipe8_io_hash_depth_0),
    .io_hash_depth_1(pipe8_io_hash_depth_1),
    .io_key_in(pipe8_io_key_in),
    .io_key_out(pipe8_io_key_out),
    .io_sum_in(pipe8_io_sum_in),
    .io_sum_out(pipe8_io_sum_out),
    .io_val_in(pipe8_io_val_in),
    .io_val_out(pipe8_io_val_out)
  );
  assign io_pipe_phv_out_data_0 = pipe8_io_pipe_phv_out_data_0; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_1 = pipe8_io_pipe_phv_out_data_1; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_2 = pipe8_io_pipe_phv_out_data_2; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_3 = pipe8_io_pipe_phv_out_data_3; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_4 = pipe8_io_pipe_phv_out_data_4; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_5 = pipe8_io_pipe_phv_out_data_5; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_6 = pipe8_io_pipe_phv_out_data_6; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_7 = pipe8_io_pipe_phv_out_data_7; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_8 = pipe8_io_pipe_phv_out_data_8; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_9 = pipe8_io_pipe_phv_out_data_9; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_10 = pipe8_io_pipe_phv_out_data_10; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_11 = pipe8_io_pipe_phv_out_data_11; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_12 = pipe8_io_pipe_phv_out_data_12; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_13 = pipe8_io_pipe_phv_out_data_13; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_14 = pipe8_io_pipe_phv_out_data_14; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_15 = pipe8_io_pipe_phv_out_data_15; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_16 = pipe8_io_pipe_phv_out_data_16; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_17 = pipe8_io_pipe_phv_out_data_17; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_18 = pipe8_io_pipe_phv_out_data_18; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_19 = pipe8_io_pipe_phv_out_data_19; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_20 = pipe8_io_pipe_phv_out_data_20; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_21 = pipe8_io_pipe_phv_out_data_21; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_22 = pipe8_io_pipe_phv_out_data_22; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_23 = pipe8_io_pipe_phv_out_data_23; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_24 = pipe8_io_pipe_phv_out_data_24; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_25 = pipe8_io_pipe_phv_out_data_25; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_26 = pipe8_io_pipe_phv_out_data_26; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_27 = pipe8_io_pipe_phv_out_data_27; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_28 = pipe8_io_pipe_phv_out_data_28; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_29 = pipe8_io_pipe_phv_out_data_29; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_30 = pipe8_io_pipe_phv_out_data_30; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_31 = pipe8_io_pipe_phv_out_data_31; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_32 = pipe8_io_pipe_phv_out_data_32; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_33 = pipe8_io_pipe_phv_out_data_33; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_34 = pipe8_io_pipe_phv_out_data_34; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_35 = pipe8_io_pipe_phv_out_data_35; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_36 = pipe8_io_pipe_phv_out_data_36; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_37 = pipe8_io_pipe_phv_out_data_37; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_38 = pipe8_io_pipe_phv_out_data_38; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_39 = pipe8_io_pipe_phv_out_data_39; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_40 = pipe8_io_pipe_phv_out_data_40; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_41 = pipe8_io_pipe_phv_out_data_41; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_42 = pipe8_io_pipe_phv_out_data_42; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_43 = pipe8_io_pipe_phv_out_data_43; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_44 = pipe8_io_pipe_phv_out_data_44; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_45 = pipe8_io_pipe_phv_out_data_45; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_46 = pipe8_io_pipe_phv_out_data_46; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_47 = pipe8_io_pipe_phv_out_data_47; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_48 = pipe8_io_pipe_phv_out_data_48; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_49 = pipe8_io_pipe_phv_out_data_49; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_50 = pipe8_io_pipe_phv_out_data_50; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_51 = pipe8_io_pipe_phv_out_data_51; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_52 = pipe8_io_pipe_phv_out_data_52; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_53 = pipe8_io_pipe_phv_out_data_53; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_54 = pipe8_io_pipe_phv_out_data_54; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_55 = pipe8_io_pipe_phv_out_data_55; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_56 = pipe8_io_pipe_phv_out_data_56; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_57 = pipe8_io_pipe_phv_out_data_57; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_58 = pipe8_io_pipe_phv_out_data_58; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_59 = pipe8_io_pipe_phv_out_data_59; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_60 = pipe8_io_pipe_phv_out_data_60; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_61 = pipe8_io_pipe_phv_out_data_61; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_62 = pipe8_io_pipe_phv_out_data_62; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_63 = pipe8_io_pipe_phv_out_data_63; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_64 = pipe8_io_pipe_phv_out_data_64; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_65 = pipe8_io_pipe_phv_out_data_65; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_66 = pipe8_io_pipe_phv_out_data_66; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_67 = pipe8_io_pipe_phv_out_data_67; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_68 = pipe8_io_pipe_phv_out_data_68; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_69 = pipe8_io_pipe_phv_out_data_69; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_70 = pipe8_io_pipe_phv_out_data_70; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_71 = pipe8_io_pipe_phv_out_data_71; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_72 = pipe8_io_pipe_phv_out_data_72; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_73 = pipe8_io_pipe_phv_out_data_73; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_74 = pipe8_io_pipe_phv_out_data_74; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_75 = pipe8_io_pipe_phv_out_data_75; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_76 = pipe8_io_pipe_phv_out_data_76; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_77 = pipe8_io_pipe_phv_out_data_77; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_78 = pipe8_io_pipe_phv_out_data_78; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_79 = pipe8_io_pipe_phv_out_data_79; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_80 = pipe8_io_pipe_phv_out_data_80; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_81 = pipe8_io_pipe_phv_out_data_81; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_82 = pipe8_io_pipe_phv_out_data_82; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_83 = pipe8_io_pipe_phv_out_data_83; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_84 = pipe8_io_pipe_phv_out_data_84; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_85 = pipe8_io_pipe_phv_out_data_85; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_86 = pipe8_io_pipe_phv_out_data_86; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_87 = pipe8_io_pipe_phv_out_data_87; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_88 = pipe8_io_pipe_phv_out_data_88; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_89 = pipe8_io_pipe_phv_out_data_89; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_90 = pipe8_io_pipe_phv_out_data_90; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_91 = pipe8_io_pipe_phv_out_data_91; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_92 = pipe8_io_pipe_phv_out_data_92; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_93 = pipe8_io_pipe_phv_out_data_93; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_94 = pipe8_io_pipe_phv_out_data_94; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_95 = pipe8_io_pipe_phv_out_data_95; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_96 = pipe8_io_pipe_phv_out_data_96; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_97 = pipe8_io_pipe_phv_out_data_97; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_98 = pipe8_io_pipe_phv_out_data_98; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_99 = pipe8_io_pipe_phv_out_data_99; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_100 = pipe8_io_pipe_phv_out_data_100; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_101 = pipe8_io_pipe_phv_out_data_101; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_102 = pipe8_io_pipe_phv_out_data_102; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_103 = pipe8_io_pipe_phv_out_data_103; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_104 = pipe8_io_pipe_phv_out_data_104; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_105 = pipe8_io_pipe_phv_out_data_105; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_106 = pipe8_io_pipe_phv_out_data_106; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_107 = pipe8_io_pipe_phv_out_data_107; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_108 = pipe8_io_pipe_phv_out_data_108; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_109 = pipe8_io_pipe_phv_out_data_109; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_110 = pipe8_io_pipe_phv_out_data_110; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_111 = pipe8_io_pipe_phv_out_data_111; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_112 = pipe8_io_pipe_phv_out_data_112; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_113 = pipe8_io_pipe_phv_out_data_113; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_114 = pipe8_io_pipe_phv_out_data_114; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_115 = pipe8_io_pipe_phv_out_data_115; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_116 = pipe8_io_pipe_phv_out_data_116; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_117 = pipe8_io_pipe_phv_out_data_117; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_118 = pipe8_io_pipe_phv_out_data_118; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_119 = pipe8_io_pipe_phv_out_data_119; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_120 = pipe8_io_pipe_phv_out_data_120; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_121 = pipe8_io_pipe_phv_out_data_121; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_122 = pipe8_io_pipe_phv_out_data_122; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_123 = pipe8_io_pipe_phv_out_data_123; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_124 = pipe8_io_pipe_phv_out_data_124; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_125 = pipe8_io_pipe_phv_out_data_125; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_126 = pipe8_io_pipe_phv_out_data_126; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_127 = pipe8_io_pipe_phv_out_data_127; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_128 = pipe8_io_pipe_phv_out_data_128; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_129 = pipe8_io_pipe_phv_out_data_129; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_130 = pipe8_io_pipe_phv_out_data_130; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_131 = pipe8_io_pipe_phv_out_data_131; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_132 = pipe8_io_pipe_phv_out_data_132; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_133 = pipe8_io_pipe_phv_out_data_133; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_134 = pipe8_io_pipe_phv_out_data_134; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_135 = pipe8_io_pipe_phv_out_data_135; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_136 = pipe8_io_pipe_phv_out_data_136; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_137 = pipe8_io_pipe_phv_out_data_137; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_138 = pipe8_io_pipe_phv_out_data_138; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_139 = pipe8_io_pipe_phv_out_data_139; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_140 = pipe8_io_pipe_phv_out_data_140; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_141 = pipe8_io_pipe_phv_out_data_141; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_142 = pipe8_io_pipe_phv_out_data_142; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_143 = pipe8_io_pipe_phv_out_data_143; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_144 = pipe8_io_pipe_phv_out_data_144; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_145 = pipe8_io_pipe_phv_out_data_145; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_146 = pipe8_io_pipe_phv_out_data_146; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_147 = pipe8_io_pipe_phv_out_data_147; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_148 = pipe8_io_pipe_phv_out_data_148; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_149 = pipe8_io_pipe_phv_out_data_149; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_150 = pipe8_io_pipe_phv_out_data_150; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_151 = pipe8_io_pipe_phv_out_data_151; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_152 = pipe8_io_pipe_phv_out_data_152; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_153 = pipe8_io_pipe_phv_out_data_153; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_154 = pipe8_io_pipe_phv_out_data_154; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_155 = pipe8_io_pipe_phv_out_data_155; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_156 = pipe8_io_pipe_phv_out_data_156; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_157 = pipe8_io_pipe_phv_out_data_157; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_158 = pipe8_io_pipe_phv_out_data_158; // @[hash.scala 176:27]
  assign io_pipe_phv_out_data_159 = pipe8_io_pipe_phv_out_data_159; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_0 = pipe8_io_pipe_phv_out_header_0; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_1 = pipe8_io_pipe_phv_out_header_1; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_2 = pipe8_io_pipe_phv_out_header_2; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_3 = pipe8_io_pipe_phv_out_header_3; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_4 = pipe8_io_pipe_phv_out_header_4; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_5 = pipe8_io_pipe_phv_out_header_5; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_6 = pipe8_io_pipe_phv_out_header_6; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_7 = pipe8_io_pipe_phv_out_header_7; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_8 = pipe8_io_pipe_phv_out_header_8; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_9 = pipe8_io_pipe_phv_out_header_9; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_10 = pipe8_io_pipe_phv_out_header_10; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_11 = pipe8_io_pipe_phv_out_header_11; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_12 = pipe8_io_pipe_phv_out_header_12; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_13 = pipe8_io_pipe_phv_out_header_13; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_14 = pipe8_io_pipe_phv_out_header_14; // @[hash.scala 176:27]
  assign io_pipe_phv_out_header_15 = pipe8_io_pipe_phv_out_header_15; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_current_state = pipe8_io_pipe_phv_out_parse_current_state; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_current_offset = pipe8_io_pipe_phv_out_parse_current_offset; // @[hash.scala 176:27]
  assign io_pipe_phv_out_parse_transition_field = pipe8_io_pipe_phv_out_parse_transition_field; // @[hash.scala 176:27]
  assign io_pipe_phv_out_next_processor_id = pipe8_io_pipe_phv_out_next_processor_id; // @[hash.scala 176:27]
  assign io_pipe_phv_out_next_config_id = pipe8_io_pipe_phv_out_next_config_id; // @[hash.scala 176:27]
  assign io_pipe_phv_out_is_valid_processor = pipe8_io_pipe_phv_out_is_valid_processor; // @[hash.scala 176:27]
  assign io_key_out = pipe8_io_key_out; // @[hash.scala 177:27]
  assign io_hash_val = pipe8_io_sum_out[7:0]; // @[hash.scala 178:46]
  assign io_hash_val_cs = pipe8_io_val_out[15:12]; // @[hash.scala 179:46]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[hash.scala 136:27]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[hash.scala 136:27]
  assign pipe1_io_key_in = io_key_in; // @[hash.scala 137:27]
  assign pipe1_io_sum_in = pipe1_io_key_in; // @[hash.scala 138:27]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[hash.scala 140:27]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[hash.scala 140:27]
  assign pipe2_io_key_in = pipe1_io_key_out; // @[hash.scala 141:27]
  assign pipe2_io_sum_in = pipe1_io_sum_out; // @[hash.scala 142:27]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[hash.scala 144:27]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[hash.scala 144:27]
  assign pipe3_io_key_in = pipe2_io_key_out; // @[hash.scala 145:27]
  assign pipe3_io_sum_in = pipe2_io_sum_out; // @[hash.scala 146:27]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[hash.scala 148:27]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[hash.scala 148:27]
  assign pipe4_io_key_in = pipe3_io_key_out; // @[hash.scala 149:27]
  assign pipe4_io_sum_in = pipe3_io_sum_out; // @[hash.scala 150:27]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_96 = pipe4_io_pipe_phv_out_data_96; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_97 = pipe4_io_pipe_phv_out_data_97; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_98 = pipe4_io_pipe_phv_out_data_98; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_99 = pipe4_io_pipe_phv_out_data_99; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_100 = pipe4_io_pipe_phv_out_data_100; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_101 = pipe4_io_pipe_phv_out_data_101; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_102 = pipe4_io_pipe_phv_out_data_102; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_103 = pipe4_io_pipe_phv_out_data_103; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_104 = pipe4_io_pipe_phv_out_data_104; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_105 = pipe4_io_pipe_phv_out_data_105; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_106 = pipe4_io_pipe_phv_out_data_106; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_107 = pipe4_io_pipe_phv_out_data_107; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_108 = pipe4_io_pipe_phv_out_data_108; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_109 = pipe4_io_pipe_phv_out_data_109; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_110 = pipe4_io_pipe_phv_out_data_110; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_111 = pipe4_io_pipe_phv_out_data_111; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_112 = pipe4_io_pipe_phv_out_data_112; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_113 = pipe4_io_pipe_phv_out_data_113; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_114 = pipe4_io_pipe_phv_out_data_114; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_115 = pipe4_io_pipe_phv_out_data_115; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_116 = pipe4_io_pipe_phv_out_data_116; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_117 = pipe4_io_pipe_phv_out_data_117; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_118 = pipe4_io_pipe_phv_out_data_118; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_119 = pipe4_io_pipe_phv_out_data_119; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_120 = pipe4_io_pipe_phv_out_data_120; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_121 = pipe4_io_pipe_phv_out_data_121; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_122 = pipe4_io_pipe_phv_out_data_122; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_123 = pipe4_io_pipe_phv_out_data_123; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_124 = pipe4_io_pipe_phv_out_data_124; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_125 = pipe4_io_pipe_phv_out_data_125; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_126 = pipe4_io_pipe_phv_out_data_126; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_127 = pipe4_io_pipe_phv_out_data_127; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_128 = pipe4_io_pipe_phv_out_data_128; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_129 = pipe4_io_pipe_phv_out_data_129; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_130 = pipe4_io_pipe_phv_out_data_130; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_131 = pipe4_io_pipe_phv_out_data_131; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_132 = pipe4_io_pipe_phv_out_data_132; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_133 = pipe4_io_pipe_phv_out_data_133; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_134 = pipe4_io_pipe_phv_out_data_134; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_135 = pipe4_io_pipe_phv_out_data_135; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_136 = pipe4_io_pipe_phv_out_data_136; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_137 = pipe4_io_pipe_phv_out_data_137; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_138 = pipe4_io_pipe_phv_out_data_138; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_139 = pipe4_io_pipe_phv_out_data_139; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_140 = pipe4_io_pipe_phv_out_data_140; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_141 = pipe4_io_pipe_phv_out_data_141; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_142 = pipe4_io_pipe_phv_out_data_142; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_143 = pipe4_io_pipe_phv_out_data_143; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_144 = pipe4_io_pipe_phv_out_data_144; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_145 = pipe4_io_pipe_phv_out_data_145; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_146 = pipe4_io_pipe_phv_out_data_146; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_147 = pipe4_io_pipe_phv_out_data_147; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_148 = pipe4_io_pipe_phv_out_data_148; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_149 = pipe4_io_pipe_phv_out_data_149; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_150 = pipe4_io_pipe_phv_out_data_150; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_151 = pipe4_io_pipe_phv_out_data_151; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_152 = pipe4_io_pipe_phv_out_data_152; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_153 = pipe4_io_pipe_phv_out_data_153; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_154 = pipe4_io_pipe_phv_out_data_154; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_155 = pipe4_io_pipe_phv_out_data_155; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_156 = pipe4_io_pipe_phv_out_data_156; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_157 = pipe4_io_pipe_phv_out_data_157; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_158 = pipe4_io_pipe_phv_out_data_158; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_data_159 = pipe4_io_pipe_phv_out_data_159; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[hash.scala 152:27]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[hash.scala 152:27]
  assign pipe5_io_hash_depth_0 = hash_depth_0; // @[hash.scala 156:27]
  assign pipe5_io_hash_depth_1 = hash_depth_1; // @[hash.scala 156:27]
  assign pipe5_io_key_in = pipe4_io_key_out; // @[hash.scala 153:27]
  assign pipe5_io_sum_in = pipe4_io_sum_out[15:0]; // @[hash.scala 154:27]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_96 = pipe5_io_pipe_phv_out_data_96; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_97 = pipe5_io_pipe_phv_out_data_97; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_98 = pipe5_io_pipe_phv_out_data_98; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_99 = pipe5_io_pipe_phv_out_data_99; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_100 = pipe5_io_pipe_phv_out_data_100; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_101 = pipe5_io_pipe_phv_out_data_101; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_102 = pipe5_io_pipe_phv_out_data_102; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_103 = pipe5_io_pipe_phv_out_data_103; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_104 = pipe5_io_pipe_phv_out_data_104; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_105 = pipe5_io_pipe_phv_out_data_105; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_106 = pipe5_io_pipe_phv_out_data_106; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_107 = pipe5_io_pipe_phv_out_data_107; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_108 = pipe5_io_pipe_phv_out_data_108; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_109 = pipe5_io_pipe_phv_out_data_109; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_110 = pipe5_io_pipe_phv_out_data_110; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_111 = pipe5_io_pipe_phv_out_data_111; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_112 = pipe5_io_pipe_phv_out_data_112; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_113 = pipe5_io_pipe_phv_out_data_113; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_114 = pipe5_io_pipe_phv_out_data_114; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_115 = pipe5_io_pipe_phv_out_data_115; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_116 = pipe5_io_pipe_phv_out_data_116; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_117 = pipe5_io_pipe_phv_out_data_117; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_118 = pipe5_io_pipe_phv_out_data_118; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_119 = pipe5_io_pipe_phv_out_data_119; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_120 = pipe5_io_pipe_phv_out_data_120; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_121 = pipe5_io_pipe_phv_out_data_121; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_122 = pipe5_io_pipe_phv_out_data_122; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_123 = pipe5_io_pipe_phv_out_data_123; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_124 = pipe5_io_pipe_phv_out_data_124; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_125 = pipe5_io_pipe_phv_out_data_125; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_126 = pipe5_io_pipe_phv_out_data_126; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_127 = pipe5_io_pipe_phv_out_data_127; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_128 = pipe5_io_pipe_phv_out_data_128; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_129 = pipe5_io_pipe_phv_out_data_129; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_130 = pipe5_io_pipe_phv_out_data_130; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_131 = pipe5_io_pipe_phv_out_data_131; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_132 = pipe5_io_pipe_phv_out_data_132; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_133 = pipe5_io_pipe_phv_out_data_133; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_134 = pipe5_io_pipe_phv_out_data_134; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_135 = pipe5_io_pipe_phv_out_data_135; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_136 = pipe5_io_pipe_phv_out_data_136; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_137 = pipe5_io_pipe_phv_out_data_137; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_138 = pipe5_io_pipe_phv_out_data_138; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_139 = pipe5_io_pipe_phv_out_data_139; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_140 = pipe5_io_pipe_phv_out_data_140; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_141 = pipe5_io_pipe_phv_out_data_141; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_142 = pipe5_io_pipe_phv_out_data_142; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_143 = pipe5_io_pipe_phv_out_data_143; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_144 = pipe5_io_pipe_phv_out_data_144; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_145 = pipe5_io_pipe_phv_out_data_145; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_146 = pipe5_io_pipe_phv_out_data_146; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_147 = pipe5_io_pipe_phv_out_data_147; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_148 = pipe5_io_pipe_phv_out_data_148; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_149 = pipe5_io_pipe_phv_out_data_149; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_150 = pipe5_io_pipe_phv_out_data_150; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_151 = pipe5_io_pipe_phv_out_data_151; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_152 = pipe5_io_pipe_phv_out_data_152; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_153 = pipe5_io_pipe_phv_out_data_153; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_154 = pipe5_io_pipe_phv_out_data_154; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_155 = pipe5_io_pipe_phv_out_data_155; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_156 = pipe5_io_pipe_phv_out_data_156; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_157 = pipe5_io_pipe_phv_out_data_157; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_158 = pipe5_io_pipe_phv_out_data_158; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_data_159 = pipe5_io_pipe_phv_out_data_159; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[hash.scala 158:27]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[hash.scala 158:27]
  assign pipe6_io_hash_depth_0 = hash_depth_0; // @[hash.scala 162:27]
  assign pipe6_io_hash_depth_1 = hash_depth_1; // @[hash.scala 162:27]
  assign pipe6_io_key_in = pipe5_io_key_out; // @[hash.scala 159:27]
  assign pipe6_io_sum_in = pipe5_io_sum_out; // @[hash.scala 160:27]
  assign pipe6_io_val_in = pipe5_io_val_out; // @[hash.scala 161:27]
  assign pipe7_clock = clock;
  assign pipe7_io_pipe_phv_in_data_0 = pipe6_io_pipe_phv_out_data_0; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_1 = pipe6_io_pipe_phv_out_data_1; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_2 = pipe6_io_pipe_phv_out_data_2; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_3 = pipe6_io_pipe_phv_out_data_3; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_4 = pipe6_io_pipe_phv_out_data_4; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_5 = pipe6_io_pipe_phv_out_data_5; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_6 = pipe6_io_pipe_phv_out_data_6; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_7 = pipe6_io_pipe_phv_out_data_7; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_8 = pipe6_io_pipe_phv_out_data_8; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_9 = pipe6_io_pipe_phv_out_data_9; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_10 = pipe6_io_pipe_phv_out_data_10; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_11 = pipe6_io_pipe_phv_out_data_11; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_12 = pipe6_io_pipe_phv_out_data_12; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_13 = pipe6_io_pipe_phv_out_data_13; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_14 = pipe6_io_pipe_phv_out_data_14; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_15 = pipe6_io_pipe_phv_out_data_15; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_16 = pipe6_io_pipe_phv_out_data_16; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_17 = pipe6_io_pipe_phv_out_data_17; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_18 = pipe6_io_pipe_phv_out_data_18; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_19 = pipe6_io_pipe_phv_out_data_19; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_20 = pipe6_io_pipe_phv_out_data_20; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_21 = pipe6_io_pipe_phv_out_data_21; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_22 = pipe6_io_pipe_phv_out_data_22; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_23 = pipe6_io_pipe_phv_out_data_23; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_24 = pipe6_io_pipe_phv_out_data_24; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_25 = pipe6_io_pipe_phv_out_data_25; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_26 = pipe6_io_pipe_phv_out_data_26; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_27 = pipe6_io_pipe_phv_out_data_27; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_28 = pipe6_io_pipe_phv_out_data_28; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_29 = pipe6_io_pipe_phv_out_data_29; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_30 = pipe6_io_pipe_phv_out_data_30; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_31 = pipe6_io_pipe_phv_out_data_31; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_32 = pipe6_io_pipe_phv_out_data_32; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_33 = pipe6_io_pipe_phv_out_data_33; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_34 = pipe6_io_pipe_phv_out_data_34; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_35 = pipe6_io_pipe_phv_out_data_35; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_36 = pipe6_io_pipe_phv_out_data_36; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_37 = pipe6_io_pipe_phv_out_data_37; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_38 = pipe6_io_pipe_phv_out_data_38; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_39 = pipe6_io_pipe_phv_out_data_39; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_40 = pipe6_io_pipe_phv_out_data_40; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_41 = pipe6_io_pipe_phv_out_data_41; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_42 = pipe6_io_pipe_phv_out_data_42; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_43 = pipe6_io_pipe_phv_out_data_43; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_44 = pipe6_io_pipe_phv_out_data_44; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_45 = pipe6_io_pipe_phv_out_data_45; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_46 = pipe6_io_pipe_phv_out_data_46; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_47 = pipe6_io_pipe_phv_out_data_47; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_48 = pipe6_io_pipe_phv_out_data_48; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_49 = pipe6_io_pipe_phv_out_data_49; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_50 = pipe6_io_pipe_phv_out_data_50; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_51 = pipe6_io_pipe_phv_out_data_51; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_52 = pipe6_io_pipe_phv_out_data_52; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_53 = pipe6_io_pipe_phv_out_data_53; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_54 = pipe6_io_pipe_phv_out_data_54; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_55 = pipe6_io_pipe_phv_out_data_55; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_56 = pipe6_io_pipe_phv_out_data_56; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_57 = pipe6_io_pipe_phv_out_data_57; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_58 = pipe6_io_pipe_phv_out_data_58; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_59 = pipe6_io_pipe_phv_out_data_59; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_60 = pipe6_io_pipe_phv_out_data_60; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_61 = pipe6_io_pipe_phv_out_data_61; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_62 = pipe6_io_pipe_phv_out_data_62; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_63 = pipe6_io_pipe_phv_out_data_63; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_64 = pipe6_io_pipe_phv_out_data_64; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_65 = pipe6_io_pipe_phv_out_data_65; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_66 = pipe6_io_pipe_phv_out_data_66; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_67 = pipe6_io_pipe_phv_out_data_67; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_68 = pipe6_io_pipe_phv_out_data_68; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_69 = pipe6_io_pipe_phv_out_data_69; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_70 = pipe6_io_pipe_phv_out_data_70; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_71 = pipe6_io_pipe_phv_out_data_71; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_72 = pipe6_io_pipe_phv_out_data_72; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_73 = pipe6_io_pipe_phv_out_data_73; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_74 = pipe6_io_pipe_phv_out_data_74; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_75 = pipe6_io_pipe_phv_out_data_75; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_76 = pipe6_io_pipe_phv_out_data_76; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_77 = pipe6_io_pipe_phv_out_data_77; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_78 = pipe6_io_pipe_phv_out_data_78; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_79 = pipe6_io_pipe_phv_out_data_79; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_80 = pipe6_io_pipe_phv_out_data_80; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_81 = pipe6_io_pipe_phv_out_data_81; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_82 = pipe6_io_pipe_phv_out_data_82; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_83 = pipe6_io_pipe_phv_out_data_83; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_84 = pipe6_io_pipe_phv_out_data_84; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_85 = pipe6_io_pipe_phv_out_data_85; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_86 = pipe6_io_pipe_phv_out_data_86; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_87 = pipe6_io_pipe_phv_out_data_87; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_88 = pipe6_io_pipe_phv_out_data_88; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_89 = pipe6_io_pipe_phv_out_data_89; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_90 = pipe6_io_pipe_phv_out_data_90; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_91 = pipe6_io_pipe_phv_out_data_91; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_92 = pipe6_io_pipe_phv_out_data_92; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_93 = pipe6_io_pipe_phv_out_data_93; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_94 = pipe6_io_pipe_phv_out_data_94; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_95 = pipe6_io_pipe_phv_out_data_95; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_96 = pipe6_io_pipe_phv_out_data_96; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_97 = pipe6_io_pipe_phv_out_data_97; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_98 = pipe6_io_pipe_phv_out_data_98; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_99 = pipe6_io_pipe_phv_out_data_99; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_100 = pipe6_io_pipe_phv_out_data_100; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_101 = pipe6_io_pipe_phv_out_data_101; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_102 = pipe6_io_pipe_phv_out_data_102; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_103 = pipe6_io_pipe_phv_out_data_103; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_104 = pipe6_io_pipe_phv_out_data_104; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_105 = pipe6_io_pipe_phv_out_data_105; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_106 = pipe6_io_pipe_phv_out_data_106; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_107 = pipe6_io_pipe_phv_out_data_107; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_108 = pipe6_io_pipe_phv_out_data_108; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_109 = pipe6_io_pipe_phv_out_data_109; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_110 = pipe6_io_pipe_phv_out_data_110; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_111 = pipe6_io_pipe_phv_out_data_111; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_112 = pipe6_io_pipe_phv_out_data_112; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_113 = pipe6_io_pipe_phv_out_data_113; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_114 = pipe6_io_pipe_phv_out_data_114; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_115 = pipe6_io_pipe_phv_out_data_115; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_116 = pipe6_io_pipe_phv_out_data_116; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_117 = pipe6_io_pipe_phv_out_data_117; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_118 = pipe6_io_pipe_phv_out_data_118; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_119 = pipe6_io_pipe_phv_out_data_119; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_120 = pipe6_io_pipe_phv_out_data_120; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_121 = pipe6_io_pipe_phv_out_data_121; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_122 = pipe6_io_pipe_phv_out_data_122; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_123 = pipe6_io_pipe_phv_out_data_123; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_124 = pipe6_io_pipe_phv_out_data_124; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_125 = pipe6_io_pipe_phv_out_data_125; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_126 = pipe6_io_pipe_phv_out_data_126; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_127 = pipe6_io_pipe_phv_out_data_127; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_128 = pipe6_io_pipe_phv_out_data_128; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_129 = pipe6_io_pipe_phv_out_data_129; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_130 = pipe6_io_pipe_phv_out_data_130; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_131 = pipe6_io_pipe_phv_out_data_131; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_132 = pipe6_io_pipe_phv_out_data_132; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_133 = pipe6_io_pipe_phv_out_data_133; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_134 = pipe6_io_pipe_phv_out_data_134; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_135 = pipe6_io_pipe_phv_out_data_135; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_136 = pipe6_io_pipe_phv_out_data_136; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_137 = pipe6_io_pipe_phv_out_data_137; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_138 = pipe6_io_pipe_phv_out_data_138; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_139 = pipe6_io_pipe_phv_out_data_139; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_140 = pipe6_io_pipe_phv_out_data_140; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_141 = pipe6_io_pipe_phv_out_data_141; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_142 = pipe6_io_pipe_phv_out_data_142; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_143 = pipe6_io_pipe_phv_out_data_143; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_144 = pipe6_io_pipe_phv_out_data_144; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_145 = pipe6_io_pipe_phv_out_data_145; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_146 = pipe6_io_pipe_phv_out_data_146; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_147 = pipe6_io_pipe_phv_out_data_147; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_148 = pipe6_io_pipe_phv_out_data_148; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_149 = pipe6_io_pipe_phv_out_data_149; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_150 = pipe6_io_pipe_phv_out_data_150; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_151 = pipe6_io_pipe_phv_out_data_151; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_152 = pipe6_io_pipe_phv_out_data_152; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_153 = pipe6_io_pipe_phv_out_data_153; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_154 = pipe6_io_pipe_phv_out_data_154; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_155 = pipe6_io_pipe_phv_out_data_155; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_156 = pipe6_io_pipe_phv_out_data_156; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_157 = pipe6_io_pipe_phv_out_data_157; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_158 = pipe6_io_pipe_phv_out_data_158; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_data_159 = pipe6_io_pipe_phv_out_data_159; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_0 = pipe6_io_pipe_phv_out_header_0; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_1 = pipe6_io_pipe_phv_out_header_1; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_2 = pipe6_io_pipe_phv_out_header_2; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_3 = pipe6_io_pipe_phv_out_header_3; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_4 = pipe6_io_pipe_phv_out_header_4; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_5 = pipe6_io_pipe_phv_out_header_5; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_6 = pipe6_io_pipe_phv_out_header_6; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_7 = pipe6_io_pipe_phv_out_header_7; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_8 = pipe6_io_pipe_phv_out_header_8; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_9 = pipe6_io_pipe_phv_out_header_9; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_10 = pipe6_io_pipe_phv_out_header_10; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_11 = pipe6_io_pipe_phv_out_header_11; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_12 = pipe6_io_pipe_phv_out_header_12; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_13 = pipe6_io_pipe_phv_out_header_13; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_14 = pipe6_io_pipe_phv_out_header_14; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_header_15 = pipe6_io_pipe_phv_out_header_15; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[hash.scala 164:27]
  assign pipe7_io_pipe_phv_in_is_valid_processor = pipe6_io_pipe_phv_out_is_valid_processor; // @[hash.scala 164:27]
  assign pipe7_io_hash_depth_0 = hash_depth_0; // @[hash.scala 168:27]
  assign pipe7_io_hash_depth_1 = hash_depth_1; // @[hash.scala 168:27]
  assign pipe7_io_key_in = pipe6_io_key_out; // @[hash.scala 165:27]
  assign pipe7_io_sum_in = pipe6_io_sum_out; // @[hash.scala 166:27]
  assign pipe7_io_val_in = pipe6_io_val_out; // @[hash.scala 167:27]
  assign pipe8_clock = clock;
  assign pipe8_io_pipe_phv_in_data_0 = pipe7_io_pipe_phv_out_data_0; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_1 = pipe7_io_pipe_phv_out_data_1; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_2 = pipe7_io_pipe_phv_out_data_2; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_3 = pipe7_io_pipe_phv_out_data_3; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_4 = pipe7_io_pipe_phv_out_data_4; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_5 = pipe7_io_pipe_phv_out_data_5; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_6 = pipe7_io_pipe_phv_out_data_6; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_7 = pipe7_io_pipe_phv_out_data_7; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_8 = pipe7_io_pipe_phv_out_data_8; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_9 = pipe7_io_pipe_phv_out_data_9; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_10 = pipe7_io_pipe_phv_out_data_10; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_11 = pipe7_io_pipe_phv_out_data_11; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_12 = pipe7_io_pipe_phv_out_data_12; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_13 = pipe7_io_pipe_phv_out_data_13; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_14 = pipe7_io_pipe_phv_out_data_14; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_15 = pipe7_io_pipe_phv_out_data_15; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_16 = pipe7_io_pipe_phv_out_data_16; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_17 = pipe7_io_pipe_phv_out_data_17; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_18 = pipe7_io_pipe_phv_out_data_18; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_19 = pipe7_io_pipe_phv_out_data_19; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_20 = pipe7_io_pipe_phv_out_data_20; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_21 = pipe7_io_pipe_phv_out_data_21; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_22 = pipe7_io_pipe_phv_out_data_22; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_23 = pipe7_io_pipe_phv_out_data_23; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_24 = pipe7_io_pipe_phv_out_data_24; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_25 = pipe7_io_pipe_phv_out_data_25; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_26 = pipe7_io_pipe_phv_out_data_26; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_27 = pipe7_io_pipe_phv_out_data_27; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_28 = pipe7_io_pipe_phv_out_data_28; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_29 = pipe7_io_pipe_phv_out_data_29; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_30 = pipe7_io_pipe_phv_out_data_30; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_31 = pipe7_io_pipe_phv_out_data_31; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_32 = pipe7_io_pipe_phv_out_data_32; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_33 = pipe7_io_pipe_phv_out_data_33; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_34 = pipe7_io_pipe_phv_out_data_34; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_35 = pipe7_io_pipe_phv_out_data_35; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_36 = pipe7_io_pipe_phv_out_data_36; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_37 = pipe7_io_pipe_phv_out_data_37; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_38 = pipe7_io_pipe_phv_out_data_38; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_39 = pipe7_io_pipe_phv_out_data_39; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_40 = pipe7_io_pipe_phv_out_data_40; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_41 = pipe7_io_pipe_phv_out_data_41; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_42 = pipe7_io_pipe_phv_out_data_42; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_43 = pipe7_io_pipe_phv_out_data_43; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_44 = pipe7_io_pipe_phv_out_data_44; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_45 = pipe7_io_pipe_phv_out_data_45; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_46 = pipe7_io_pipe_phv_out_data_46; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_47 = pipe7_io_pipe_phv_out_data_47; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_48 = pipe7_io_pipe_phv_out_data_48; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_49 = pipe7_io_pipe_phv_out_data_49; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_50 = pipe7_io_pipe_phv_out_data_50; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_51 = pipe7_io_pipe_phv_out_data_51; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_52 = pipe7_io_pipe_phv_out_data_52; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_53 = pipe7_io_pipe_phv_out_data_53; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_54 = pipe7_io_pipe_phv_out_data_54; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_55 = pipe7_io_pipe_phv_out_data_55; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_56 = pipe7_io_pipe_phv_out_data_56; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_57 = pipe7_io_pipe_phv_out_data_57; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_58 = pipe7_io_pipe_phv_out_data_58; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_59 = pipe7_io_pipe_phv_out_data_59; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_60 = pipe7_io_pipe_phv_out_data_60; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_61 = pipe7_io_pipe_phv_out_data_61; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_62 = pipe7_io_pipe_phv_out_data_62; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_63 = pipe7_io_pipe_phv_out_data_63; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_64 = pipe7_io_pipe_phv_out_data_64; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_65 = pipe7_io_pipe_phv_out_data_65; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_66 = pipe7_io_pipe_phv_out_data_66; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_67 = pipe7_io_pipe_phv_out_data_67; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_68 = pipe7_io_pipe_phv_out_data_68; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_69 = pipe7_io_pipe_phv_out_data_69; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_70 = pipe7_io_pipe_phv_out_data_70; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_71 = pipe7_io_pipe_phv_out_data_71; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_72 = pipe7_io_pipe_phv_out_data_72; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_73 = pipe7_io_pipe_phv_out_data_73; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_74 = pipe7_io_pipe_phv_out_data_74; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_75 = pipe7_io_pipe_phv_out_data_75; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_76 = pipe7_io_pipe_phv_out_data_76; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_77 = pipe7_io_pipe_phv_out_data_77; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_78 = pipe7_io_pipe_phv_out_data_78; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_79 = pipe7_io_pipe_phv_out_data_79; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_80 = pipe7_io_pipe_phv_out_data_80; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_81 = pipe7_io_pipe_phv_out_data_81; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_82 = pipe7_io_pipe_phv_out_data_82; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_83 = pipe7_io_pipe_phv_out_data_83; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_84 = pipe7_io_pipe_phv_out_data_84; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_85 = pipe7_io_pipe_phv_out_data_85; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_86 = pipe7_io_pipe_phv_out_data_86; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_87 = pipe7_io_pipe_phv_out_data_87; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_88 = pipe7_io_pipe_phv_out_data_88; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_89 = pipe7_io_pipe_phv_out_data_89; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_90 = pipe7_io_pipe_phv_out_data_90; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_91 = pipe7_io_pipe_phv_out_data_91; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_92 = pipe7_io_pipe_phv_out_data_92; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_93 = pipe7_io_pipe_phv_out_data_93; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_94 = pipe7_io_pipe_phv_out_data_94; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_95 = pipe7_io_pipe_phv_out_data_95; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_96 = pipe7_io_pipe_phv_out_data_96; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_97 = pipe7_io_pipe_phv_out_data_97; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_98 = pipe7_io_pipe_phv_out_data_98; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_99 = pipe7_io_pipe_phv_out_data_99; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_100 = pipe7_io_pipe_phv_out_data_100; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_101 = pipe7_io_pipe_phv_out_data_101; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_102 = pipe7_io_pipe_phv_out_data_102; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_103 = pipe7_io_pipe_phv_out_data_103; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_104 = pipe7_io_pipe_phv_out_data_104; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_105 = pipe7_io_pipe_phv_out_data_105; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_106 = pipe7_io_pipe_phv_out_data_106; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_107 = pipe7_io_pipe_phv_out_data_107; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_108 = pipe7_io_pipe_phv_out_data_108; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_109 = pipe7_io_pipe_phv_out_data_109; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_110 = pipe7_io_pipe_phv_out_data_110; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_111 = pipe7_io_pipe_phv_out_data_111; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_112 = pipe7_io_pipe_phv_out_data_112; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_113 = pipe7_io_pipe_phv_out_data_113; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_114 = pipe7_io_pipe_phv_out_data_114; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_115 = pipe7_io_pipe_phv_out_data_115; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_116 = pipe7_io_pipe_phv_out_data_116; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_117 = pipe7_io_pipe_phv_out_data_117; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_118 = pipe7_io_pipe_phv_out_data_118; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_119 = pipe7_io_pipe_phv_out_data_119; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_120 = pipe7_io_pipe_phv_out_data_120; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_121 = pipe7_io_pipe_phv_out_data_121; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_122 = pipe7_io_pipe_phv_out_data_122; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_123 = pipe7_io_pipe_phv_out_data_123; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_124 = pipe7_io_pipe_phv_out_data_124; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_125 = pipe7_io_pipe_phv_out_data_125; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_126 = pipe7_io_pipe_phv_out_data_126; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_127 = pipe7_io_pipe_phv_out_data_127; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_128 = pipe7_io_pipe_phv_out_data_128; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_129 = pipe7_io_pipe_phv_out_data_129; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_130 = pipe7_io_pipe_phv_out_data_130; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_131 = pipe7_io_pipe_phv_out_data_131; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_132 = pipe7_io_pipe_phv_out_data_132; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_133 = pipe7_io_pipe_phv_out_data_133; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_134 = pipe7_io_pipe_phv_out_data_134; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_135 = pipe7_io_pipe_phv_out_data_135; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_136 = pipe7_io_pipe_phv_out_data_136; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_137 = pipe7_io_pipe_phv_out_data_137; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_138 = pipe7_io_pipe_phv_out_data_138; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_139 = pipe7_io_pipe_phv_out_data_139; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_140 = pipe7_io_pipe_phv_out_data_140; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_141 = pipe7_io_pipe_phv_out_data_141; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_142 = pipe7_io_pipe_phv_out_data_142; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_143 = pipe7_io_pipe_phv_out_data_143; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_144 = pipe7_io_pipe_phv_out_data_144; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_145 = pipe7_io_pipe_phv_out_data_145; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_146 = pipe7_io_pipe_phv_out_data_146; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_147 = pipe7_io_pipe_phv_out_data_147; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_148 = pipe7_io_pipe_phv_out_data_148; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_149 = pipe7_io_pipe_phv_out_data_149; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_150 = pipe7_io_pipe_phv_out_data_150; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_151 = pipe7_io_pipe_phv_out_data_151; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_152 = pipe7_io_pipe_phv_out_data_152; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_153 = pipe7_io_pipe_phv_out_data_153; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_154 = pipe7_io_pipe_phv_out_data_154; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_155 = pipe7_io_pipe_phv_out_data_155; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_156 = pipe7_io_pipe_phv_out_data_156; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_157 = pipe7_io_pipe_phv_out_data_157; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_158 = pipe7_io_pipe_phv_out_data_158; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_data_159 = pipe7_io_pipe_phv_out_data_159; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_0 = pipe7_io_pipe_phv_out_header_0; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_1 = pipe7_io_pipe_phv_out_header_1; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_2 = pipe7_io_pipe_phv_out_header_2; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_3 = pipe7_io_pipe_phv_out_header_3; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_4 = pipe7_io_pipe_phv_out_header_4; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_5 = pipe7_io_pipe_phv_out_header_5; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_6 = pipe7_io_pipe_phv_out_header_6; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_7 = pipe7_io_pipe_phv_out_header_7; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_8 = pipe7_io_pipe_phv_out_header_8; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_9 = pipe7_io_pipe_phv_out_header_9; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_10 = pipe7_io_pipe_phv_out_header_10; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_11 = pipe7_io_pipe_phv_out_header_11; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_12 = pipe7_io_pipe_phv_out_header_12; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_13 = pipe7_io_pipe_phv_out_header_13; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_14 = pipe7_io_pipe_phv_out_header_14; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_header_15 = pipe7_io_pipe_phv_out_header_15; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_current_state = pipe7_io_pipe_phv_out_parse_current_state; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_current_offset = pipe7_io_pipe_phv_out_parse_current_offset; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_parse_transition_field = pipe7_io_pipe_phv_out_parse_transition_field; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_next_processor_id = pipe7_io_pipe_phv_out_next_processor_id; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_next_config_id = pipe7_io_pipe_phv_out_next_config_id; // @[hash.scala 170:27]
  assign pipe8_io_pipe_phv_in_is_valid_processor = pipe7_io_pipe_phv_out_is_valid_processor; // @[hash.scala 170:27]
  assign pipe8_io_hash_depth_0 = hash_depth_0; // @[hash.scala 174:27]
  assign pipe8_io_hash_depth_1 = hash_depth_1; // @[hash.scala 174:27]
  assign pipe8_io_key_in = pipe7_io_key_out; // @[hash.scala 171:27]
  assign pipe8_io_sum_in = pipe7_io_sum_out; // @[hash.scala 172:27]
  assign pipe8_io_val_in = pipe7_io_val_out; // @[hash.scala 173:27]
  always @(posedge clock) begin
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (~io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_0 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
    if (io_mod_hash_depth_mod) begin // @[hash.scala 19:34]
      if (io_mod_config_id) begin // @[hash.scala 20:38]
        hash_depth_1 <= io_mod_hash_depth; // @[hash.scala 20:38]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hash_depth_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  hash_depth_1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
