module Executor(
  input         clock,
  input  [7:0]  io_pipe_phv_in_data_0,
  input  [7:0]  io_pipe_phv_in_data_1,
  input  [7:0]  io_pipe_phv_in_data_2,
  input  [7:0]  io_pipe_phv_in_data_3,
  input  [7:0]  io_pipe_phv_in_data_4,
  input  [7:0]  io_pipe_phv_in_data_5,
  input  [7:0]  io_pipe_phv_in_data_6,
  input  [7:0]  io_pipe_phv_in_data_7,
  input  [7:0]  io_pipe_phv_in_data_8,
  input  [7:0]  io_pipe_phv_in_data_9,
  input  [7:0]  io_pipe_phv_in_data_10,
  input  [7:0]  io_pipe_phv_in_data_11,
  input  [7:0]  io_pipe_phv_in_data_12,
  input  [7:0]  io_pipe_phv_in_data_13,
  input  [7:0]  io_pipe_phv_in_data_14,
  input  [7:0]  io_pipe_phv_in_data_15,
  input  [7:0]  io_pipe_phv_in_data_16,
  input  [7:0]  io_pipe_phv_in_data_17,
  input  [7:0]  io_pipe_phv_in_data_18,
  input  [7:0]  io_pipe_phv_in_data_19,
  input  [7:0]  io_pipe_phv_in_data_20,
  input  [7:0]  io_pipe_phv_in_data_21,
  input  [7:0]  io_pipe_phv_in_data_22,
  input  [7:0]  io_pipe_phv_in_data_23,
  input  [7:0]  io_pipe_phv_in_data_24,
  input  [7:0]  io_pipe_phv_in_data_25,
  input  [7:0]  io_pipe_phv_in_data_26,
  input  [7:0]  io_pipe_phv_in_data_27,
  input  [7:0]  io_pipe_phv_in_data_28,
  input  [7:0]  io_pipe_phv_in_data_29,
  input  [7:0]  io_pipe_phv_in_data_30,
  input  [7:0]  io_pipe_phv_in_data_31,
  input  [7:0]  io_pipe_phv_in_data_32,
  input  [7:0]  io_pipe_phv_in_data_33,
  input  [7:0]  io_pipe_phv_in_data_34,
  input  [7:0]  io_pipe_phv_in_data_35,
  input  [7:0]  io_pipe_phv_in_data_36,
  input  [7:0]  io_pipe_phv_in_data_37,
  input  [7:0]  io_pipe_phv_in_data_38,
  input  [7:0]  io_pipe_phv_in_data_39,
  input  [7:0]  io_pipe_phv_in_data_40,
  input  [7:0]  io_pipe_phv_in_data_41,
  input  [7:0]  io_pipe_phv_in_data_42,
  input  [7:0]  io_pipe_phv_in_data_43,
  input  [7:0]  io_pipe_phv_in_data_44,
  input  [7:0]  io_pipe_phv_in_data_45,
  input  [7:0]  io_pipe_phv_in_data_46,
  input  [7:0]  io_pipe_phv_in_data_47,
  input  [7:0]  io_pipe_phv_in_data_48,
  input  [7:0]  io_pipe_phv_in_data_49,
  input  [7:0]  io_pipe_phv_in_data_50,
  input  [7:0]  io_pipe_phv_in_data_51,
  input  [7:0]  io_pipe_phv_in_data_52,
  input  [7:0]  io_pipe_phv_in_data_53,
  input  [7:0]  io_pipe_phv_in_data_54,
  input  [7:0]  io_pipe_phv_in_data_55,
  input  [7:0]  io_pipe_phv_in_data_56,
  input  [7:0]  io_pipe_phv_in_data_57,
  input  [7:0]  io_pipe_phv_in_data_58,
  input  [7:0]  io_pipe_phv_in_data_59,
  input  [7:0]  io_pipe_phv_in_data_60,
  input  [7:0]  io_pipe_phv_in_data_61,
  input  [7:0]  io_pipe_phv_in_data_62,
  input  [7:0]  io_pipe_phv_in_data_63,
  input  [7:0]  io_pipe_phv_in_data_64,
  input  [7:0]  io_pipe_phv_in_data_65,
  input  [7:0]  io_pipe_phv_in_data_66,
  input  [7:0]  io_pipe_phv_in_data_67,
  input  [7:0]  io_pipe_phv_in_data_68,
  input  [7:0]  io_pipe_phv_in_data_69,
  input  [7:0]  io_pipe_phv_in_data_70,
  input  [7:0]  io_pipe_phv_in_data_71,
  input  [7:0]  io_pipe_phv_in_data_72,
  input  [7:0]  io_pipe_phv_in_data_73,
  input  [7:0]  io_pipe_phv_in_data_74,
  input  [7:0]  io_pipe_phv_in_data_75,
  input  [7:0]  io_pipe_phv_in_data_76,
  input  [7:0]  io_pipe_phv_in_data_77,
  input  [7:0]  io_pipe_phv_in_data_78,
  input  [7:0]  io_pipe_phv_in_data_79,
  input  [7:0]  io_pipe_phv_in_data_80,
  input  [7:0]  io_pipe_phv_in_data_81,
  input  [7:0]  io_pipe_phv_in_data_82,
  input  [7:0]  io_pipe_phv_in_data_83,
  input  [7:0]  io_pipe_phv_in_data_84,
  input  [7:0]  io_pipe_phv_in_data_85,
  input  [7:0]  io_pipe_phv_in_data_86,
  input  [7:0]  io_pipe_phv_in_data_87,
  input  [7:0]  io_pipe_phv_in_data_88,
  input  [7:0]  io_pipe_phv_in_data_89,
  input  [7:0]  io_pipe_phv_in_data_90,
  input  [7:0]  io_pipe_phv_in_data_91,
  input  [7:0]  io_pipe_phv_in_data_92,
  input  [7:0]  io_pipe_phv_in_data_93,
  input  [7:0]  io_pipe_phv_in_data_94,
  input  [7:0]  io_pipe_phv_in_data_95,
  input  [7:0]  io_pipe_phv_in_data_96,
  input  [7:0]  io_pipe_phv_in_data_97,
  input  [7:0]  io_pipe_phv_in_data_98,
  input  [7:0]  io_pipe_phv_in_data_99,
  input  [7:0]  io_pipe_phv_in_data_100,
  input  [7:0]  io_pipe_phv_in_data_101,
  input  [7:0]  io_pipe_phv_in_data_102,
  input  [7:0]  io_pipe_phv_in_data_103,
  input  [7:0]  io_pipe_phv_in_data_104,
  input  [7:0]  io_pipe_phv_in_data_105,
  input  [7:0]  io_pipe_phv_in_data_106,
  input  [7:0]  io_pipe_phv_in_data_107,
  input  [7:0]  io_pipe_phv_in_data_108,
  input  [7:0]  io_pipe_phv_in_data_109,
  input  [7:0]  io_pipe_phv_in_data_110,
  input  [7:0]  io_pipe_phv_in_data_111,
  input  [7:0]  io_pipe_phv_in_data_112,
  input  [7:0]  io_pipe_phv_in_data_113,
  input  [7:0]  io_pipe_phv_in_data_114,
  input  [7:0]  io_pipe_phv_in_data_115,
  input  [7:0]  io_pipe_phv_in_data_116,
  input  [7:0]  io_pipe_phv_in_data_117,
  input  [7:0]  io_pipe_phv_in_data_118,
  input  [7:0]  io_pipe_phv_in_data_119,
  input  [7:0]  io_pipe_phv_in_data_120,
  input  [7:0]  io_pipe_phv_in_data_121,
  input  [7:0]  io_pipe_phv_in_data_122,
  input  [7:0]  io_pipe_phv_in_data_123,
  input  [7:0]  io_pipe_phv_in_data_124,
  input  [7:0]  io_pipe_phv_in_data_125,
  input  [7:0]  io_pipe_phv_in_data_126,
  input  [7:0]  io_pipe_phv_in_data_127,
  input  [7:0]  io_pipe_phv_in_data_128,
  input  [7:0]  io_pipe_phv_in_data_129,
  input  [7:0]  io_pipe_phv_in_data_130,
  input  [7:0]  io_pipe_phv_in_data_131,
  input  [7:0]  io_pipe_phv_in_data_132,
  input  [7:0]  io_pipe_phv_in_data_133,
  input  [7:0]  io_pipe_phv_in_data_134,
  input  [7:0]  io_pipe_phv_in_data_135,
  input  [7:0]  io_pipe_phv_in_data_136,
  input  [7:0]  io_pipe_phv_in_data_137,
  input  [7:0]  io_pipe_phv_in_data_138,
  input  [7:0]  io_pipe_phv_in_data_139,
  input  [7:0]  io_pipe_phv_in_data_140,
  input  [7:0]  io_pipe_phv_in_data_141,
  input  [7:0]  io_pipe_phv_in_data_142,
  input  [7:0]  io_pipe_phv_in_data_143,
  input  [7:0]  io_pipe_phv_in_data_144,
  input  [7:0]  io_pipe_phv_in_data_145,
  input  [7:0]  io_pipe_phv_in_data_146,
  input  [7:0]  io_pipe_phv_in_data_147,
  input  [7:0]  io_pipe_phv_in_data_148,
  input  [7:0]  io_pipe_phv_in_data_149,
  input  [7:0]  io_pipe_phv_in_data_150,
  input  [7:0]  io_pipe_phv_in_data_151,
  input  [7:0]  io_pipe_phv_in_data_152,
  input  [7:0]  io_pipe_phv_in_data_153,
  input  [7:0]  io_pipe_phv_in_data_154,
  input  [7:0]  io_pipe_phv_in_data_155,
  input  [7:0]  io_pipe_phv_in_data_156,
  input  [7:0]  io_pipe_phv_in_data_157,
  input  [7:0]  io_pipe_phv_in_data_158,
  input  [7:0]  io_pipe_phv_in_data_159,
  input  [7:0]  io_pipe_phv_in_data_160,
  input  [7:0]  io_pipe_phv_in_data_161,
  input  [7:0]  io_pipe_phv_in_data_162,
  input  [7:0]  io_pipe_phv_in_data_163,
  input  [7:0]  io_pipe_phv_in_data_164,
  input  [7:0]  io_pipe_phv_in_data_165,
  input  [7:0]  io_pipe_phv_in_data_166,
  input  [7:0]  io_pipe_phv_in_data_167,
  input  [7:0]  io_pipe_phv_in_data_168,
  input  [7:0]  io_pipe_phv_in_data_169,
  input  [7:0]  io_pipe_phv_in_data_170,
  input  [7:0]  io_pipe_phv_in_data_171,
  input  [7:0]  io_pipe_phv_in_data_172,
  input  [7:0]  io_pipe_phv_in_data_173,
  input  [7:0]  io_pipe_phv_in_data_174,
  input  [7:0]  io_pipe_phv_in_data_175,
  input  [7:0]  io_pipe_phv_in_data_176,
  input  [7:0]  io_pipe_phv_in_data_177,
  input  [7:0]  io_pipe_phv_in_data_178,
  input  [7:0]  io_pipe_phv_in_data_179,
  input  [7:0]  io_pipe_phv_in_data_180,
  input  [7:0]  io_pipe_phv_in_data_181,
  input  [7:0]  io_pipe_phv_in_data_182,
  input  [7:0]  io_pipe_phv_in_data_183,
  input  [7:0]  io_pipe_phv_in_data_184,
  input  [7:0]  io_pipe_phv_in_data_185,
  input  [7:0]  io_pipe_phv_in_data_186,
  input  [7:0]  io_pipe_phv_in_data_187,
  input  [7:0]  io_pipe_phv_in_data_188,
  input  [7:0]  io_pipe_phv_in_data_189,
  input  [7:0]  io_pipe_phv_in_data_190,
  input  [7:0]  io_pipe_phv_in_data_191,
  input  [7:0]  io_pipe_phv_in_data_192,
  input  [7:0]  io_pipe_phv_in_data_193,
  input  [7:0]  io_pipe_phv_in_data_194,
  input  [7:0]  io_pipe_phv_in_data_195,
  input  [7:0]  io_pipe_phv_in_data_196,
  input  [7:0]  io_pipe_phv_in_data_197,
  input  [7:0]  io_pipe_phv_in_data_198,
  input  [7:0]  io_pipe_phv_in_data_199,
  input  [7:0]  io_pipe_phv_in_data_200,
  input  [7:0]  io_pipe_phv_in_data_201,
  input  [7:0]  io_pipe_phv_in_data_202,
  input  [7:0]  io_pipe_phv_in_data_203,
  input  [7:0]  io_pipe_phv_in_data_204,
  input  [7:0]  io_pipe_phv_in_data_205,
  input  [7:0]  io_pipe_phv_in_data_206,
  input  [7:0]  io_pipe_phv_in_data_207,
  input  [7:0]  io_pipe_phv_in_data_208,
  input  [7:0]  io_pipe_phv_in_data_209,
  input  [7:0]  io_pipe_phv_in_data_210,
  input  [7:0]  io_pipe_phv_in_data_211,
  input  [7:0]  io_pipe_phv_in_data_212,
  input  [7:0]  io_pipe_phv_in_data_213,
  input  [7:0]  io_pipe_phv_in_data_214,
  input  [7:0]  io_pipe_phv_in_data_215,
  input  [7:0]  io_pipe_phv_in_data_216,
  input  [7:0]  io_pipe_phv_in_data_217,
  input  [7:0]  io_pipe_phv_in_data_218,
  input  [7:0]  io_pipe_phv_in_data_219,
  input  [7:0]  io_pipe_phv_in_data_220,
  input  [7:0]  io_pipe_phv_in_data_221,
  input  [7:0]  io_pipe_phv_in_data_222,
  input  [7:0]  io_pipe_phv_in_data_223,
  input  [7:0]  io_pipe_phv_in_data_224,
  input  [7:0]  io_pipe_phv_in_data_225,
  input  [7:0]  io_pipe_phv_in_data_226,
  input  [7:0]  io_pipe_phv_in_data_227,
  input  [7:0]  io_pipe_phv_in_data_228,
  input  [7:0]  io_pipe_phv_in_data_229,
  input  [7:0]  io_pipe_phv_in_data_230,
  input  [7:0]  io_pipe_phv_in_data_231,
  input  [7:0]  io_pipe_phv_in_data_232,
  input  [7:0]  io_pipe_phv_in_data_233,
  input  [7:0]  io_pipe_phv_in_data_234,
  input  [7:0]  io_pipe_phv_in_data_235,
  input  [7:0]  io_pipe_phv_in_data_236,
  input  [7:0]  io_pipe_phv_in_data_237,
  input  [7:0]  io_pipe_phv_in_data_238,
  input  [7:0]  io_pipe_phv_in_data_239,
  input  [7:0]  io_pipe_phv_in_data_240,
  input  [7:0]  io_pipe_phv_in_data_241,
  input  [7:0]  io_pipe_phv_in_data_242,
  input  [7:0]  io_pipe_phv_in_data_243,
  input  [7:0]  io_pipe_phv_in_data_244,
  input  [7:0]  io_pipe_phv_in_data_245,
  input  [7:0]  io_pipe_phv_in_data_246,
  input  [7:0]  io_pipe_phv_in_data_247,
  input  [7:0]  io_pipe_phv_in_data_248,
  input  [7:0]  io_pipe_phv_in_data_249,
  input  [7:0]  io_pipe_phv_in_data_250,
  input  [7:0]  io_pipe_phv_in_data_251,
  input  [7:0]  io_pipe_phv_in_data_252,
  input  [7:0]  io_pipe_phv_in_data_253,
  input  [7:0]  io_pipe_phv_in_data_254,
  input  [7:0]  io_pipe_phv_in_data_255,
  input  [7:0]  io_pipe_phv_in_data_256,
  input  [7:0]  io_pipe_phv_in_data_257,
  input  [7:0]  io_pipe_phv_in_data_258,
  input  [7:0]  io_pipe_phv_in_data_259,
  input  [7:0]  io_pipe_phv_in_data_260,
  input  [7:0]  io_pipe_phv_in_data_261,
  input  [7:0]  io_pipe_phv_in_data_262,
  input  [7:0]  io_pipe_phv_in_data_263,
  input  [7:0]  io_pipe_phv_in_data_264,
  input  [7:0]  io_pipe_phv_in_data_265,
  input  [7:0]  io_pipe_phv_in_data_266,
  input  [7:0]  io_pipe_phv_in_data_267,
  input  [7:0]  io_pipe_phv_in_data_268,
  input  [7:0]  io_pipe_phv_in_data_269,
  input  [7:0]  io_pipe_phv_in_data_270,
  input  [7:0]  io_pipe_phv_in_data_271,
  input  [7:0]  io_pipe_phv_in_data_272,
  input  [7:0]  io_pipe_phv_in_data_273,
  input  [7:0]  io_pipe_phv_in_data_274,
  input  [7:0]  io_pipe_phv_in_data_275,
  input  [7:0]  io_pipe_phv_in_data_276,
  input  [7:0]  io_pipe_phv_in_data_277,
  input  [7:0]  io_pipe_phv_in_data_278,
  input  [7:0]  io_pipe_phv_in_data_279,
  input  [7:0]  io_pipe_phv_in_data_280,
  input  [7:0]  io_pipe_phv_in_data_281,
  input  [7:0]  io_pipe_phv_in_data_282,
  input  [7:0]  io_pipe_phv_in_data_283,
  input  [7:0]  io_pipe_phv_in_data_284,
  input  [7:0]  io_pipe_phv_in_data_285,
  input  [7:0]  io_pipe_phv_in_data_286,
  input  [7:0]  io_pipe_phv_in_data_287,
  input  [7:0]  io_pipe_phv_in_data_288,
  input  [7:0]  io_pipe_phv_in_data_289,
  input  [7:0]  io_pipe_phv_in_data_290,
  input  [7:0]  io_pipe_phv_in_data_291,
  input  [7:0]  io_pipe_phv_in_data_292,
  input  [7:0]  io_pipe_phv_in_data_293,
  input  [7:0]  io_pipe_phv_in_data_294,
  input  [7:0]  io_pipe_phv_in_data_295,
  input  [7:0]  io_pipe_phv_in_data_296,
  input  [7:0]  io_pipe_phv_in_data_297,
  input  [7:0]  io_pipe_phv_in_data_298,
  input  [7:0]  io_pipe_phv_in_data_299,
  input  [7:0]  io_pipe_phv_in_data_300,
  input  [7:0]  io_pipe_phv_in_data_301,
  input  [7:0]  io_pipe_phv_in_data_302,
  input  [7:0]  io_pipe_phv_in_data_303,
  input  [7:0]  io_pipe_phv_in_data_304,
  input  [7:0]  io_pipe_phv_in_data_305,
  input  [7:0]  io_pipe_phv_in_data_306,
  input  [7:0]  io_pipe_phv_in_data_307,
  input  [7:0]  io_pipe_phv_in_data_308,
  input  [7:0]  io_pipe_phv_in_data_309,
  input  [7:0]  io_pipe_phv_in_data_310,
  input  [7:0]  io_pipe_phv_in_data_311,
  input  [7:0]  io_pipe_phv_in_data_312,
  input  [7:0]  io_pipe_phv_in_data_313,
  input  [7:0]  io_pipe_phv_in_data_314,
  input  [7:0]  io_pipe_phv_in_data_315,
  input  [7:0]  io_pipe_phv_in_data_316,
  input  [7:0]  io_pipe_phv_in_data_317,
  input  [7:0]  io_pipe_phv_in_data_318,
  input  [7:0]  io_pipe_phv_in_data_319,
  input  [7:0]  io_pipe_phv_in_data_320,
  input  [7:0]  io_pipe_phv_in_data_321,
  input  [7:0]  io_pipe_phv_in_data_322,
  input  [7:0]  io_pipe_phv_in_data_323,
  input  [7:0]  io_pipe_phv_in_data_324,
  input  [7:0]  io_pipe_phv_in_data_325,
  input  [7:0]  io_pipe_phv_in_data_326,
  input  [7:0]  io_pipe_phv_in_data_327,
  input  [7:0]  io_pipe_phv_in_data_328,
  input  [7:0]  io_pipe_phv_in_data_329,
  input  [7:0]  io_pipe_phv_in_data_330,
  input  [7:0]  io_pipe_phv_in_data_331,
  input  [7:0]  io_pipe_phv_in_data_332,
  input  [7:0]  io_pipe_phv_in_data_333,
  input  [7:0]  io_pipe_phv_in_data_334,
  input  [7:0]  io_pipe_phv_in_data_335,
  input  [7:0]  io_pipe_phv_in_data_336,
  input  [7:0]  io_pipe_phv_in_data_337,
  input  [7:0]  io_pipe_phv_in_data_338,
  input  [7:0]  io_pipe_phv_in_data_339,
  input  [7:0]  io_pipe_phv_in_data_340,
  input  [7:0]  io_pipe_phv_in_data_341,
  input  [7:0]  io_pipe_phv_in_data_342,
  input  [7:0]  io_pipe_phv_in_data_343,
  input  [7:0]  io_pipe_phv_in_data_344,
  input  [7:0]  io_pipe_phv_in_data_345,
  input  [7:0]  io_pipe_phv_in_data_346,
  input  [7:0]  io_pipe_phv_in_data_347,
  input  [7:0]  io_pipe_phv_in_data_348,
  input  [7:0]  io_pipe_phv_in_data_349,
  input  [7:0]  io_pipe_phv_in_data_350,
  input  [7:0]  io_pipe_phv_in_data_351,
  input  [7:0]  io_pipe_phv_in_data_352,
  input  [7:0]  io_pipe_phv_in_data_353,
  input  [7:0]  io_pipe_phv_in_data_354,
  input  [7:0]  io_pipe_phv_in_data_355,
  input  [7:0]  io_pipe_phv_in_data_356,
  input  [7:0]  io_pipe_phv_in_data_357,
  input  [7:0]  io_pipe_phv_in_data_358,
  input  [7:0]  io_pipe_phv_in_data_359,
  input  [7:0]  io_pipe_phv_in_data_360,
  input  [7:0]  io_pipe_phv_in_data_361,
  input  [7:0]  io_pipe_phv_in_data_362,
  input  [7:0]  io_pipe_phv_in_data_363,
  input  [7:0]  io_pipe_phv_in_data_364,
  input  [7:0]  io_pipe_phv_in_data_365,
  input  [7:0]  io_pipe_phv_in_data_366,
  input  [7:0]  io_pipe_phv_in_data_367,
  input  [7:0]  io_pipe_phv_in_data_368,
  input  [7:0]  io_pipe_phv_in_data_369,
  input  [7:0]  io_pipe_phv_in_data_370,
  input  [7:0]  io_pipe_phv_in_data_371,
  input  [7:0]  io_pipe_phv_in_data_372,
  input  [7:0]  io_pipe_phv_in_data_373,
  input  [7:0]  io_pipe_phv_in_data_374,
  input  [7:0]  io_pipe_phv_in_data_375,
  input  [7:0]  io_pipe_phv_in_data_376,
  input  [7:0]  io_pipe_phv_in_data_377,
  input  [7:0]  io_pipe_phv_in_data_378,
  input  [7:0]  io_pipe_phv_in_data_379,
  input  [7:0]  io_pipe_phv_in_data_380,
  input  [7:0]  io_pipe_phv_in_data_381,
  input  [7:0]  io_pipe_phv_in_data_382,
  input  [7:0]  io_pipe_phv_in_data_383,
  input  [7:0]  io_pipe_phv_in_data_384,
  input  [7:0]  io_pipe_phv_in_data_385,
  input  [7:0]  io_pipe_phv_in_data_386,
  input  [7:0]  io_pipe_phv_in_data_387,
  input  [7:0]  io_pipe_phv_in_data_388,
  input  [7:0]  io_pipe_phv_in_data_389,
  input  [7:0]  io_pipe_phv_in_data_390,
  input  [7:0]  io_pipe_phv_in_data_391,
  input  [7:0]  io_pipe_phv_in_data_392,
  input  [7:0]  io_pipe_phv_in_data_393,
  input  [7:0]  io_pipe_phv_in_data_394,
  input  [7:0]  io_pipe_phv_in_data_395,
  input  [7:0]  io_pipe_phv_in_data_396,
  input  [7:0]  io_pipe_phv_in_data_397,
  input  [7:0]  io_pipe_phv_in_data_398,
  input  [7:0]  io_pipe_phv_in_data_399,
  input  [7:0]  io_pipe_phv_in_data_400,
  input  [7:0]  io_pipe_phv_in_data_401,
  input  [7:0]  io_pipe_phv_in_data_402,
  input  [7:0]  io_pipe_phv_in_data_403,
  input  [7:0]  io_pipe_phv_in_data_404,
  input  [7:0]  io_pipe_phv_in_data_405,
  input  [7:0]  io_pipe_phv_in_data_406,
  input  [7:0]  io_pipe_phv_in_data_407,
  input  [7:0]  io_pipe_phv_in_data_408,
  input  [7:0]  io_pipe_phv_in_data_409,
  input  [7:0]  io_pipe_phv_in_data_410,
  input  [7:0]  io_pipe_phv_in_data_411,
  input  [7:0]  io_pipe_phv_in_data_412,
  input  [7:0]  io_pipe_phv_in_data_413,
  input  [7:0]  io_pipe_phv_in_data_414,
  input  [7:0]  io_pipe_phv_in_data_415,
  input  [7:0]  io_pipe_phv_in_data_416,
  input  [7:0]  io_pipe_phv_in_data_417,
  input  [7:0]  io_pipe_phv_in_data_418,
  input  [7:0]  io_pipe_phv_in_data_419,
  input  [7:0]  io_pipe_phv_in_data_420,
  input  [7:0]  io_pipe_phv_in_data_421,
  input  [7:0]  io_pipe_phv_in_data_422,
  input  [7:0]  io_pipe_phv_in_data_423,
  input  [7:0]  io_pipe_phv_in_data_424,
  input  [7:0]  io_pipe_phv_in_data_425,
  input  [7:0]  io_pipe_phv_in_data_426,
  input  [7:0]  io_pipe_phv_in_data_427,
  input  [7:0]  io_pipe_phv_in_data_428,
  input  [7:0]  io_pipe_phv_in_data_429,
  input  [7:0]  io_pipe_phv_in_data_430,
  input  [7:0]  io_pipe_phv_in_data_431,
  input  [7:0]  io_pipe_phv_in_data_432,
  input  [7:0]  io_pipe_phv_in_data_433,
  input  [7:0]  io_pipe_phv_in_data_434,
  input  [7:0]  io_pipe_phv_in_data_435,
  input  [7:0]  io_pipe_phv_in_data_436,
  input  [7:0]  io_pipe_phv_in_data_437,
  input  [7:0]  io_pipe_phv_in_data_438,
  input  [7:0]  io_pipe_phv_in_data_439,
  input  [7:0]  io_pipe_phv_in_data_440,
  input  [7:0]  io_pipe_phv_in_data_441,
  input  [7:0]  io_pipe_phv_in_data_442,
  input  [7:0]  io_pipe_phv_in_data_443,
  input  [7:0]  io_pipe_phv_in_data_444,
  input  [7:0]  io_pipe_phv_in_data_445,
  input  [7:0]  io_pipe_phv_in_data_446,
  input  [7:0]  io_pipe_phv_in_data_447,
  input  [7:0]  io_pipe_phv_in_data_448,
  input  [7:0]  io_pipe_phv_in_data_449,
  input  [7:0]  io_pipe_phv_in_data_450,
  input  [7:0]  io_pipe_phv_in_data_451,
  input  [7:0]  io_pipe_phv_in_data_452,
  input  [7:0]  io_pipe_phv_in_data_453,
  input  [7:0]  io_pipe_phv_in_data_454,
  input  [7:0]  io_pipe_phv_in_data_455,
  input  [7:0]  io_pipe_phv_in_data_456,
  input  [7:0]  io_pipe_phv_in_data_457,
  input  [7:0]  io_pipe_phv_in_data_458,
  input  [7:0]  io_pipe_phv_in_data_459,
  input  [7:0]  io_pipe_phv_in_data_460,
  input  [7:0]  io_pipe_phv_in_data_461,
  input  [7:0]  io_pipe_phv_in_data_462,
  input  [7:0]  io_pipe_phv_in_data_463,
  input  [7:0]  io_pipe_phv_in_data_464,
  input  [7:0]  io_pipe_phv_in_data_465,
  input  [7:0]  io_pipe_phv_in_data_466,
  input  [7:0]  io_pipe_phv_in_data_467,
  input  [7:0]  io_pipe_phv_in_data_468,
  input  [7:0]  io_pipe_phv_in_data_469,
  input  [7:0]  io_pipe_phv_in_data_470,
  input  [7:0]  io_pipe_phv_in_data_471,
  input  [7:0]  io_pipe_phv_in_data_472,
  input  [7:0]  io_pipe_phv_in_data_473,
  input  [7:0]  io_pipe_phv_in_data_474,
  input  [7:0]  io_pipe_phv_in_data_475,
  input  [7:0]  io_pipe_phv_in_data_476,
  input  [7:0]  io_pipe_phv_in_data_477,
  input  [7:0]  io_pipe_phv_in_data_478,
  input  [7:0]  io_pipe_phv_in_data_479,
  input  [7:0]  io_pipe_phv_in_data_480,
  input  [7:0]  io_pipe_phv_in_data_481,
  input  [7:0]  io_pipe_phv_in_data_482,
  input  [7:0]  io_pipe_phv_in_data_483,
  input  [7:0]  io_pipe_phv_in_data_484,
  input  [7:0]  io_pipe_phv_in_data_485,
  input  [7:0]  io_pipe_phv_in_data_486,
  input  [7:0]  io_pipe_phv_in_data_487,
  input  [7:0]  io_pipe_phv_in_data_488,
  input  [7:0]  io_pipe_phv_in_data_489,
  input  [7:0]  io_pipe_phv_in_data_490,
  input  [7:0]  io_pipe_phv_in_data_491,
  input  [7:0]  io_pipe_phv_in_data_492,
  input  [7:0]  io_pipe_phv_in_data_493,
  input  [7:0]  io_pipe_phv_in_data_494,
  input  [7:0]  io_pipe_phv_in_data_495,
  input  [7:0]  io_pipe_phv_in_data_496,
  input  [7:0]  io_pipe_phv_in_data_497,
  input  [7:0]  io_pipe_phv_in_data_498,
  input  [7:0]  io_pipe_phv_in_data_499,
  input  [7:0]  io_pipe_phv_in_data_500,
  input  [7:0]  io_pipe_phv_in_data_501,
  input  [7:0]  io_pipe_phv_in_data_502,
  input  [7:0]  io_pipe_phv_in_data_503,
  input  [7:0]  io_pipe_phv_in_data_504,
  input  [7:0]  io_pipe_phv_in_data_505,
  input  [7:0]  io_pipe_phv_in_data_506,
  input  [7:0]  io_pipe_phv_in_data_507,
  input  [7:0]  io_pipe_phv_in_data_508,
  input  [7:0]  io_pipe_phv_in_data_509,
  input  [7:0]  io_pipe_phv_in_data_510,
  input  [7:0]  io_pipe_phv_in_data_511,
  input  [15:0] io_pipe_phv_in_header_0,
  input  [15:0] io_pipe_phv_in_header_1,
  input  [15:0] io_pipe_phv_in_header_2,
  input  [15:0] io_pipe_phv_in_header_3,
  input  [15:0] io_pipe_phv_in_header_4,
  input  [15:0] io_pipe_phv_in_header_5,
  input  [15:0] io_pipe_phv_in_header_6,
  input  [15:0] io_pipe_phv_in_header_7,
  input  [15:0] io_pipe_phv_in_header_8,
  input  [15:0] io_pipe_phv_in_header_9,
  input  [15:0] io_pipe_phv_in_header_10,
  input  [15:0] io_pipe_phv_in_header_11,
  input  [15:0] io_pipe_phv_in_header_12,
  input  [15:0] io_pipe_phv_in_header_13,
  input  [15:0] io_pipe_phv_in_header_14,
  input  [15:0] io_pipe_phv_in_header_15,
  input  [7:0]  io_pipe_phv_in_parse_current_state,
  input  [7:0]  io_pipe_phv_in_parse_current_offset,
  input  [15:0] io_pipe_phv_in_parse_transition_field,
  input  [3:0]  io_pipe_phv_in_next_processor_id,
  input         io_pipe_phv_in_next_config_id,
  input         io_pipe_phv_in_is_valid_processor,
  output [7:0]  io_pipe_phv_out_data_0,
  output [7:0]  io_pipe_phv_out_data_1,
  output [7:0]  io_pipe_phv_out_data_2,
  output [7:0]  io_pipe_phv_out_data_3,
  output [7:0]  io_pipe_phv_out_data_4,
  output [7:0]  io_pipe_phv_out_data_5,
  output [7:0]  io_pipe_phv_out_data_6,
  output [7:0]  io_pipe_phv_out_data_7,
  output [7:0]  io_pipe_phv_out_data_8,
  output [7:0]  io_pipe_phv_out_data_9,
  output [7:0]  io_pipe_phv_out_data_10,
  output [7:0]  io_pipe_phv_out_data_11,
  output [7:0]  io_pipe_phv_out_data_12,
  output [7:0]  io_pipe_phv_out_data_13,
  output [7:0]  io_pipe_phv_out_data_14,
  output [7:0]  io_pipe_phv_out_data_15,
  output [7:0]  io_pipe_phv_out_data_16,
  output [7:0]  io_pipe_phv_out_data_17,
  output [7:0]  io_pipe_phv_out_data_18,
  output [7:0]  io_pipe_phv_out_data_19,
  output [7:0]  io_pipe_phv_out_data_20,
  output [7:0]  io_pipe_phv_out_data_21,
  output [7:0]  io_pipe_phv_out_data_22,
  output [7:0]  io_pipe_phv_out_data_23,
  output [7:0]  io_pipe_phv_out_data_24,
  output [7:0]  io_pipe_phv_out_data_25,
  output [7:0]  io_pipe_phv_out_data_26,
  output [7:0]  io_pipe_phv_out_data_27,
  output [7:0]  io_pipe_phv_out_data_28,
  output [7:0]  io_pipe_phv_out_data_29,
  output [7:0]  io_pipe_phv_out_data_30,
  output [7:0]  io_pipe_phv_out_data_31,
  output [7:0]  io_pipe_phv_out_data_32,
  output [7:0]  io_pipe_phv_out_data_33,
  output [7:0]  io_pipe_phv_out_data_34,
  output [7:0]  io_pipe_phv_out_data_35,
  output [7:0]  io_pipe_phv_out_data_36,
  output [7:0]  io_pipe_phv_out_data_37,
  output [7:0]  io_pipe_phv_out_data_38,
  output [7:0]  io_pipe_phv_out_data_39,
  output [7:0]  io_pipe_phv_out_data_40,
  output [7:0]  io_pipe_phv_out_data_41,
  output [7:0]  io_pipe_phv_out_data_42,
  output [7:0]  io_pipe_phv_out_data_43,
  output [7:0]  io_pipe_phv_out_data_44,
  output [7:0]  io_pipe_phv_out_data_45,
  output [7:0]  io_pipe_phv_out_data_46,
  output [7:0]  io_pipe_phv_out_data_47,
  output [7:0]  io_pipe_phv_out_data_48,
  output [7:0]  io_pipe_phv_out_data_49,
  output [7:0]  io_pipe_phv_out_data_50,
  output [7:0]  io_pipe_phv_out_data_51,
  output [7:0]  io_pipe_phv_out_data_52,
  output [7:0]  io_pipe_phv_out_data_53,
  output [7:0]  io_pipe_phv_out_data_54,
  output [7:0]  io_pipe_phv_out_data_55,
  output [7:0]  io_pipe_phv_out_data_56,
  output [7:0]  io_pipe_phv_out_data_57,
  output [7:0]  io_pipe_phv_out_data_58,
  output [7:0]  io_pipe_phv_out_data_59,
  output [7:0]  io_pipe_phv_out_data_60,
  output [7:0]  io_pipe_phv_out_data_61,
  output [7:0]  io_pipe_phv_out_data_62,
  output [7:0]  io_pipe_phv_out_data_63,
  output [7:0]  io_pipe_phv_out_data_64,
  output [7:0]  io_pipe_phv_out_data_65,
  output [7:0]  io_pipe_phv_out_data_66,
  output [7:0]  io_pipe_phv_out_data_67,
  output [7:0]  io_pipe_phv_out_data_68,
  output [7:0]  io_pipe_phv_out_data_69,
  output [7:0]  io_pipe_phv_out_data_70,
  output [7:0]  io_pipe_phv_out_data_71,
  output [7:0]  io_pipe_phv_out_data_72,
  output [7:0]  io_pipe_phv_out_data_73,
  output [7:0]  io_pipe_phv_out_data_74,
  output [7:0]  io_pipe_phv_out_data_75,
  output [7:0]  io_pipe_phv_out_data_76,
  output [7:0]  io_pipe_phv_out_data_77,
  output [7:0]  io_pipe_phv_out_data_78,
  output [7:0]  io_pipe_phv_out_data_79,
  output [7:0]  io_pipe_phv_out_data_80,
  output [7:0]  io_pipe_phv_out_data_81,
  output [7:0]  io_pipe_phv_out_data_82,
  output [7:0]  io_pipe_phv_out_data_83,
  output [7:0]  io_pipe_phv_out_data_84,
  output [7:0]  io_pipe_phv_out_data_85,
  output [7:0]  io_pipe_phv_out_data_86,
  output [7:0]  io_pipe_phv_out_data_87,
  output [7:0]  io_pipe_phv_out_data_88,
  output [7:0]  io_pipe_phv_out_data_89,
  output [7:0]  io_pipe_phv_out_data_90,
  output [7:0]  io_pipe_phv_out_data_91,
  output [7:0]  io_pipe_phv_out_data_92,
  output [7:0]  io_pipe_phv_out_data_93,
  output [7:0]  io_pipe_phv_out_data_94,
  output [7:0]  io_pipe_phv_out_data_95,
  output [7:0]  io_pipe_phv_out_data_96,
  output [7:0]  io_pipe_phv_out_data_97,
  output [7:0]  io_pipe_phv_out_data_98,
  output [7:0]  io_pipe_phv_out_data_99,
  output [7:0]  io_pipe_phv_out_data_100,
  output [7:0]  io_pipe_phv_out_data_101,
  output [7:0]  io_pipe_phv_out_data_102,
  output [7:0]  io_pipe_phv_out_data_103,
  output [7:0]  io_pipe_phv_out_data_104,
  output [7:0]  io_pipe_phv_out_data_105,
  output [7:0]  io_pipe_phv_out_data_106,
  output [7:0]  io_pipe_phv_out_data_107,
  output [7:0]  io_pipe_phv_out_data_108,
  output [7:0]  io_pipe_phv_out_data_109,
  output [7:0]  io_pipe_phv_out_data_110,
  output [7:0]  io_pipe_phv_out_data_111,
  output [7:0]  io_pipe_phv_out_data_112,
  output [7:0]  io_pipe_phv_out_data_113,
  output [7:0]  io_pipe_phv_out_data_114,
  output [7:0]  io_pipe_phv_out_data_115,
  output [7:0]  io_pipe_phv_out_data_116,
  output [7:0]  io_pipe_phv_out_data_117,
  output [7:0]  io_pipe_phv_out_data_118,
  output [7:0]  io_pipe_phv_out_data_119,
  output [7:0]  io_pipe_phv_out_data_120,
  output [7:0]  io_pipe_phv_out_data_121,
  output [7:0]  io_pipe_phv_out_data_122,
  output [7:0]  io_pipe_phv_out_data_123,
  output [7:0]  io_pipe_phv_out_data_124,
  output [7:0]  io_pipe_phv_out_data_125,
  output [7:0]  io_pipe_phv_out_data_126,
  output [7:0]  io_pipe_phv_out_data_127,
  output [7:0]  io_pipe_phv_out_data_128,
  output [7:0]  io_pipe_phv_out_data_129,
  output [7:0]  io_pipe_phv_out_data_130,
  output [7:0]  io_pipe_phv_out_data_131,
  output [7:0]  io_pipe_phv_out_data_132,
  output [7:0]  io_pipe_phv_out_data_133,
  output [7:0]  io_pipe_phv_out_data_134,
  output [7:0]  io_pipe_phv_out_data_135,
  output [7:0]  io_pipe_phv_out_data_136,
  output [7:0]  io_pipe_phv_out_data_137,
  output [7:0]  io_pipe_phv_out_data_138,
  output [7:0]  io_pipe_phv_out_data_139,
  output [7:0]  io_pipe_phv_out_data_140,
  output [7:0]  io_pipe_phv_out_data_141,
  output [7:0]  io_pipe_phv_out_data_142,
  output [7:0]  io_pipe_phv_out_data_143,
  output [7:0]  io_pipe_phv_out_data_144,
  output [7:0]  io_pipe_phv_out_data_145,
  output [7:0]  io_pipe_phv_out_data_146,
  output [7:0]  io_pipe_phv_out_data_147,
  output [7:0]  io_pipe_phv_out_data_148,
  output [7:0]  io_pipe_phv_out_data_149,
  output [7:0]  io_pipe_phv_out_data_150,
  output [7:0]  io_pipe_phv_out_data_151,
  output [7:0]  io_pipe_phv_out_data_152,
  output [7:0]  io_pipe_phv_out_data_153,
  output [7:0]  io_pipe_phv_out_data_154,
  output [7:0]  io_pipe_phv_out_data_155,
  output [7:0]  io_pipe_phv_out_data_156,
  output [7:0]  io_pipe_phv_out_data_157,
  output [7:0]  io_pipe_phv_out_data_158,
  output [7:0]  io_pipe_phv_out_data_159,
  output [7:0]  io_pipe_phv_out_data_160,
  output [7:0]  io_pipe_phv_out_data_161,
  output [7:0]  io_pipe_phv_out_data_162,
  output [7:0]  io_pipe_phv_out_data_163,
  output [7:0]  io_pipe_phv_out_data_164,
  output [7:0]  io_pipe_phv_out_data_165,
  output [7:0]  io_pipe_phv_out_data_166,
  output [7:0]  io_pipe_phv_out_data_167,
  output [7:0]  io_pipe_phv_out_data_168,
  output [7:0]  io_pipe_phv_out_data_169,
  output [7:0]  io_pipe_phv_out_data_170,
  output [7:0]  io_pipe_phv_out_data_171,
  output [7:0]  io_pipe_phv_out_data_172,
  output [7:0]  io_pipe_phv_out_data_173,
  output [7:0]  io_pipe_phv_out_data_174,
  output [7:0]  io_pipe_phv_out_data_175,
  output [7:0]  io_pipe_phv_out_data_176,
  output [7:0]  io_pipe_phv_out_data_177,
  output [7:0]  io_pipe_phv_out_data_178,
  output [7:0]  io_pipe_phv_out_data_179,
  output [7:0]  io_pipe_phv_out_data_180,
  output [7:0]  io_pipe_phv_out_data_181,
  output [7:0]  io_pipe_phv_out_data_182,
  output [7:0]  io_pipe_phv_out_data_183,
  output [7:0]  io_pipe_phv_out_data_184,
  output [7:0]  io_pipe_phv_out_data_185,
  output [7:0]  io_pipe_phv_out_data_186,
  output [7:0]  io_pipe_phv_out_data_187,
  output [7:0]  io_pipe_phv_out_data_188,
  output [7:0]  io_pipe_phv_out_data_189,
  output [7:0]  io_pipe_phv_out_data_190,
  output [7:0]  io_pipe_phv_out_data_191,
  output [7:0]  io_pipe_phv_out_data_192,
  output [7:0]  io_pipe_phv_out_data_193,
  output [7:0]  io_pipe_phv_out_data_194,
  output [7:0]  io_pipe_phv_out_data_195,
  output [7:0]  io_pipe_phv_out_data_196,
  output [7:0]  io_pipe_phv_out_data_197,
  output [7:0]  io_pipe_phv_out_data_198,
  output [7:0]  io_pipe_phv_out_data_199,
  output [7:0]  io_pipe_phv_out_data_200,
  output [7:0]  io_pipe_phv_out_data_201,
  output [7:0]  io_pipe_phv_out_data_202,
  output [7:0]  io_pipe_phv_out_data_203,
  output [7:0]  io_pipe_phv_out_data_204,
  output [7:0]  io_pipe_phv_out_data_205,
  output [7:0]  io_pipe_phv_out_data_206,
  output [7:0]  io_pipe_phv_out_data_207,
  output [7:0]  io_pipe_phv_out_data_208,
  output [7:0]  io_pipe_phv_out_data_209,
  output [7:0]  io_pipe_phv_out_data_210,
  output [7:0]  io_pipe_phv_out_data_211,
  output [7:0]  io_pipe_phv_out_data_212,
  output [7:0]  io_pipe_phv_out_data_213,
  output [7:0]  io_pipe_phv_out_data_214,
  output [7:0]  io_pipe_phv_out_data_215,
  output [7:0]  io_pipe_phv_out_data_216,
  output [7:0]  io_pipe_phv_out_data_217,
  output [7:0]  io_pipe_phv_out_data_218,
  output [7:0]  io_pipe_phv_out_data_219,
  output [7:0]  io_pipe_phv_out_data_220,
  output [7:0]  io_pipe_phv_out_data_221,
  output [7:0]  io_pipe_phv_out_data_222,
  output [7:0]  io_pipe_phv_out_data_223,
  output [7:0]  io_pipe_phv_out_data_224,
  output [7:0]  io_pipe_phv_out_data_225,
  output [7:0]  io_pipe_phv_out_data_226,
  output [7:0]  io_pipe_phv_out_data_227,
  output [7:0]  io_pipe_phv_out_data_228,
  output [7:0]  io_pipe_phv_out_data_229,
  output [7:0]  io_pipe_phv_out_data_230,
  output [7:0]  io_pipe_phv_out_data_231,
  output [7:0]  io_pipe_phv_out_data_232,
  output [7:0]  io_pipe_phv_out_data_233,
  output [7:0]  io_pipe_phv_out_data_234,
  output [7:0]  io_pipe_phv_out_data_235,
  output [7:0]  io_pipe_phv_out_data_236,
  output [7:0]  io_pipe_phv_out_data_237,
  output [7:0]  io_pipe_phv_out_data_238,
  output [7:0]  io_pipe_phv_out_data_239,
  output [7:0]  io_pipe_phv_out_data_240,
  output [7:0]  io_pipe_phv_out_data_241,
  output [7:0]  io_pipe_phv_out_data_242,
  output [7:0]  io_pipe_phv_out_data_243,
  output [7:0]  io_pipe_phv_out_data_244,
  output [7:0]  io_pipe_phv_out_data_245,
  output [7:0]  io_pipe_phv_out_data_246,
  output [7:0]  io_pipe_phv_out_data_247,
  output [7:0]  io_pipe_phv_out_data_248,
  output [7:0]  io_pipe_phv_out_data_249,
  output [7:0]  io_pipe_phv_out_data_250,
  output [7:0]  io_pipe_phv_out_data_251,
  output [7:0]  io_pipe_phv_out_data_252,
  output [7:0]  io_pipe_phv_out_data_253,
  output [7:0]  io_pipe_phv_out_data_254,
  output [7:0]  io_pipe_phv_out_data_255,
  output [7:0]  io_pipe_phv_out_data_256,
  output [7:0]  io_pipe_phv_out_data_257,
  output [7:0]  io_pipe_phv_out_data_258,
  output [7:0]  io_pipe_phv_out_data_259,
  output [7:0]  io_pipe_phv_out_data_260,
  output [7:0]  io_pipe_phv_out_data_261,
  output [7:0]  io_pipe_phv_out_data_262,
  output [7:0]  io_pipe_phv_out_data_263,
  output [7:0]  io_pipe_phv_out_data_264,
  output [7:0]  io_pipe_phv_out_data_265,
  output [7:0]  io_pipe_phv_out_data_266,
  output [7:0]  io_pipe_phv_out_data_267,
  output [7:0]  io_pipe_phv_out_data_268,
  output [7:0]  io_pipe_phv_out_data_269,
  output [7:0]  io_pipe_phv_out_data_270,
  output [7:0]  io_pipe_phv_out_data_271,
  output [7:0]  io_pipe_phv_out_data_272,
  output [7:0]  io_pipe_phv_out_data_273,
  output [7:0]  io_pipe_phv_out_data_274,
  output [7:0]  io_pipe_phv_out_data_275,
  output [7:0]  io_pipe_phv_out_data_276,
  output [7:0]  io_pipe_phv_out_data_277,
  output [7:0]  io_pipe_phv_out_data_278,
  output [7:0]  io_pipe_phv_out_data_279,
  output [7:0]  io_pipe_phv_out_data_280,
  output [7:0]  io_pipe_phv_out_data_281,
  output [7:0]  io_pipe_phv_out_data_282,
  output [7:0]  io_pipe_phv_out_data_283,
  output [7:0]  io_pipe_phv_out_data_284,
  output [7:0]  io_pipe_phv_out_data_285,
  output [7:0]  io_pipe_phv_out_data_286,
  output [7:0]  io_pipe_phv_out_data_287,
  output [7:0]  io_pipe_phv_out_data_288,
  output [7:0]  io_pipe_phv_out_data_289,
  output [7:0]  io_pipe_phv_out_data_290,
  output [7:0]  io_pipe_phv_out_data_291,
  output [7:0]  io_pipe_phv_out_data_292,
  output [7:0]  io_pipe_phv_out_data_293,
  output [7:0]  io_pipe_phv_out_data_294,
  output [7:0]  io_pipe_phv_out_data_295,
  output [7:0]  io_pipe_phv_out_data_296,
  output [7:0]  io_pipe_phv_out_data_297,
  output [7:0]  io_pipe_phv_out_data_298,
  output [7:0]  io_pipe_phv_out_data_299,
  output [7:0]  io_pipe_phv_out_data_300,
  output [7:0]  io_pipe_phv_out_data_301,
  output [7:0]  io_pipe_phv_out_data_302,
  output [7:0]  io_pipe_phv_out_data_303,
  output [7:0]  io_pipe_phv_out_data_304,
  output [7:0]  io_pipe_phv_out_data_305,
  output [7:0]  io_pipe_phv_out_data_306,
  output [7:0]  io_pipe_phv_out_data_307,
  output [7:0]  io_pipe_phv_out_data_308,
  output [7:0]  io_pipe_phv_out_data_309,
  output [7:0]  io_pipe_phv_out_data_310,
  output [7:0]  io_pipe_phv_out_data_311,
  output [7:0]  io_pipe_phv_out_data_312,
  output [7:0]  io_pipe_phv_out_data_313,
  output [7:0]  io_pipe_phv_out_data_314,
  output [7:0]  io_pipe_phv_out_data_315,
  output [7:0]  io_pipe_phv_out_data_316,
  output [7:0]  io_pipe_phv_out_data_317,
  output [7:0]  io_pipe_phv_out_data_318,
  output [7:0]  io_pipe_phv_out_data_319,
  output [7:0]  io_pipe_phv_out_data_320,
  output [7:0]  io_pipe_phv_out_data_321,
  output [7:0]  io_pipe_phv_out_data_322,
  output [7:0]  io_pipe_phv_out_data_323,
  output [7:0]  io_pipe_phv_out_data_324,
  output [7:0]  io_pipe_phv_out_data_325,
  output [7:0]  io_pipe_phv_out_data_326,
  output [7:0]  io_pipe_phv_out_data_327,
  output [7:0]  io_pipe_phv_out_data_328,
  output [7:0]  io_pipe_phv_out_data_329,
  output [7:0]  io_pipe_phv_out_data_330,
  output [7:0]  io_pipe_phv_out_data_331,
  output [7:0]  io_pipe_phv_out_data_332,
  output [7:0]  io_pipe_phv_out_data_333,
  output [7:0]  io_pipe_phv_out_data_334,
  output [7:0]  io_pipe_phv_out_data_335,
  output [7:0]  io_pipe_phv_out_data_336,
  output [7:0]  io_pipe_phv_out_data_337,
  output [7:0]  io_pipe_phv_out_data_338,
  output [7:0]  io_pipe_phv_out_data_339,
  output [7:0]  io_pipe_phv_out_data_340,
  output [7:0]  io_pipe_phv_out_data_341,
  output [7:0]  io_pipe_phv_out_data_342,
  output [7:0]  io_pipe_phv_out_data_343,
  output [7:0]  io_pipe_phv_out_data_344,
  output [7:0]  io_pipe_phv_out_data_345,
  output [7:0]  io_pipe_phv_out_data_346,
  output [7:0]  io_pipe_phv_out_data_347,
  output [7:0]  io_pipe_phv_out_data_348,
  output [7:0]  io_pipe_phv_out_data_349,
  output [7:0]  io_pipe_phv_out_data_350,
  output [7:0]  io_pipe_phv_out_data_351,
  output [7:0]  io_pipe_phv_out_data_352,
  output [7:0]  io_pipe_phv_out_data_353,
  output [7:0]  io_pipe_phv_out_data_354,
  output [7:0]  io_pipe_phv_out_data_355,
  output [7:0]  io_pipe_phv_out_data_356,
  output [7:0]  io_pipe_phv_out_data_357,
  output [7:0]  io_pipe_phv_out_data_358,
  output [7:0]  io_pipe_phv_out_data_359,
  output [7:0]  io_pipe_phv_out_data_360,
  output [7:0]  io_pipe_phv_out_data_361,
  output [7:0]  io_pipe_phv_out_data_362,
  output [7:0]  io_pipe_phv_out_data_363,
  output [7:0]  io_pipe_phv_out_data_364,
  output [7:0]  io_pipe_phv_out_data_365,
  output [7:0]  io_pipe_phv_out_data_366,
  output [7:0]  io_pipe_phv_out_data_367,
  output [7:0]  io_pipe_phv_out_data_368,
  output [7:0]  io_pipe_phv_out_data_369,
  output [7:0]  io_pipe_phv_out_data_370,
  output [7:0]  io_pipe_phv_out_data_371,
  output [7:0]  io_pipe_phv_out_data_372,
  output [7:0]  io_pipe_phv_out_data_373,
  output [7:0]  io_pipe_phv_out_data_374,
  output [7:0]  io_pipe_phv_out_data_375,
  output [7:0]  io_pipe_phv_out_data_376,
  output [7:0]  io_pipe_phv_out_data_377,
  output [7:0]  io_pipe_phv_out_data_378,
  output [7:0]  io_pipe_phv_out_data_379,
  output [7:0]  io_pipe_phv_out_data_380,
  output [7:0]  io_pipe_phv_out_data_381,
  output [7:0]  io_pipe_phv_out_data_382,
  output [7:0]  io_pipe_phv_out_data_383,
  output [7:0]  io_pipe_phv_out_data_384,
  output [7:0]  io_pipe_phv_out_data_385,
  output [7:0]  io_pipe_phv_out_data_386,
  output [7:0]  io_pipe_phv_out_data_387,
  output [7:0]  io_pipe_phv_out_data_388,
  output [7:0]  io_pipe_phv_out_data_389,
  output [7:0]  io_pipe_phv_out_data_390,
  output [7:0]  io_pipe_phv_out_data_391,
  output [7:0]  io_pipe_phv_out_data_392,
  output [7:0]  io_pipe_phv_out_data_393,
  output [7:0]  io_pipe_phv_out_data_394,
  output [7:0]  io_pipe_phv_out_data_395,
  output [7:0]  io_pipe_phv_out_data_396,
  output [7:0]  io_pipe_phv_out_data_397,
  output [7:0]  io_pipe_phv_out_data_398,
  output [7:0]  io_pipe_phv_out_data_399,
  output [7:0]  io_pipe_phv_out_data_400,
  output [7:0]  io_pipe_phv_out_data_401,
  output [7:0]  io_pipe_phv_out_data_402,
  output [7:0]  io_pipe_phv_out_data_403,
  output [7:0]  io_pipe_phv_out_data_404,
  output [7:0]  io_pipe_phv_out_data_405,
  output [7:0]  io_pipe_phv_out_data_406,
  output [7:0]  io_pipe_phv_out_data_407,
  output [7:0]  io_pipe_phv_out_data_408,
  output [7:0]  io_pipe_phv_out_data_409,
  output [7:0]  io_pipe_phv_out_data_410,
  output [7:0]  io_pipe_phv_out_data_411,
  output [7:0]  io_pipe_phv_out_data_412,
  output [7:0]  io_pipe_phv_out_data_413,
  output [7:0]  io_pipe_phv_out_data_414,
  output [7:0]  io_pipe_phv_out_data_415,
  output [7:0]  io_pipe_phv_out_data_416,
  output [7:0]  io_pipe_phv_out_data_417,
  output [7:0]  io_pipe_phv_out_data_418,
  output [7:0]  io_pipe_phv_out_data_419,
  output [7:0]  io_pipe_phv_out_data_420,
  output [7:0]  io_pipe_phv_out_data_421,
  output [7:0]  io_pipe_phv_out_data_422,
  output [7:0]  io_pipe_phv_out_data_423,
  output [7:0]  io_pipe_phv_out_data_424,
  output [7:0]  io_pipe_phv_out_data_425,
  output [7:0]  io_pipe_phv_out_data_426,
  output [7:0]  io_pipe_phv_out_data_427,
  output [7:0]  io_pipe_phv_out_data_428,
  output [7:0]  io_pipe_phv_out_data_429,
  output [7:0]  io_pipe_phv_out_data_430,
  output [7:0]  io_pipe_phv_out_data_431,
  output [7:0]  io_pipe_phv_out_data_432,
  output [7:0]  io_pipe_phv_out_data_433,
  output [7:0]  io_pipe_phv_out_data_434,
  output [7:0]  io_pipe_phv_out_data_435,
  output [7:0]  io_pipe_phv_out_data_436,
  output [7:0]  io_pipe_phv_out_data_437,
  output [7:0]  io_pipe_phv_out_data_438,
  output [7:0]  io_pipe_phv_out_data_439,
  output [7:0]  io_pipe_phv_out_data_440,
  output [7:0]  io_pipe_phv_out_data_441,
  output [7:0]  io_pipe_phv_out_data_442,
  output [7:0]  io_pipe_phv_out_data_443,
  output [7:0]  io_pipe_phv_out_data_444,
  output [7:0]  io_pipe_phv_out_data_445,
  output [7:0]  io_pipe_phv_out_data_446,
  output [7:0]  io_pipe_phv_out_data_447,
  output [7:0]  io_pipe_phv_out_data_448,
  output [7:0]  io_pipe_phv_out_data_449,
  output [7:0]  io_pipe_phv_out_data_450,
  output [7:0]  io_pipe_phv_out_data_451,
  output [7:0]  io_pipe_phv_out_data_452,
  output [7:0]  io_pipe_phv_out_data_453,
  output [7:0]  io_pipe_phv_out_data_454,
  output [7:0]  io_pipe_phv_out_data_455,
  output [7:0]  io_pipe_phv_out_data_456,
  output [7:0]  io_pipe_phv_out_data_457,
  output [7:0]  io_pipe_phv_out_data_458,
  output [7:0]  io_pipe_phv_out_data_459,
  output [7:0]  io_pipe_phv_out_data_460,
  output [7:0]  io_pipe_phv_out_data_461,
  output [7:0]  io_pipe_phv_out_data_462,
  output [7:0]  io_pipe_phv_out_data_463,
  output [7:0]  io_pipe_phv_out_data_464,
  output [7:0]  io_pipe_phv_out_data_465,
  output [7:0]  io_pipe_phv_out_data_466,
  output [7:0]  io_pipe_phv_out_data_467,
  output [7:0]  io_pipe_phv_out_data_468,
  output [7:0]  io_pipe_phv_out_data_469,
  output [7:0]  io_pipe_phv_out_data_470,
  output [7:0]  io_pipe_phv_out_data_471,
  output [7:0]  io_pipe_phv_out_data_472,
  output [7:0]  io_pipe_phv_out_data_473,
  output [7:0]  io_pipe_phv_out_data_474,
  output [7:0]  io_pipe_phv_out_data_475,
  output [7:0]  io_pipe_phv_out_data_476,
  output [7:0]  io_pipe_phv_out_data_477,
  output [7:0]  io_pipe_phv_out_data_478,
  output [7:0]  io_pipe_phv_out_data_479,
  output [7:0]  io_pipe_phv_out_data_480,
  output [7:0]  io_pipe_phv_out_data_481,
  output [7:0]  io_pipe_phv_out_data_482,
  output [7:0]  io_pipe_phv_out_data_483,
  output [7:0]  io_pipe_phv_out_data_484,
  output [7:0]  io_pipe_phv_out_data_485,
  output [7:0]  io_pipe_phv_out_data_486,
  output [7:0]  io_pipe_phv_out_data_487,
  output [7:0]  io_pipe_phv_out_data_488,
  output [7:0]  io_pipe_phv_out_data_489,
  output [7:0]  io_pipe_phv_out_data_490,
  output [7:0]  io_pipe_phv_out_data_491,
  output [7:0]  io_pipe_phv_out_data_492,
  output [7:0]  io_pipe_phv_out_data_493,
  output [7:0]  io_pipe_phv_out_data_494,
  output [7:0]  io_pipe_phv_out_data_495,
  output [7:0]  io_pipe_phv_out_data_496,
  output [7:0]  io_pipe_phv_out_data_497,
  output [7:0]  io_pipe_phv_out_data_498,
  output [7:0]  io_pipe_phv_out_data_499,
  output [7:0]  io_pipe_phv_out_data_500,
  output [7:0]  io_pipe_phv_out_data_501,
  output [7:0]  io_pipe_phv_out_data_502,
  output [7:0]  io_pipe_phv_out_data_503,
  output [7:0]  io_pipe_phv_out_data_504,
  output [7:0]  io_pipe_phv_out_data_505,
  output [7:0]  io_pipe_phv_out_data_506,
  output [7:0]  io_pipe_phv_out_data_507,
  output [7:0]  io_pipe_phv_out_data_508,
  output [7:0]  io_pipe_phv_out_data_509,
  output [7:0]  io_pipe_phv_out_data_510,
  output [7:0]  io_pipe_phv_out_data_511,
  output [15:0] io_pipe_phv_out_header_0,
  output [15:0] io_pipe_phv_out_header_1,
  output [15:0] io_pipe_phv_out_header_2,
  output [15:0] io_pipe_phv_out_header_3,
  output [15:0] io_pipe_phv_out_header_4,
  output [15:0] io_pipe_phv_out_header_5,
  output [15:0] io_pipe_phv_out_header_6,
  output [15:0] io_pipe_phv_out_header_7,
  output [15:0] io_pipe_phv_out_header_8,
  output [15:0] io_pipe_phv_out_header_9,
  output [15:0] io_pipe_phv_out_header_10,
  output [15:0] io_pipe_phv_out_header_11,
  output [15:0] io_pipe_phv_out_header_12,
  output [15:0] io_pipe_phv_out_header_13,
  output [15:0] io_pipe_phv_out_header_14,
  output [15:0] io_pipe_phv_out_header_15,
  output [7:0]  io_pipe_phv_out_parse_current_state,
  output [7:0]  io_pipe_phv_out_parse_current_offset,
  output [15:0] io_pipe_phv_out_parse_transition_field,
  output [3:0]  io_pipe_phv_out_next_processor_id,
  output        io_pipe_phv_out_next_config_id,
  input         io_hit,
  input  [63:0] io_match_value,
  input         io_action_mod_en_0,
  input         io_action_mod_en_1,
  input  [7:0]  io_action_mod_addr,
  input  [63:0] io_action_mod_data_0,
  input  [63:0] io_action_mod_data_1
);
  wire  pipe1_clock; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_0; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_2; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_3; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_4; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_5; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_6; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_7; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_8; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_9; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_10; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_11; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_12; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_13; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_14; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_16; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_17; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_18; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_19; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_20; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_21; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_22; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_23; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_24; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_25; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_26; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_27; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_28; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_29; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_30; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_31; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_32; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_33; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_34; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_35; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_36; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_37; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_38; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_39; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_40; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_41; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_42; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_43; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_44; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_45; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_46; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_47; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_48; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_49; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_50; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_51; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_52; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_53; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_54; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_55; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_56; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_57; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_58; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_59; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_60; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_61; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_62; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_63; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_64; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_65; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_66; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_67; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_68; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_69; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_70; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_71; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_72; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_73; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_74; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_75; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_76; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_77; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_78; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_79; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_80; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_81; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_82; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_83; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_84; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_85; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_86; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_87; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_88; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_89; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_90; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_91; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_92; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_93; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_94; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_95; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_96; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_97; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_98; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_99; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_100; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_101; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_102; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_103; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_104; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_105; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_106; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_107; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_108; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_109; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_110; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_111; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_112; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_113; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_114; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_115; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_116; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_117; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_118; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_119; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_120; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_121; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_122; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_123; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_124; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_125; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_126; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_127; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_128; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_129; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_130; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_131; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_132; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_133; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_134; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_135; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_136; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_137; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_138; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_139; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_140; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_141; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_142; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_143; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_144; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_145; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_146; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_147; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_148; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_149; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_150; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_151; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_152; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_153; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_154; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_155; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_156; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_157; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_158; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_159; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_160; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_161; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_162; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_163; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_164; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_165; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_166; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_167; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_168; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_169; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_170; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_171; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_172; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_173; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_174; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_175; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_176; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_177; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_178; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_179; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_180; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_181; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_182; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_183; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_184; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_185; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_186; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_187; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_188; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_189; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_190; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_191; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_192; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_193; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_194; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_195; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_196; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_197; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_198; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_199; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_200; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_201; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_202; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_203; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_204; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_205; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_206; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_207; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_208; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_209; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_210; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_211; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_212; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_213; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_214; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_215; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_216; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_217; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_218; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_219; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_220; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_221; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_222; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_223; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_224; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_225; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_226; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_227; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_228; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_229; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_230; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_231; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_232; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_233; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_234; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_235; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_236; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_237; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_238; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_239; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_240; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_241; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_242; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_243; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_244; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_245; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_246; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_247; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_248; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_249; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_250; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_251; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_252; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_253; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_254; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_255; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_256; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_257; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_258; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_259; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_260; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_261; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_262; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_263; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_264; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_265; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_266; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_267; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_268; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_269; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_270; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_271; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_272; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_273; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_274; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_275; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_276; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_277; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_278; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_279; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_280; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_281; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_282; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_283; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_284; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_285; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_286; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_287; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_288; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_289; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_290; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_291; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_292; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_293; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_294; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_295; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_296; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_297; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_298; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_299; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_300; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_301; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_302; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_303; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_304; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_305; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_306; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_307; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_308; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_309; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_310; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_311; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_312; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_313; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_314; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_315; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_316; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_317; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_318; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_319; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_320; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_321; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_322; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_323; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_324; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_325; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_326; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_327; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_328; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_329; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_330; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_331; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_332; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_333; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_334; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_335; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_336; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_337; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_338; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_339; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_340; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_341; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_342; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_343; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_344; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_345; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_346; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_347; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_348; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_349; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_350; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_351; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_352; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_353; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_354; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_355; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_356; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_357; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_358; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_359; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_360; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_361; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_362; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_363; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_364; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_365; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_366; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_367; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_368; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_369; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_370; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_371; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_372; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_373; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_374; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_375; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_376; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_377; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_378; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_379; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_380; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_381; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_382; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_383; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_384; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_385; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_386; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_387; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_388; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_389; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_390; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_391; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_392; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_393; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_394; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_395; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_396; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_397; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_398; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_399; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_400; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_401; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_402; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_403; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_404; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_405; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_406; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_407; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_408; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_409; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_410; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_411; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_412; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_413; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_414; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_415; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_416; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_417; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_418; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_419; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_420; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_421; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_422; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_423; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_424; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_425; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_426; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_427; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_428; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_429; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_430; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_431; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_432; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_433; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_434; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_435; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_436; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_437; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_438; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_439; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_440; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_441; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_442; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_443; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_444; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_445; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_446; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_447; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_448; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_449; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_450; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_451; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_452; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_453; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_454; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_455; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_456; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_457; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_458; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_459; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_460; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_461; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_462; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_463; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_464; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_465; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_466; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_467; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_468; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_469; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_470; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_471; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_472; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_473; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_474; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_475; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_476; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_477; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_478; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_479; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_480; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_481; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_482; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_483; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_484; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_485; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_486; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_487; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_488; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_489; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_490; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_491; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_492; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_493; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_494; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_495; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_496; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_497; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_498; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_499; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_500; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_501; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_502; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_503; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_504; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_505; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_506; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_507; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_508; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_509; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_510; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_data_511; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_0; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_1; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_2; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_3; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_4; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_5; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_6; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_7; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_8; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_9; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_10; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_11; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_12; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_13; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_14; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_header_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_state; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_in_parse_current_offset; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_in_parse_transition_field; // @[executor.scala 489:23]
  wire [3:0] pipe1_io_pipe_phv_in_next_processor_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_in_next_config_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_in_is_valid_processor; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_0; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_2; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_3; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_4; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_5; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_6; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_7; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_8; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_9; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_10; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_11; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_12; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_13; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_14; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_16; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_17; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_18; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_19; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_20; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_21; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_22; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_23; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_24; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_25; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_26; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_27; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_28; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_29; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_30; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_31; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_32; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_33; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_34; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_35; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_36; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_37; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_38; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_39; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_40; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_41; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_42; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_43; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_44; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_45; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_46; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_47; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_48; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_49; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_50; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_51; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_52; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_53; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_54; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_55; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_56; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_57; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_58; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_59; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_60; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_61; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_62; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_63; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_64; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_65; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_66; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_67; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_68; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_69; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_70; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_71; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_72; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_73; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_74; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_75; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_76; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_77; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_78; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_79; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_80; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_81; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_82; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_83; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_84; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_85; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_86; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_87; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_88; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_89; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_90; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_91; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_92; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_93; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_94; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_95; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_96; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_97; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_98; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_99; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_100; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_101; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_102; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_103; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_104; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_105; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_106; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_107; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_108; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_109; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_110; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_111; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_112; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_113; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_114; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_115; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_116; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_117; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_118; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_119; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_120; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_121; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_122; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_123; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_124; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_125; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_126; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_127; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_128; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_129; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_130; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_131; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_132; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_133; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_134; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_135; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_136; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_137; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_138; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_139; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_140; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_141; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_142; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_143; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_144; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_145; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_146; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_147; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_148; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_149; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_150; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_151; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_152; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_153; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_154; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_155; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_156; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_157; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_158; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_159; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_160; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_161; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_162; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_163; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_164; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_165; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_166; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_167; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_168; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_169; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_170; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_171; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_172; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_173; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_174; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_175; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_176; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_177; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_178; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_179; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_180; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_181; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_182; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_183; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_184; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_185; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_186; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_187; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_188; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_189; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_190; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_191; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_192; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_193; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_194; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_195; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_196; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_197; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_198; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_199; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_200; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_201; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_202; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_203; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_204; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_205; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_206; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_207; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_208; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_209; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_210; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_211; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_212; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_213; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_214; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_215; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_216; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_217; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_218; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_219; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_220; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_221; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_222; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_223; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_224; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_225; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_226; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_227; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_228; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_229; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_230; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_231; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_232; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_233; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_234; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_235; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_236; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_237; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_238; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_239; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_240; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_241; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_242; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_243; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_244; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_245; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_246; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_247; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_248; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_249; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_250; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_251; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_252; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_253; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_254; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_255; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_256; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_257; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_258; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_259; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_260; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_261; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_262; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_263; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_264; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_265; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_266; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_267; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_268; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_269; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_270; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_271; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_272; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_273; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_274; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_275; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_276; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_277; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_278; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_279; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_280; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_281; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_282; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_283; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_284; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_285; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_286; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_287; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_288; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_289; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_290; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_291; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_292; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_293; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_294; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_295; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_296; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_297; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_298; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_299; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_300; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_301; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_302; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_303; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_304; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_305; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_306; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_307; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_308; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_309; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_310; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_311; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_312; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_313; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_314; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_315; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_316; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_317; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_318; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_319; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_320; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_321; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_322; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_323; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_324; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_325; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_326; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_327; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_328; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_329; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_330; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_331; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_332; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_333; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_334; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_335; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_336; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_337; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_338; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_339; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_340; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_341; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_342; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_343; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_344; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_345; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_346; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_347; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_348; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_349; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_350; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_351; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_352; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_353; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_354; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_355; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_356; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_357; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_358; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_359; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_360; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_361; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_362; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_363; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_364; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_365; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_366; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_367; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_368; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_369; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_370; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_371; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_372; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_373; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_374; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_375; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_376; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_377; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_378; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_379; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_380; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_381; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_382; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_383; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_384; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_385; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_386; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_387; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_388; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_389; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_390; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_391; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_392; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_393; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_394; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_395; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_396; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_397; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_398; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_399; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_400; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_401; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_402; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_403; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_404; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_405; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_406; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_407; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_408; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_409; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_410; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_411; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_412; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_413; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_414; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_415; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_416; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_417; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_418; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_419; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_420; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_421; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_422; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_423; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_424; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_425; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_426; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_427; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_428; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_429; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_430; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_431; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_432; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_433; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_434; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_435; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_436; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_437; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_438; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_439; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_440; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_441; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_442; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_443; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_444; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_445; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_446; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_447; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_448; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_449; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_450; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_451; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_452; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_453; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_454; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_455; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_456; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_457; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_458; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_459; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_460; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_461; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_462; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_463; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_464; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_465; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_466; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_467; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_468; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_469; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_470; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_471; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_472; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_473; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_474; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_475; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_476; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_477; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_478; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_479; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_480; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_481; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_482; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_483; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_484; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_485; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_486; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_487; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_488; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_489; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_490; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_491; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_492; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_493; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_494; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_495; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_496; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_497; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_498; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_499; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_500; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_501; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_502; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_503; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_504; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_505; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_506; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_507; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_508; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_509; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_510; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_data_511; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_0; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_1; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_2; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_3; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_4; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_5; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_6; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_7; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_8; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_9; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_10; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_11; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_12; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_13; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_14; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_header_15; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 489:23]
  wire [15:0] pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 489:23]
  wire [3:0] pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_out_next_config_id; // @[executor.scala 489:23]
  wire  pipe1_io_pipe_phv_out_is_valid_processor; // @[executor.scala 489:23]
  wire  pipe1_io_hit; // @[executor.scala 489:23]
  wire [63:0] pipe1_io_match_value; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_0; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_2; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_3; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_4; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_5; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_args_out_6; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_0; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_1; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_2; // @[executor.scala 489:23]
  wire [31:0] pipe1_io_vliw_out_3; // @[executor.scala 489:23]
  wire  pipe1_io_action_mod_en_0; // @[executor.scala 489:23]
  wire  pipe1_io_action_mod_en_1; // @[executor.scala 489:23]
  wire [7:0] pipe1_io_action_mod_addr; // @[executor.scala 489:23]
  wire [63:0] pipe1_io_action_mod_data_0; // @[executor.scala 489:23]
  wire [63:0] pipe1_io_action_mod_data_1; // @[executor.scala 489:23]
  wire  pipe2_clock; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_6; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_7; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_8; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_9; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_10; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_11; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_12; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_13; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_14; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_16; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_17; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_18; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_19; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_20; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_21; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_22; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_23; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_24; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_25; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_26; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_27; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_28; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_29; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_30; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_31; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_32; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_33; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_34; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_35; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_36; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_37; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_38; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_39; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_40; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_41; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_42; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_43; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_44; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_45; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_46; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_47; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_48; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_49; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_50; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_51; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_52; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_53; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_54; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_55; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_56; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_57; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_58; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_59; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_60; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_61; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_62; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_63; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_64; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_65; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_66; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_67; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_68; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_69; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_70; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_71; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_72; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_73; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_74; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_75; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_76; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_77; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_78; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_79; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_80; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_81; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_82; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_83; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_84; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_85; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_86; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_87; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_88; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_89; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_90; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_91; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_92; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_93; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_94; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_95; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_96; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_97; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_98; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_99; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_100; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_101; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_102; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_103; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_104; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_105; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_106; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_107; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_108; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_109; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_110; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_111; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_112; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_113; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_114; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_115; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_116; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_117; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_118; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_119; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_120; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_121; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_122; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_123; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_124; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_125; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_126; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_127; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_128; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_129; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_130; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_131; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_132; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_133; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_134; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_135; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_136; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_137; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_138; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_139; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_140; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_141; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_142; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_143; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_144; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_145; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_146; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_147; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_148; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_149; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_150; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_151; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_152; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_153; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_154; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_155; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_156; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_157; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_158; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_159; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_160; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_161; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_162; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_163; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_164; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_165; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_166; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_167; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_168; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_169; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_170; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_171; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_172; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_173; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_174; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_175; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_176; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_177; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_178; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_179; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_180; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_181; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_182; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_183; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_184; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_185; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_186; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_187; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_188; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_189; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_190; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_191; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_192; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_193; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_194; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_195; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_196; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_197; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_198; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_199; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_200; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_201; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_202; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_203; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_204; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_205; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_206; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_207; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_208; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_209; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_210; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_211; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_212; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_213; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_214; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_215; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_216; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_217; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_218; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_219; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_220; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_221; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_222; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_223; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_224; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_225; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_226; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_227; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_228; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_229; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_230; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_231; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_232; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_233; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_234; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_235; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_236; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_237; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_238; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_239; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_240; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_241; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_242; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_243; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_244; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_245; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_246; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_247; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_248; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_249; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_250; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_251; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_252; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_253; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_254; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_255; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_256; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_257; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_258; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_259; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_260; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_261; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_262; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_263; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_264; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_265; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_266; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_267; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_268; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_269; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_270; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_271; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_272; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_273; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_274; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_275; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_276; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_277; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_278; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_279; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_280; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_281; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_282; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_283; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_284; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_285; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_286; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_287; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_288; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_289; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_290; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_291; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_292; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_293; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_294; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_295; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_296; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_297; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_298; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_299; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_300; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_301; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_302; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_303; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_304; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_305; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_306; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_307; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_308; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_309; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_310; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_311; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_312; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_313; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_314; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_315; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_316; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_317; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_318; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_319; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_320; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_321; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_322; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_323; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_324; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_325; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_326; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_327; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_328; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_329; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_330; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_331; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_332; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_333; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_334; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_335; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_336; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_337; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_338; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_339; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_340; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_341; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_342; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_343; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_344; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_345; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_346; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_347; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_348; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_349; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_350; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_351; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_352; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_353; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_354; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_355; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_356; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_357; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_358; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_359; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_360; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_361; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_362; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_363; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_364; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_365; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_366; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_367; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_368; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_369; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_370; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_371; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_372; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_373; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_374; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_375; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_376; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_377; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_378; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_379; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_380; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_381; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_382; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_383; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_384; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_385; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_386; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_387; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_388; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_389; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_390; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_391; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_392; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_393; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_394; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_395; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_396; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_397; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_398; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_399; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_400; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_401; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_402; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_403; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_404; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_405; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_406; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_407; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_408; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_409; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_410; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_411; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_412; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_413; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_414; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_415; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_416; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_417; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_418; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_419; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_420; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_421; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_422; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_423; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_424; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_425; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_426; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_427; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_428; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_429; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_430; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_431; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_432; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_433; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_434; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_435; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_436; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_437; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_438; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_439; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_440; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_441; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_442; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_443; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_444; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_445; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_446; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_447; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_448; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_449; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_450; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_451; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_452; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_453; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_454; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_455; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_456; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_457; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_458; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_459; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_460; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_461; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_462; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_463; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_464; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_465; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_466; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_467; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_468; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_469; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_470; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_471; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_472; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_473; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_474; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_475; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_476; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_477; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_478; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_479; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_480; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_481; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_482; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_483; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_484; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_485; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_486; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_487; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_488; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_489; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_490; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_491; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_492; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_493; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_494; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_495; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_496; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_497; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_498; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_499; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_500; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_501; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_502; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_503; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_504; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_505; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_506; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_507; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_508; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_509; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_510; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_data_511; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_0; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_1; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_2; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_3; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_4; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_5; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_6; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_7; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_8; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_9; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_10; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_11; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_12; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_13; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_14; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_header_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_state; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_in_parse_current_offset; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_in_parse_transition_field; // @[executor.scala 490:23]
  wire [3:0] pipe2_io_pipe_phv_in_next_processor_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_in_next_config_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_in_is_valid_processor; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_6; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_7; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_8; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_9; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_10; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_11; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_12; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_13; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_14; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_16; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_17; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_18; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_19; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_20; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_21; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_22; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_23; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_24; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_25; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_26; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_27; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_28; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_29; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_30; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_31; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_32; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_33; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_34; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_35; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_36; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_37; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_38; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_39; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_40; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_41; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_42; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_43; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_44; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_45; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_46; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_47; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_48; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_49; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_50; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_51; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_52; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_53; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_54; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_55; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_56; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_57; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_58; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_59; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_60; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_61; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_62; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_63; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_64; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_65; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_66; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_67; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_68; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_69; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_70; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_71; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_72; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_73; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_74; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_75; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_76; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_77; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_78; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_79; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_80; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_81; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_82; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_83; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_84; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_85; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_86; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_87; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_88; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_89; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_90; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_91; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_92; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_93; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_94; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_95; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_96; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_97; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_98; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_99; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_100; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_101; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_102; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_103; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_104; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_105; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_106; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_107; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_108; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_109; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_110; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_111; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_112; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_113; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_114; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_115; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_116; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_117; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_118; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_119; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_120; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_121; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_122; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_123; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_124; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_125; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_126; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_127; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_128; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_129; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_130; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_131; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_132; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_133; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_134; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_135; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_136; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_137; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_138; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_139; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_140; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_141; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_142; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_143; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_144; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_145; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_146; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_147; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_148; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_149; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_150; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_151; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_152; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_153; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_154; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_155; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_156; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_157; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_158; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_159; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_160; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_161; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_162; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_163; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_164; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_165; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_166; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_167; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_168; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_169; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_170; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_171; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_172; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_173; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_174; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_175; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_176; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_177; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_178; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_179; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_180; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_181; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_182; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_183; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_184; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_185; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_186; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_187; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_188; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_189; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_190; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_191; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_192; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_193; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_194; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_195; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_196; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_197; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_198; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_199; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_200; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_201; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_202; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_203; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_204; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_205; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_206; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_207; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_208; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_209; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_210; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_211; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_212; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_213; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_214; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_215; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_216; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_217; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_218; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_219; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_220; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_221; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_222; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_223; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_224; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_225; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_226; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_227; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_228; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_229; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_230; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_231; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_232; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_233; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_234; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_235; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_236; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_237; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_238; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_239; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_240; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_241; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_242; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_243; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_244; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_245; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_246; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_247; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_248; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_249; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_250; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_251; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_252; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_253; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_254; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_255; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_256; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_257; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_258; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_259; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_260; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_261; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_262; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_263; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_264; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_265; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_266; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_267; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_268; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_269; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_270; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_271; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_272; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_273; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_274; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_275; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_276; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_277; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_278; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_279; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_280; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_281; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_282; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_283; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_284; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_285; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_286; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_287; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_288; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_289; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_290; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_291; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_292; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_293; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_294; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_295; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_296; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_297; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_298; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_299; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_300; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_301; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_302; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_303; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_304; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_305; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_306; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_307; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_308; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_309; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_310; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_311; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_312; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_313; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_314; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_315; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_316; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_317; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_318; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_319; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_320; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_321; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_322; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_323; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_324; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_325; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_326; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_327; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_328; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_329; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_330; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_331; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_332; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_333; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_334; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_335; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_336; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_337; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_338; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_339; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_340; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_341; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_342; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_343; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_344; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_345; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_346; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_347; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_348; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_349; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_350; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_351; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_352; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_353; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_354; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_355; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_356; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_357; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_358; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_359; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_360; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_361; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_362; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_363; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_364; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_365; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_366; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_367; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_368; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_369; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_370; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_371; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_372; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_373; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_374; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_375; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_376; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_377; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_378; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_379; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_380; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_381; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_382; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_383; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_384; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_385; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_386; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_387; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_388; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_389; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_390; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_391; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_392; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_393; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_394; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_395; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_396; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_397; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_398; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_399; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_400; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_401; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_402; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_403; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_404; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_405; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_406; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_407; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_408; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_409; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_410; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_411; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_412; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_413; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_414; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_415; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_416; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_417; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_418; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_419; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_420; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_421; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_422; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_423; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_424; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_425; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_426; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_427; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_428; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_429; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_430; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_431; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_432; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_433; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_434; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_435; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_436; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_437; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_438; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_439; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_440; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_441; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_442; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_443; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_444; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_445; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_446; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_447; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_448; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_449; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_450; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_451; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_452; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_453; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_454; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_455; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_456; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_457; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_458; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_459; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_460; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_461; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_462; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_463; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_464; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_465; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_466; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_467; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_468; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_469; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_470; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_471; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_472; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_473; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_474; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_475; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_476; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_477; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_478; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_479; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_480; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_481; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_482; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_483; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_484; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_485; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_486; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_487; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_488; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_489; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_490; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_491; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_492; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_493; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_494; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_495; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_496; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_497; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_498; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_499; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_500; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_501; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_502; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_503; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_504; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_505; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_506; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_507; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_508; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_509; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_510; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_data_511; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_0; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_1; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_2; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_3; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_4; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_5; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_6; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_7; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_8; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_9; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_10; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_11; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_12; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_13; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_14; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_header_15; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 490:23]
  wire [15:0] pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 490:23]
  wire [3:0] pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_out_next_config_id; // @[executor.scala 490:23]
  wire  pipe2_io_pipe_phv_out_is_valid_processor; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_in_6; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_0; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_1; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_2; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_in_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_4; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_5; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_args_out_6; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_0; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_1; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_2; // @[executor.scala 490:23]
  wire [31:0] pipe2_io_vliw_out_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_offset_out_3; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_0; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_1; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_2; // @[executor.scala 490:23]
  wire [7:0] pipe2_io_length_out_3; // @[executor.scala 490:23]
  wire  pipe3_clock; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_4; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_5; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_6; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_7; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_8; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_9; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_10; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_11; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_12; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_13; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_14; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_16; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_17; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_18; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_19; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_20; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_21; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_22; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_23; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_24; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_25; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_26; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_27; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_28; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_29; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_30; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_31; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_32; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_33; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_34; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_35; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_36; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_37; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_38; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_39; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_40; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_41; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_42; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_43; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_44; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_45; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_46; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_47; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_48; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_49; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_50; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_51; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_52; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_53; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_54; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_55; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_56; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_57; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_58; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_59; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_60; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_61; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_62; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_63; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_64; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_65; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_66; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_67; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_68; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_69; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_70; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_71; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_72; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_73; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_74; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_75; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_76; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_77; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_78; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_79; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_80; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_81; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_82; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_83; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_84; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_85; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_86; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_87; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_88; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_89; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_90; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_91; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_92; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_93; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_94; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_95; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_96; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_97; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_98; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_99; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_100; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_101; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_102; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_103; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_104; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_105; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_106; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_107; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_108; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_109; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_110; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_111; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_112; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_113; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_114; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_115; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_116; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_117; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_118; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_119; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_120; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_121; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_122; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_123; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_124; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_125; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_126; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_127; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_128; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_129; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_130; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_131; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_132; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_133; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_134; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_135; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_136; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_137; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_138; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_139; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_140; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_141; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_142; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_143; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_144; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_145; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_146; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_147; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_148; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_149; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_150; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_151; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_152; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_153; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_154; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_155; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_156; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_157; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_158; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_159; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_160; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_161; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_162; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_163; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_164; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_165; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_166; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_167; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_168; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_169; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_170; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_171; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_172; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_173; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_174; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_175; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_176; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_177; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_178; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_179; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_180; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_181; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_182; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_183; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_184; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_185; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_186; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_187; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_188; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_189; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_190; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_191; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_192; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_193; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_194; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_195; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_196; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_197; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_198; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_199; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_200; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_201; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_202; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_203; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_204; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_205; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_206; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_207; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_208; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_209; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_210; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_211; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_212; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_213; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_214; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_215; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_216; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_217; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_218; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_219; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_220; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_221; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_222; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_223; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_224; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_225; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_226; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_227; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_228; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_229; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_230; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_231; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_232; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_233; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_234; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_235; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_236; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_237; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_238; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_239; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_240; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_241; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_242; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_243; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_244; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_245; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_246; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_247; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_248; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_249; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_250; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_251; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_252; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_253; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_254; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_255; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_256; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_257; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_258; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_259; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_260; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_261; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_262; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_263; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_264; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_265; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_266; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_267; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_268; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_269; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_270; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_271; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_272; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_273; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_274; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_275; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_276; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_277; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_278; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_279; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_280; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_281; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_282; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_283; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_284; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_285; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_286; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_287; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_288; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_289; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_290; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_291; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_292; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_293; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_294; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_295; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_296; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_297; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_298; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_299; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_300; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_301; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_302; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_303; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_304; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_305; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_306; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_307; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_308; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_309; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_310; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_311; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_312; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_313; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_314; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_315; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_316; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_317; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_318; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_319; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_320; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_321; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_322; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_323; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_324; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_325; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_326; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_327; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_328; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_329; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_330; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_331; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_332; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_333; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_334; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_335; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_336; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_337; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_338; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_339; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_340; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_341; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_342; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_343; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_344; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_345; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_346; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_347; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_348; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_349; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_350; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_351; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_352; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_353; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_354; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_355; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_356; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_357; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_358; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_359; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_360; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_361; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_362; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_363; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_364; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_365; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_366; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_367; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_368; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_369; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_370; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_371; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_372; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_373; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_374; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_375; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_376; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_377; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_378; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_379; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_380; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_381; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_382; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_383; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_384; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_385; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_386; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_387; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_388; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_389; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_390; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_391; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_392; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_393; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_394; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_395; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_396; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_397; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_398; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_399; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_400; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_401; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_402; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_403; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_404; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_405; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_406; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_407; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_408; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_409; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_410; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_411; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_412; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_413; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_414; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_415; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_416; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_417; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_418; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_419; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_420; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_421; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_422; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_423; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_424; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_425; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_426; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_427; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_428; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_429; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_430; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_431; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_432; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_433; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_434; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_435; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_436; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_437; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_438; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_439; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_440; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_441; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_442; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_443; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_444; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_445; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_446; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_447; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_448; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_449; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_450; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_451; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_452; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_453; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_454; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_455; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_456; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_457; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_458; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_459; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_460; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_461; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_462; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_463; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_464; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_465; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_466; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_467; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_468; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_469; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_470; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_471; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_472; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_473; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_474; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_475; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_476; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_477; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_478; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_479; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_480; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_481; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_482; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_483; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_484; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_485; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_486; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_487; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_488; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_489; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_490; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_491; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_492; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_493; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_494; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_495; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_496; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_497; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_498; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_499; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_500; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_501; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_502; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_503; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_504; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_505; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_506; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_507; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_508; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_509; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_510; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_data_511; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_0; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_1; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_2; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_3; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_4; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_5; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_6; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_7; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_8; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_9; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_10; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_11; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_12; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_13; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_14; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_header_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_state; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_in_parse_current_offset; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_in_parse_transition_field; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_pipe_phv_in_next_processor_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_in_next_config_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_in_is_valid_processor; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_4; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_5; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_6; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_7; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_8; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_9; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_10; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_11; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_12; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_13; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_14; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_16; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_17; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_18; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_19; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_20; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_21; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_22; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_23; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_24; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_25; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_26; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_27; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_28; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_29; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_30; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_31; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_32; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_33; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_34; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_35; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_36; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_37; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_38; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_39; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_40; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_41; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_42; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_43; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_44; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_45; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_46; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_47; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_48; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_49; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_50; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_51; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_52; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_53; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_54; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_55; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_56; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_57; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_58; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_59; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_60; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_61; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_62; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_63; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_64; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_65; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_66; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_67; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_68; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_69; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_70; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_71; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_72; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_73; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_74; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_75; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_76; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_77; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_78; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_79; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_80; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_81; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_82; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_83; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_84; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_85; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_86; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_87; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_88; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_89; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_90; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_91; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_92; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_93; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_94; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_95; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_96; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_97; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_98; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_99; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_100; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_101; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_102; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_103; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_104; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_105; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_106; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_107; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_108; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_109; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_110; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_111; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_112; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_113; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_114; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_115; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_116; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_117; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_118; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_119; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_120; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_121; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_122; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_123; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_124; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_125; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_126; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_127; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_128; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_129; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_130; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_131; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_132; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_133; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_134; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_135; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_136; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_137; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_138; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_139; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_140; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_141; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_142; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_143; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_144; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_145; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_146; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_147; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_148; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_149; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_150; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_151; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_152; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_153; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_154; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_155; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_156; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_157; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_158; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_159; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_160; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_161; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_162; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_163; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_164; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_165; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_166; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_167; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_168; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_169; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_170; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_171; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_172; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_173; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_174; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_175; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_176; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_177; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_178; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_179; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_180; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_181; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_182; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_183; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_184; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_185; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_186; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_187; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_188; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_189; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_190; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_191; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_192; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_193; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_194; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_195; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_196; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_197; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_198; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_199; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_200; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_201; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_202; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_203; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_204; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_205; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_206; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_207; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_208; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_209; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_210; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_211; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_212; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_213; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_214; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_215; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_216; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_217; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_218; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_219; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_220; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_221; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_222; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_223; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_224; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_225; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_226; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_227; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_228; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_229; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_230; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_231; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_232; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_233; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_234; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_235; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_236; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_237; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_238; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_239; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_240; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_241; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_242; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_243; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_244; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_245; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_246; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_247; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_248; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_249; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_250; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_251; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_252; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_253; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_254; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_255; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_256; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_257; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_258; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_259; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_260; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_261; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_262; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_263; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_264; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_265; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_266; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_267; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_268; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_269; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_270; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_271; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_272; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_273; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_274; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_275; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_276; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_277; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_278; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_279; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_280; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_281; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_282; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_283; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_284; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_285; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_286; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_287; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_288; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_289; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_290; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_291; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_292; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_293; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_294; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_295; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_296; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_297; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_298; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_299; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_300; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_301; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_302; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_303; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_304; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_305; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_306; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_307; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_308; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_309; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_310; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_311; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_312; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_313; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_314; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_315; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_316; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_317; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_318; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_319; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_320; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_321; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_322; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_323; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_324; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_325; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_326; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_327; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_328; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_329; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_330; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_331; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_332; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_333; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_334; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_335; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_336; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_337; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_338; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_339; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_340; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_341; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_342; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_343; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_344; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_345; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_346; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_347; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_348; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_349; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_350; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_351; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_352; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_353; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_354; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_355; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_356; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_357; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_358; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_359; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_360; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_361; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_362; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_363; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_364; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_365; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_366; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_367; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_368; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_369; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_370; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_371; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_372; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_373; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_374; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_375; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_376; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_377; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_378; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_379; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_380; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_381; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_382; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_383; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_384; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_385; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_386; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_387; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_388; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_389; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_390; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_391; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_392; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_393; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_394; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_395; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_396; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_397; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_398; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_399; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_400; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_401; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_402; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_403; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_404; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_405; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_406; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_407; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_408; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_409; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_410; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_411; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_412; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_413; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_414; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_415; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_416; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_417; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_418; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_419; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_420; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_421; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_422; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_423; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_424; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_425; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_426; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_427; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_428; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_429; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_430; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_431; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_432; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_433; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_434; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_435; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_436; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_437; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_438; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_439; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_440; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_441; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_442; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_443; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_444; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_445; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_446; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_447; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_448; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_449; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_450; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_451; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_452; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_453; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_454; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_455; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_456; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_457; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_458; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_459; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_460; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_461; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_462; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_463; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_464; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_465; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_466; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_467; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_468; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_469; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_470; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_471; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_472; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_473; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_474; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_475; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_476; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_477; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_478; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_479; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_480; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_481; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_482; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_483; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_484; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_485; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_486; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_487; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_488; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_489; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_490; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_491; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_492; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_493; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_494; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_495; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_496; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_497; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_498; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_499; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_500; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_501; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_502; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_503; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_504; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_505; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_506; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_507; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_508; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_509; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_510; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_data_511; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_0; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_1; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_2; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_3; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_4; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_5; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_6; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_7; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_8; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_9; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_10; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_11; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_12; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_13; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_14; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_header_15; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 491:23]
  wire [15:0] pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_out_next_config_id; // @[executor.scala 491:23]
  wire  pipe3_io_pipe_phv_out_is_valid_processor; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_4; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_5; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_args_in_6; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_0; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_1; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_2; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_in_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_offset_in_3; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_0; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_1; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_2; // @[executor.scala 491:23]
  wire [7:0] pipe3_io_length_in_3; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_0; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_1; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_2; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_vliw_out_3; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_0; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_1; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_2; // @[executor.scala 491:23]
  wire [31:0] pipe3_io_field_out_3; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_0; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_1; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_2; // @[executor.scala 491:23]
  wire [3:0] pipe3_io_mask_out_3; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_0; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_1; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_2; // @[executor.scala 491:23]
  wire [1:0] pipe3_io_bias_out_3; // @[executor.scala 491:23]
  wire  pipe4_clock; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_0; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_1; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_2; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_3; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_4; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_5; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_6; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_7; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_8; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_9; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_10; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_11; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_12; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_13; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_14; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_16; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_17; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_18; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_19; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_20; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_21; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_22; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_23; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_24; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_25; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_26; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_27; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_28; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_29; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_30; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_31; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_32; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_33; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_34; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_35; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_36; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_37; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_38; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_39; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_40; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_41; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_42; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_43; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_44; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_45; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_46; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_47; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_48; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_49; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_50; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_51; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_52; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_53; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_54; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_55; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_56; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_57; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_58; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_59; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_60; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_61; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_62; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_63; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_64; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_65; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_66; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_67; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_68; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_69; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_70; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_71; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_72; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_73; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_74; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_75; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_76; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_77; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_78; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_79; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_80; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_81; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_82; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_83; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_84; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_85; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_86; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_87; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_88; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_89; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_90; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_91; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_92; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_93; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_94; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_95; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_96; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_97; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_98; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_99; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_100; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_101; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_102; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_103; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_104; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_105; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_106; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_107; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_108; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_109; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_110; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_111; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_112; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_113; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_114; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_115; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_116; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_117; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_118; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_119; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_120; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_121; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_122; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_123; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_124; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_125; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_126; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_127; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_128; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_129; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_130; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_131; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_132; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_133; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_134; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_135; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_136; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_137; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_138; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_139; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_140; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_141; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_142; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_143; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_144; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_145; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_146; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_147; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_148; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_149; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_150; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_151; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_152; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_153; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_154; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_155; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_156; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_157; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_158; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_159; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_160; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_161; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_162; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_163; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_164; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_165; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_166; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_167; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_168; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_169; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_170; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_171; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_172; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_173; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_174; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_175; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_176; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_177; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_178; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_179; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_180; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_181; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_182; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_183; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_184; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_185; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_186; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_187; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_188; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_189; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_190; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_191; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_192; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_193; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_194; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_195; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_196; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_197; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_198; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_199; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_200; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_201; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_202; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_203; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_204; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_205; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_206; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_207; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_208; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_209; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_210; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_211; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_212; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_213; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_214; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_215; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_216; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_217; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_218; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_219; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_220; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_221; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_222; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_223; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_224; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_225; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_226; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_227; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_228; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_229; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_230; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_231; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_232; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_233; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_234; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_235; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_236; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_237; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_238; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_239; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_240; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_241; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_242; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_243; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_244; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_245; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_246; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_247; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_248; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_249; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_250; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_251; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_252; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_253; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_254; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_255; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_256; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_257; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_258; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_259; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_260; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_261; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_262; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_263; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_264; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_265; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_266; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_267; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_268; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_269; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_270; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_271; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_272; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_273; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_274; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_275; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_276; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_277; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_278; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_279; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_280; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_281; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_282; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_283; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_284; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_285; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_286; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_287; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_288; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_289; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_290; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_291; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_292; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_293; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_294; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_295; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_296; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_297; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_298; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_299; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_300; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_301; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_302; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_303; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_304; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_305; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_306; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_307; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_308; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_309; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_310; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_311; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_312; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_313; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_314; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_315; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_316; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_317; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_318; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_319; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_320; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_321; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_322; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_323; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_324; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_325; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_326; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_327; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_328; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_329; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_330; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_331; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_332; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_333; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_334; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_335; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_336; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_337; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_338; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_339; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_340; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_341; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_342; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_343; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_344; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_345; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_346; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_347; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_348; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_349; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_350; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_351; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_352; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_353; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_354; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_355; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_356; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_357; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_358; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_359; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_360; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_361; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_362; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_363; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_364; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_365; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_366; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_367; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_368; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_369; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_370; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_371; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_372; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_373; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_374; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_375; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_376; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_377; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_378; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_379; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_380; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_381; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_382; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_383; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_384; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_385; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_386; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_387; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_388; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_389; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_390; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_391; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_392; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_393; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_394; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_395; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_396; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_397; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_398; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_399; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_400; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_401; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_402; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_403; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_404; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_405; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_406; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_407; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_408; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_409; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_410; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_411; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_412; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_413; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_414; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_415; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_416; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_417; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_418; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_419; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_420; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_421; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_422; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_423; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_424; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_425; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_426; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_427; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_428; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_429; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_430; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_431; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_432; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_433; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_434; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_435; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_436; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_437; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_438; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_439; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_440; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_441; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_442; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_443; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_444; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_445; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_446; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_447; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_448; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_449; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_450; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_451; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_452; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_453; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_454; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_455; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_456; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_457; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_458; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_459; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_460; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_461; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_462; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_463; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_464; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_465; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_466; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_467; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_468; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_469; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_470; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_471; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_472; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_473; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_474; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_475; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_476; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_477; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_478; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_479; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_480; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_481; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_482; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_483; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_484; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_485; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_486; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_487; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_488; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_489; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_490; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_491; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_492; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_493; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_494; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_495; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_496; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_497; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_498; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_499; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_500; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_501; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_502; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_503; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_504; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_505; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_506; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_507; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_508; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_509; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_510; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_data_511; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_0; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_1; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_2; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_3; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_4; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_5; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_6; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_7; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_8; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_9; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_10; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_11; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_12; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_13; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_14; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_header_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_state; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_in_parse_current_offset; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_in_parse_transition_field; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_pipe_phv_in_next_processor_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_in_next_config_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_in_is_valid_processor; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_0; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_1; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_2; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_3; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_4; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_5; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_6; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_7; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_8; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_9; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_10; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_11; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_12; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_13; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_14; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_16; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_17; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_18; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_19; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_20; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_21; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_22; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_23; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_24; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_25; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_26; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_27; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_28; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_29; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_30; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_31; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_32; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_33; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_34; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_35; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_36; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_37; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_38; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_39; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_40; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_41; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_42; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_43; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_44; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_45; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_46; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_47; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_48; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_49; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_50; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_51; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_52; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_53; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_54; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_55; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_56; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_57; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_58; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_59; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_60; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_61; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_62; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_63; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_64; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_65; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_66; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_67; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_68; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_69; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_70; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_71; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_72; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_73; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_74; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_75; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_76; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_77; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_78; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_79; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_80; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_81; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_82; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_83; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_84; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_85; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_86; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_87; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_88; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_89; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_90; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_91; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_92; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_93; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_94; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_95; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_96; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_97; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_98; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_99; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_100; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_101; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_102; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_103; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_104; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_105; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_106; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_107; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_108; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_109; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_110; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_111; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_112; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_113; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_114; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_115; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_116; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_117; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_118; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_119; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_120; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_121; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_122; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_123; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_124; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_125; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_126; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_127; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_128; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_129; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_130; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_131; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_132; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_133; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_134; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_135; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_136; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_137; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_138; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_139; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_140; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_141; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_142; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_143; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_144; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_145; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_146; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_147; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_148; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_149; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_150; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_151; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_152; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_153; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_154; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_155; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_156; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_157; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_158; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_159; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_160; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_161; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_162; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_163; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_164; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_165; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_166; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_167; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_168; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_169; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_170; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_171; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_172; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_173; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_174; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_175; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_176; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_177; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_178; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_179; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_180; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_181; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_182; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_183; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_184; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_185; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_186; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_187; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_188; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_189; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_190; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_191; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_192; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_193; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_194; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_195; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_196; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_197; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_198; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_199; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_200; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_201; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_202; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_203; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_204; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_205; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_206; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_207; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_208; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_209; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_210; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_211; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_212; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_213; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_214; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_215; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_216; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_217; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_218; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_219; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_220; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_221; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_222; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_223; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_224; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_225; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_226; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_227; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_228; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_229; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_230; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_231; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_232; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_233; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_234; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_235; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_236; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_237; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_238; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_239; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_240; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_241; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_242; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_243; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_244; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_245; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_246; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_247; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_248; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_249; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_250; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_251; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_252; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_253; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_254; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_255; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_256; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_257; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_258; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_259; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_260; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_261; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_262; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_263; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_264; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_265; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_266; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_267; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_268; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_269; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_270; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_271; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_272; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_273; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_274; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_275; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_276; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_277; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_278; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_279; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_280; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_281; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_282; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_283; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_284; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_285; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_286; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_287; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_288; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_289; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_290; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_291; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_292; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_293; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_294; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_295; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_296; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_297; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_298; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_299; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_300; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_301; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_302; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_303; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_304; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_305; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_306; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_307; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_308; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_309; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_310; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_311; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_312; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_313; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_314; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_315; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_316; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_317; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_318; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_319; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_320; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_321; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_322; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_323; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_324; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_325; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_326; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_327; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_328; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_329; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_330; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_331; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_332; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_333; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_334; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_335; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_336; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_337; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_338; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_339; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_340; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_341; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_342; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_343; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_344; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_345; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_346; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_347; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_348; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_349; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_350; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_351; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_352; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_353; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_354; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_355; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_356; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_357; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_358; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_359; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_360; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_361; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_362; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_363; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_364; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_365; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_366; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_367; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_368; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_369; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_370; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_371; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_372; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_373; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_374; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_375; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_376; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_377; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_378; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_379; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_380; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_381; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_382; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_383; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_384; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_385; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_386; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_387; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_388; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_389; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_390; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_391; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_392; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_393; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_394; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_395; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_396; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_397; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_398; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_399; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_400; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_401; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_402; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_403; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_404; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_405; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_406; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_407; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_408; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_409; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_410; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_411; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_412; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_413; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_414; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_415; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_416; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_417; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_418; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_419; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_420; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_421; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_422; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_423; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_424; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_425; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_426; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_427; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_428; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_429; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_430; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_431; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_432; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_433; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_434; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_435; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_436; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_437; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_438; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_439; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_440; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_441; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_442; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_443; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_444; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_445; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_446; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_447; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_448; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_449; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_450; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_451; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_452; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_453; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_454; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_455; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_456; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_457; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_458; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_459; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_460; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_461; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_462; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_463; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_464; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_465; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_466; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_467; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_468; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_469; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_470; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_471; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_472; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_473; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_474; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_475; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_476; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_477; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_478; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_479; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_480; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_481; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_482; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_483; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_484; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_485; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_486; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_487; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_488; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_489; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_490; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_491; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_492; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_493; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_494; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_495; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_496; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_497; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_498; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_499; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_500; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_501; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_502; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_503; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_504; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_505; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_506; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_507; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_508; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_509; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_510; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_data_511; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_0; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_1; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_2; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_3; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_4; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_5; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_6; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_7; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_8; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_9; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_10; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_11; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_12; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_13; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_14; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_header_15; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 492:23]
  wire [7:0] pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 492:23]
  wire [15:0] pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_out_next_config_id; // @[executor.scala 492:23]
  wire  pipe4_io_pipe_phv_out_is_valid_processor; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_in_3; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_in_3; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_0; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_1; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_2; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_in_3; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_0; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_1; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_2; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_in_3; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_vliw_out_3; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_0; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_1; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_2; // @[executor.scala 492:23]
  wire [31:0] pipe4_io_field_out_3; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_0; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_1; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_2; // @[executor.scala 492:23]
  wire [3:0] pipe4_io_mask_out_3; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_0; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_1; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_2; // @[executor.scala 492:23]
  wire [1:0] pipe4_io_bias_out_3; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_0; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_1; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_2; // @[executor.scala 492:23]
  wire [5:0] pipe4_io_dst_offset_out_3; // @[executor.scala 492:23]
  wire  pipe5_clock; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_0; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_1; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_2; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_3; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_4; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_5; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_6; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_7; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_8; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_9; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_10; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_11; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_12; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_13; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_14; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_16; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_17; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_18; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_19; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_20; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_21; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_22; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_23; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_24; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_25; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_26; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_27; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_28; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_29; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_30; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_31; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_32; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_33; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_34; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_35; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_36; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_37; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_38; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_39; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_40; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_41; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_42; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_43; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_44; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_45; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_46; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_47; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_48; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_49; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_50; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_51; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_52; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_53; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_54; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_55; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_56; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_57; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_58; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_59; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_60; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_61; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_62; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_63; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_64; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_65; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_66; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_67; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_68; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_69; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_70; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_71; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_72; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_73; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_74; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_75; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_76; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_77; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_78; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_79; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_80; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_81; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_82; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_83; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_84; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_85; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_86; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_87; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_88; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_89; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_90; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_91; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_92; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_93; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_94; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_95; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_96; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_97; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_98; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_99; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_100; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_101; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_102; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_103; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_104; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_105; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_106; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_107; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_108; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_109; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_110; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_111; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_112; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_113; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_114; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_115; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_116; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_117; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_118; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_119; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_120; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_121; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_122; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_123; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_124; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_125; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_126; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_127; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_128; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_129; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_130; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_131; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_132; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_133; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_134; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_135; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_136; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_137; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_138; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_139; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_140; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_141; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_142; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_143; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_144; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_145; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_146; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_147; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_148; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_149; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_150; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_151; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_152; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_153; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_154; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_155; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_156; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_157; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_158; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_159; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_160; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_161; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_162; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_163; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_164; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_165; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_166; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_167; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_168; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_169; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_170; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_171; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_172; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_173; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_174; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_175; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_176; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_177; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_178; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_179; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_180; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_181; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_182; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_183; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_184; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_185; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_186; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_187; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_188; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_189; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_190; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_191; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_192; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_193; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_194; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_195; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_196; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_197; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_198; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_199; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_200; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_201; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_202; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_203; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_204; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_205; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_206; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_207; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_208; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_209; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_210; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_211; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_212; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_213; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_214; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_215; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_216; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_217; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_218; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_219; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_220; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_221; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_222; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_223; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_224; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_225; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_226; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_227; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_228; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_229; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_230; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_231; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_232; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_233; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_234; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_235; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_236; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_237; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_238; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_239; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_240; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_241; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_242; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_243; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_244; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_245; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_246; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_247; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_248; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_249; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_250; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_251; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_252; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_253; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_254; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_255; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_256; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_257; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_258; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_259; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_260; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_261; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_262; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_263; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_264; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_265; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_266; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_267; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_268; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_269; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_270; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_271; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_272; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_273; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_274; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_275; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_276; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_277; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_278; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_279; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_280; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_281; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_282; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_283; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_284; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_285; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_286; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_287; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_288; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_289; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_290; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_291; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_292; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_293; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_294; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_295; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_296; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_297; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_298; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_299; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_300; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_301; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_302; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_303; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_304; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_305; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_306; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_307; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_308; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_309; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_310; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_311; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_312; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_313; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_314; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_315; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_316; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_317; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_318; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_319; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_320; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_321; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_322; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_323; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_324; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_325; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_326; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_327; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_328; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_329; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_330; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_331; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_332; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_333; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_334; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_335; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_336; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_337; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_338; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_339; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_340; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_341; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_342; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_343; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_344; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_345; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_346; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_347; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_348; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_349; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_350; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_351; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_352; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_353; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_354; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_355; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_356; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_357; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_358; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_359; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_360; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_361; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_362; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_363; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_364; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_365; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_366; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_367; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_368; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_369; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_370; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_371; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_372; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_373; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_374; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_375; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_376; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_377; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_378; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_379; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_380; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_381; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_382; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_383; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_384; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_385; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_386; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_387; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_388; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_389; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_390; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_391; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_392; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_393; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_394; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_395; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_396; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_397; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_398; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_399; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_400; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_401; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_402; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_403; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_404; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_405; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_406; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_407; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_408; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_409; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_410; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_411; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_412; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_413; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_414; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_415; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_416; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_417; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_418; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_419; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_420; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_421; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_422; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_423; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_424; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_425; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_426; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_427; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_428; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_429; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_430; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_431; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_432; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_433; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_434; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_435; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_436; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_437; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_438; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_439; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_440; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_441; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_442; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_443; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_444; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_445; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_446; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_447; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_448; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_449; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_450; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_451; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_452; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_453; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_454; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_455; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_456; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_457; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_458; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_459; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_460; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_461; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_462; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_463; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_464; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_465; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_466; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_467; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_468; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_469; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_470; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_471; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_472; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_473; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_474; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_475; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_476; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_477; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_478; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_479; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_480; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_481; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_482; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_483; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_484; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_485; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_486; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_487; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_488; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_489; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_490; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_491; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_492; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_493; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_494; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_495; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_496; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_497; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_498; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_499; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_500; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_501; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_502; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_503; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_504; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_505; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_506; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_507; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_508; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_509; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_510; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_data_511; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_0; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_1; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_2; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_3; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_4; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_5; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_6; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_7; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_8; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_9; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_10; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_11; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_12; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_13; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_14; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_header_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_state; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_in_parse_current_offset; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_in_parse_transition_field; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_pipe_phv_in_next_processor_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_in_next_config_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_in_is_valid_processor; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_0; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_1; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_2; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_3; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_4; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_5; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_6; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_7; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_8; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_9; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_10; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_11; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_12; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_13; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_14; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_16; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_17; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_18; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_19; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_20; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_21; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_22; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_23; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_24; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_25; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_26; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_27; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_28; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_29; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_30; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_31; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_32; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_33; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_34; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_35; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_36; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_37; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_38; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_39; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_40; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_41; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_42; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_43; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_44; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_45; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_46; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_47; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_48; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_49; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_50; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_51; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_52; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_53; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_54; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_55; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_56; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_57; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_58; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_59; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_60; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_61; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_62; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_63; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_64; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_65; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_66; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_67; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_68; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_69; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_70; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_71; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_72; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_73; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_74; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_75; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_76; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_77; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_78; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_79; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_80; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_81; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_82; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_83; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_84; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_85; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_86; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_87; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_88; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_89; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_90; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_91; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_92; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_93; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_94; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_95; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_96; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_97; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_98; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_99; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_100; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_101; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_102; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_103; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_104; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_105; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_106; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_107; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_108; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_109; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_110; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_111; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_112; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_113; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_114; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_115; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_116; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_117; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_118; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_119; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_120; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_121; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_122; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_123; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_124; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_125; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_126; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_127; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_128; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_129; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_130; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_131; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_132; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_133; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_134; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_135; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_136; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_137; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_138; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_139; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_140; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_141; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_142; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_143; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_144; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_145; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_146; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_147; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_148; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_149; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_150; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_151; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_152; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_153; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_154; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_155; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_156; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_157; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_158; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_159; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_160; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_161; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_162; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_163; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_164; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_165; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_166; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_167; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_168; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_169; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_170; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_171; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_172; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_173; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_174; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_175; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_176; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_177; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_178; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_179; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_180; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_181; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_182; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_183; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_184; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_185; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_186; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_187; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_188; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_189; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_190; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_191; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_192; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_193; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_194; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_195; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_196; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_197; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_198; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_199; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_200; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_201; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_202; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_203; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_204; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_205; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_206; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_207; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_208; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_209; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_210; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_211; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_212; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_213; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_214; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_215; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_216; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_217; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_218; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_219; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_220; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_221; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_222; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_223; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_224; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_225; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_226; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_227; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_228; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_229; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_230; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_231; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_232; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_233; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_234; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_235; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_236; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_237; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_238; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_239; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_240; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_241; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_242; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_243; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_244; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_245; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_246; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_247; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_248; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_249; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_250; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_251; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_252; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_253; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_254; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_255; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_256; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_257; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_258; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_259; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_260; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_261; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_262; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_263; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_264; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_265; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_266; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_267; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_268; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_269; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_270; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_271; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_272; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_273; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_274; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_275; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_276; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_277; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_278; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_279; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_280; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_281; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_282; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_283; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_284; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_285; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_286; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_287; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_288; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_289; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_290; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_291; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_292; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_293; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_294; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_295; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_296; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_297; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_298; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_299; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_300; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_301; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_302; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_303; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_304; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_305; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_306; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_307; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_308; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_309; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_310; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_311; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_312; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_313; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_314; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_315; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_316; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_317; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_318; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_319; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_320; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_321; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_322; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_323; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_324; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_325; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_326; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_327; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_328; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_329; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_330; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_331; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_332; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_333; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_334; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_335; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_336; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_337; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_338; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_339; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_340; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_341; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_342; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_343; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_344; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_345; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_346; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_347; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_348; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_349; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_350; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_351; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_352; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_353; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_354; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_355; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_356; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_357; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_358; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_359; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_360; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_361; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_362; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_363; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_364; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_365; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_366; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_367; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_368; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_369; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_370; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_371; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_372; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_373; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_374; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_375; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_376; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_377; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_378; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_379; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_380; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_381; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_382; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_383; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_384; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_385; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_386; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_387; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_388; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_389; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_390; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_391; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_392; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_393; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_394; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_395; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_396; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_397; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_398; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_399; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_400; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_401; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_402; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_403; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_404; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_405; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_406; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_407; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_408; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_409; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_410; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_411; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_412; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_413; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_414; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_415; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_416; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_417; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_418; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_419; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_420; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_421; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_422; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_423; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_424; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_425; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_426; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_427; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_428; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_429; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_430; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_431; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_432; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_433; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_434; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_435; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_436; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_437; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_438; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_439; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_440; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_441; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_442; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_443; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_444; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_445; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_446; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_447; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_448; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_449; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_450; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_451; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_452; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_453; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_454; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_455; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_456; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_457; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_458; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_459; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_460; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_461; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_462; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_463; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_464; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_465; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_466; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_467; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_468; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_469; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_470; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_471; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_472; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_473; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_474; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_475; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_476; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_477; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_478; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_479; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_480; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_481; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_482; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_483; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_484; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_485; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_486; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_487; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_488; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_489; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_490; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_491; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_492; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_493; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_494; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_495; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_496; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_497; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_498; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_499; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_500; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_501; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_502; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_503; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_504; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_505; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_506; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_507; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_508; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_509; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_510; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_data_511; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_0; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_1; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_2; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_3; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_4; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_5; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_6; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_7; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_8; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_9; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_10; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_11; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_12; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_13; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_14; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_header_15; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 493:23]
  wire [7:0] pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 493:23]
  wire [15:0] pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_out_next_config_id; // @[executor.scala 493:23]
  wire  pipe5_io_pipe_phv_out_is_valid_processor; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_in_3; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_in_3; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_0; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_1; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_2; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_in_3; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_0; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_1; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_2; // @[executor.scala 493:23]
  wire [1:0] pipe5_io_bias_in_3; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_0; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_1; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_2; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_in_3; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_vliw_out_3; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_0; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_1; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_2; // @[executor.scala 493:23]
  wire [31:0] pipe5_io_field_out_3; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_0; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_1; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_2; // @[executor.scala 493:23]
  wire [3:0] pipe5_io_mask_out_3; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_0; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_1; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_2; // @[executor.scala 493:23]
  wire [5:0] pipe5_io_dst_offset_out_3; // @[executor.scala 493:23]
  wire  pipe6_clock; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_0; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_1; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_2; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_3; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_4; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_5; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_6; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_7; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_8; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_9; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_10; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_11; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_12; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_13; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_14; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_16; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_17; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_18; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_19; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_20; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_21; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_22; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_23; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_24; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_25; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_26; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_27; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_28; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_29; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_30; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_31; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_32; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_33; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_34; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_35; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_36; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_37; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_38; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_39; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_40; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_41; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_42; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_43; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_44; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_45; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_46; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_47; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_48; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_49; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_50; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_51; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_52; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_53; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_54; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_55; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_56; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_57; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_58; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_59; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_60; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_61; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_62; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_63; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_64; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_65; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_66; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_67; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_68; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_69; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_70; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_71; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_72; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_73; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_74; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_75; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_76; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_77; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_78; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_79; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_80; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_81; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_82; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_83; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_84; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_85; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_86; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_87; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_88; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_89; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_90; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_91; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_92; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_93; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_94; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_95; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_96; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_97; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_98; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_99; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_100; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_101; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_102; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_103; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_104; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_105; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_106; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_107; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_108; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_109; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_110; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_111; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_112; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_113; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_114; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_115; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_116; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_117; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_118; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_119; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_120; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_121; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_122; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_123; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_124; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_125; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_126; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_127; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_128; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_129; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_130; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_131; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_132; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_133; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_134; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_135; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_136; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_137; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_138; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_139; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_140; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_141; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_142; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_143; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_144; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_145; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_146; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_147; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_148; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_149; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_150; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_151; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_152; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_153; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_154; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_155; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_156; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_157; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_158; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_159; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_160; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_161; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_162; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_163; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_164; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_165; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_166; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_167; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_168; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_169; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_170; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_171; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_172; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_173; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_174; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_175; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_176; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_177; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_178; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_179; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_180; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_181; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_182; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_183; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_184; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_185; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_186; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_187; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_188; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_189; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_190; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_191; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_192; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_193; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_194; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_195; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_196; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_197; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_198; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_199; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_200; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_201; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_202; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_203; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_204; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_205; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_206; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_207; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_208; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_209; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_210; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_211; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_212; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_213; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_214; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_215; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_216; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_217; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_218; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_219; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_220; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_221; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_222; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_223; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_224; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_225; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_226; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_227; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_228; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_229; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_230; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_231; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_232; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_233; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_234; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_235; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_236; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_237; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_238; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_239; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_240; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_241; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_242; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_243; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_244; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_245; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_246; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_247; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_248; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_249; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_250; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_251; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_252; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_253; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_254; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_255; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_256; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_257; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_258; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_259; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_260; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_261; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_262; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_263; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_264; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_265; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_266; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_267; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_268; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_269; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_270; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_271; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_272; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_273; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_274; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_275; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_276; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_277; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_278; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_279; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_280; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_281; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_282; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_283; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_284; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_285; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_286; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_287; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_288; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_289; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_290; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_291; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_292; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_293; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_294; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_295; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_296; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_297; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_298; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_299; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_300; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_301; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_302; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_303; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_304; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_305; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_306; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_307; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_308; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_309; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_310; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_311; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_312; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_313; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_314; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_315; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_316; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_317; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_318; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_319; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_320; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_321; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_322; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_323; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_324; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_325; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_326; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_327; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_328; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_329; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_330; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_331; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_332; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_333; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_334; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_335; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_336; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_337; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_338; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_339; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_340; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_341; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_342; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_343; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_344; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_345; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_346; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_347; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_348; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_349; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_350; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_351; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_352; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_353; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_354; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_355; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_356; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_357; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_358; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_359; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_360; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_361; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_362; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_363; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_364; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_365; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_366; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_367; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_368; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_369; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_370; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_371; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_372; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_373; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_374; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_375; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_376; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_377; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_378; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_379; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_380; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_381; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_382; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_383; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_384; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_385; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_386; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_387; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_388; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_389; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_390; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_391; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_392; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_393; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_394; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_395; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_396; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_397; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_398; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_399; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_400; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_401; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_402; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_403; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_404; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_405; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_406; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_407; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_408; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_409; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_410; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_411; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_412; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_413; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_414; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_415; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_416; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_417; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_418; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_419; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_420; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_421; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_422; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_423; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_424; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_425; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_426; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_427; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_428; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_429; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_430; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_431; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_432; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_433; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_434; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_435; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_436; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_437; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_438; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_439; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_440; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_441; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_442; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_443; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_444; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_445; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_446; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_447; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_448; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_449; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_450; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_451; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_452; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_453; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_454; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_455; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_456; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_457; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_458; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_459; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_460; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_461; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_462; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_463; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_464; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_465; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_466; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_467; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_468; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_469; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_470; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_471; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_472; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_473; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_474; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_475; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_476; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_477; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_478; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_479; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_480; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_481; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_482; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_483; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_484; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_485; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_486; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_487; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_488; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_489; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_490; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_491; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_492; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_493; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_494; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_495; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_496; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_497; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_498; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_499; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_500; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_501; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_502; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_503; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_504; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_505; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_506; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_507; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_508; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_509; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_510; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_data_511; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_0; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_1; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_2; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_3; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_4; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_5; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_6; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_7; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_8; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_9; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_10; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_11; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_12; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_13; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_14; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_header_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_state; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_in_parse_current_offset; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_in_parse_transition_field; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_pipe_phv_in_next_processor_id; // @[executor.scala 494:23]
  wire  pipe6_io_pipe_phv_in_next_config_id; // @[executor.scala 494:23]
  wire  pipe6_io_pipe_phv_in_is_valid_processor; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_0; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_1; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_2; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_3; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_4; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_5; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_6; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_7; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_8; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_9; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_10; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_11; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_12; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_13; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_14; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_16; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_17; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_18; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_19; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_20; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_21; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_22; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_23; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_24; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_25; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_26; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_27; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_28; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_29; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_30; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_31; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_32; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_33; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_34; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_35; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_36; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_37; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_38; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_39; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_40; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_41; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_42; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_43; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_44; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_45; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_46; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_47; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_48; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_49; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_50; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_51; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_52; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_53; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_54; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_55; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_56; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_57; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_58; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_59; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_60; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_61; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_62; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_63; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_64; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_65; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_66; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_67; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_68; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_69; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_70; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_71; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_72; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_73; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_74; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_75; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_76; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_77; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_78; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_79; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_80; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_81; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_82; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_83; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_84; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_85; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_86; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_87; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_88; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_89; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_90; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_91; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_92; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_93; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_94; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_95; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_96; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_97; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_98; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_99; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_100; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_101; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_102; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_103; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_104; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_105; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_106; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_107; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_108; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_109; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_110; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_111; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_112; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_113; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_114; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_115; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_116; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_117; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_118; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_119; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_120; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_121; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_122; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_123; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_124; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_125; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_126; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_127; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_128; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_129; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_130; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_131; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_132; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_133; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_134; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_135; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_136; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_137; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_138; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_139; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_140; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_141; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_142; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_143; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_144; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_145; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_146; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_147; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_148; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_149; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_150; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_151; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_152; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_153; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_154; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_155; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_156; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_157; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_158; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_159; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_160; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_161; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_162; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_163; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_164; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_165; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_166; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_167; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_168; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_169; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_170; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_171; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_172; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_173; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_174; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_175; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_176; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_177; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_178; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_179; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_180; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_181; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_182; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_183; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_184; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_185; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_186; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_187; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_188; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_189; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_190; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_191; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_192; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_193; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_194; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_195; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_196; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_197; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_198; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_199; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_200; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_201; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_202; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_203; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_204; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_205; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_206; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_207; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_208; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_209; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_210; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_211; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_212; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_213; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_214; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_215; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_216; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_217; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_218; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_219; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_220; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_221; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_222; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_223; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_224; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_225; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_226; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_227; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_228; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_229; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_230; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_231; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_232; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_233; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_234; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_235; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_236; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_237; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_238; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_239; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_240; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_241; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_242; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_243; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_244; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_245; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_246; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_247; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_248; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_249; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_250; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_251; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_252; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_253; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_254; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_255; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_256; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_257; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_258; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_259; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_260; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_261; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_262; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_263; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_264; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_265; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_266; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_267; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_268; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_269; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_270; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_271; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_272; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_273; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_274; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_275; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_276; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_277; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_278; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_279; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_280; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_281; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_282; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_283; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_284; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_285; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_286; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_287; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_288; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_289; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_290; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_291; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_292; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_293; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_294; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_295; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_296; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_297; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_298; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_299; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_300; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_301; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_302; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_303; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_304; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_305; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_306; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_307; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_308; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_309; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_310; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_311; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_312; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_313; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_314; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_315; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_316; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_317; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_318; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_319; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_320; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_321; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_322; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_323; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_324; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_325; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_326; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_327; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_328; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_329; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_330; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_331; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_332; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_333; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_334; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_335; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_336; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_337; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_338; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_339; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_340; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_341; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_342; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_343; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_344; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_345; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_346; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_347; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_348; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_349; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_350; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_351; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_352; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_353; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_354; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_355; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_356; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_357; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_358; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_359; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_360; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_361; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_362; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_363; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_364; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_365; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_366; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_367; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_368; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_369; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_370; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_371; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_372; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_373; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_374; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_375; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_376; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_377; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_378; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_379; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_380; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_381; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_382; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_383; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_384; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_385; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_386; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_387; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_388; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_389; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_390; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_391; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_392; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_393; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_394; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_395; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_396; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_397; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_398; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_399; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_400; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_401; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_402; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_403; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_404; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_405; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_406; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_407; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_408; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_409; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_410; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_411; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_412; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_413; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_414; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_415; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_416; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_417; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_418; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_419; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_420; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_421; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_422; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_423; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_424; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_425; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_426; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_427; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_428; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_429; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_430; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_431; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_432; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_433; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_434; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_435; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_436; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_437; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_438; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_439; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_440; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_441; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_442; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_443; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_444; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_445; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_446; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_447; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_448; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_449; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_450; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_451; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_452; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_453; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_454; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_455; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_456; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_457; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_458; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_459; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_460; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_461; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_462; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_463; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_464; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_465; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_466; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_467; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_468; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_469; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_470; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_471; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_472; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_473; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_474; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_475; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_476; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_477; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_478; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_479; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_480; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_481; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_482; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_483; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_484; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_485; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_486; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_487; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_488; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_489; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_490; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_491; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_492; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_493; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_494; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_495; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_496; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_497; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_498; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_499; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_500; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_501; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_502; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_503; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_504; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_505; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_506; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_507; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_508; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_509; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_510; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_data_511; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_0; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_1; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_2; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_3; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_4; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_5; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_6; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_7; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_8; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_9; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_10; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_11; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_12; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_13; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_14; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_header_15; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 494:23]
  wire [7:0] pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 494:23]
  wire [15:0] pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 494:23]
  wire  pipe6_io_pipe_phv_out_next_config_id; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_0; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_1; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_2; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_vliw_in_3; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_0; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_1; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_2; // @[executor.scala 494:23]
  wire [31:0] pipe6_io_field_in_3; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_0; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_1; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_2; // @[executor.scala 494:23]
  wire [3:0] pipe6_io_mask_in_3; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_0; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_1; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_2; // @[executor.scala 494:23]
  wire [5:0] pipe6_io_dst_offset_in_3; // @[executor.scala 494:23]
  ActionReader pipe1 ( // @[executor.scala 489:23]
    .clock(pipe1_clock),
    .io_pipe_phv_in_data_0(pipe1_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe1_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe1_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe1_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe1_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe1_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe1_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe1_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe1_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe1_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe1_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe1_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe1_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe1_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe1_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe1_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe1_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe1_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe1_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe1_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe1_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe1_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe1_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe1_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe1_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe1_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe1_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe1_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe1_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe1_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe1_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe1_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe1_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe1_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe1_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe1_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe1_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe1_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe1_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe1_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe1_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe1_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe1_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe1_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe1_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe1_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe1_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe1_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe1_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe1_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe1_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe1_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe1_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe1_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe1_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe1_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe1_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe1_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe1_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe1_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe1_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe1_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe1_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe1_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe1_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe1_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe1_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe1_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe1_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe1_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe1_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe1_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe1_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe1_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe1_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe1_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe1_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe1_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe1_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe1_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe1_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe1_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe1_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe1_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe1_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe1_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe1_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe1_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe1_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe1_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe1_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe1_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe1_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe1_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe1_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe1_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe1_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe1_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe1_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe1_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe1_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe1_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe1_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe1_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe1_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe1_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe1_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe1_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe1_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe1_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe1_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe1_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe1_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe1_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe1_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe1_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe1_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe1_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe1_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe1_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe1_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe1_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe1_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe1_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe1_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe1_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe1_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe1_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe1_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe1_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe1_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe1_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe1_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe1_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe1_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe1_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe1_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe1_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe1_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe1_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe1_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe1_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe1_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe1_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe1_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe1_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe1_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe1_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe1_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe1_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe1_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe1_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe1_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe1_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe1_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe1_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe1_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe1_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe1_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe1_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe1_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe1_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe1_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe1_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe1_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe1_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe1_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe1_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe1_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe1_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe1_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe1_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe1_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe1_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe1_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe1_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe1_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe1_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe1_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe1_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe1_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe1_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe1_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe1_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe1_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe1_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe1_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe1_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe1_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe1_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe1_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe1_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe1_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe1_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe1_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe1_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe1_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe1_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe1_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe1_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe1_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe1_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe1_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe1_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe1_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe1_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe1_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe1_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe1_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe1_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe1_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe1_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe1_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe1_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe1_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe1_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe1_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe1_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe1_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe1_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe1_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe1_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe1_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe1_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe1_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe1_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe1_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe1_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe1_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe1_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe1_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe1_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe1_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe1_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe1_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe1_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe1_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe1_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe1_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe1_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe1_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe1_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe1_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe1_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe1_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe1_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe1_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe1_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe1_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe1_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe1_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe1_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe1_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe1_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe1_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe1_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe1_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe1_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe1_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe1_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe1_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe1_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe1_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe1_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe1_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe1_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe1_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe1_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe1_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe1_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe1_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe1_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe1_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe1_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe1_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe1_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe1_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe1_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe1_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe1_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe1_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe1_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe1_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe1_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe1_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe1_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe1_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe1_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe1_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe1_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe1_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe1_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe1_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe1_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe1_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe1_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe1_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe1_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe1_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe1_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe1_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe1_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe1_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe1_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe1_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe1_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe1_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe1_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe1_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe1_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe1_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe1_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe1_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe1_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe1_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe1_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe1_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe1_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe1_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe1_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe1_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe1_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe1_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe1_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe1_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe1_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe1_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe1_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe1_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe1_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe1_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe1_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe1_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe1_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe1_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe1_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe1_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe1_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe1_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe1_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe1_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe1_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe1_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe1_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe1_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe1_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe1_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe1_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe1_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe1_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe1_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe1_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe1_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe1_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe1_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe1_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe1_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe1_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe1_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe1_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe1_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe1_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe1_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe1_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe1_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe1_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe1_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe1_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe1_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe1_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe1_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe1_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe1_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe1_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe1_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe1_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe1_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe1_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe1_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe1_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe1_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe1_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe1_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe1_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe1_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe1_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe1_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe1_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe1_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe1_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe1_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe1_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe1_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe1_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe1_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe1_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe1_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe1_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe1_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe1_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe1_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe1_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe1_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe1_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe1_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe1_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe1_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe1_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe1_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe1_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe1_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe1_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe1_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe1_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe1_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe1_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe1_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe1_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe1_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe1_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe1_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe1_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe1_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe1_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe1_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe1_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe1_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe1_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe1_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe1_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe1_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe1_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe1_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe1_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe1_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe1_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe1_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe1_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe1_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe1_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe1_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe1_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe1_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe1_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe1_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe1_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe1_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe1_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe1_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe1_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe1_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe1_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe1_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe1_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe1_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe1_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe1_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe1_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe1_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe1_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe1_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe1_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe1_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe1_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe1_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe1_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe1_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe1_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe1_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe1_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe1_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe1_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe1_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe1_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe1_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe1_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe1_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe1_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe1_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe1_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe1_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe1_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe1_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe1_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe1_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe1_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe1_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe1_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe1_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe1_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe1_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe1_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe1_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe1_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe1_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe1_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe1_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe1_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe1_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe1_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe1_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe1_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe1_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe1_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe1_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe1_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe1_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe1_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe1_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe1_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe1_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe1_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe1_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe1_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe1_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe1_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe1_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe1_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe1_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe1_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe1_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe1_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe1_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe1_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe1_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe1_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe1_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe1_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe1_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe1_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe1_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe1_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe1_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe1_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe1_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe1_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe1_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe1_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe1_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe1_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe1_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe1_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe1_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe1_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe1_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe1_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe1_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe1_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe1_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe1_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe1_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe1_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe1_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe1_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe1_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe1_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe1_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe1_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe1_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe1_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe1_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe1_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe1_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe1_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe1_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe1_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe1_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe1_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe1_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe1_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe1_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe1_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe1_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe1_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe1_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe1_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe1_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe1_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe1_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe1_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe1_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe1_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe1_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe1_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe1_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe1_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe1_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe1_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe1_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe1_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe1_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe1_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe1_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe1_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe1_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe1_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe1_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe1_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe1_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe1_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe1_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe1_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe1_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe1_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe1_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe1_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe1_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe1_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe1_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe1_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe1_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe1_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe1_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe1_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe1_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe1_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe1_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe1_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe1_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe1_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe1_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe1_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe1_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe1_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe1_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe1_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe1_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe1_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe1_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe1_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe1_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe1_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe1_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe1_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe1_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe1_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe1_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe1_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe1_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe1_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe1_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe1_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe1_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe1_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe1_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe1_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe1_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe1_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe1_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe1_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe1_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe1_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe1_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe1_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe1_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe1_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe1_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe1_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe1_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe1_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe1_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe1_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe1_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe1_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe1_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe1_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe1_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe1_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe1_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe1_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe1_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe1_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe1_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe1_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe1_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe1_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe1_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe1_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe1_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe1_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe1_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe1_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe1_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe1_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe1_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe1_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe1_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe1_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe1_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe1_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe1_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe1_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe1_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe1_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe1_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe1_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe1_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe1_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe1_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe1_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe1_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe1_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe1_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe1_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe1_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe1_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe1_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe1_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe1_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe1_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe1_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe1_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe1_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe1_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe1_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe1_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe1_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe1_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe1_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe1_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe1_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe1_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe1_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe1_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe1_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe1_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe1_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe1_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe1_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe1_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe1_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe1_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe1_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe1_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe1_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe1_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe1_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe1_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe1_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe1_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe1_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe1_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe1_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe1_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe1_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe1_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe1_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe1_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe1_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe1_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe1_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe1_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe1_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe1_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe1_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe1_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe1_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe1_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe1_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe1_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe1_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe1_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe1_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe1_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe1_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe1_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe1_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe1_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe1_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe1_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe1_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe1_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe1_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe1_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe1_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe1_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe1_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe1_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe1_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe1_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe1_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe1_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe1_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe1_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe1_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe1_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe1_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe1_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe1_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe1_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe1_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe1_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe1_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe1_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe1_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe1_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe1_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe1_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe1_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe1_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe1_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe1_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe1_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe1_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe1_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe1_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe1_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe1_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe1_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe1_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe1_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe1_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe1_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe1_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe1_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe1_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe1_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe1_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe1_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe1_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe1_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe1_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe1_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe1_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe1_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe1_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe1_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe1_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe1_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe1_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe1_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe1_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe1_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe1_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe1_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe1_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe1_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe1_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe1_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe1_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe1_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe1_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe1_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe1_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe1_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe1_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe1_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe1_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe1_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe1_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe1_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe1_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe1_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe1_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe1_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe1_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe1_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe1_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe1_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe1_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe1_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe1_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe1_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe1_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe1_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe1_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe1_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe1_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe1_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe1_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe1_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe1_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe1_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe1_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe1_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe1_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe1_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe1_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe1_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe1_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe1_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe1_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe1_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe1_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe1_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe1_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe1_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe1_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe1_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe1_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe1_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe1_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe1_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe1_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe1_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe1_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe1_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe1_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe1_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe1_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe1_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe1_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe1_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe1_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe1_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe1_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe1_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe1_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe1_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe1_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe1_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe1_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe1_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe1_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe1_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe1_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe1_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe1_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe1_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe1_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe1_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe1_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe1_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe1_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe1_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe1_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe1_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe1_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe1_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe1_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe1_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe1_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe1_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe1_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe1_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe1_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe1_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe1_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe1_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe1_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe1_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe1_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe1_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe1_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe1_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe1_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe1_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe1_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe1_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe1_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe1_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe1_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe1_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe1_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe1_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe1_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe1_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe1_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe1_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe1_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe1_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe1_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe1_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe1_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe1_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe1_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe1_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe1_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe1_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe1_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe1_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe1_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe1_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe1_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe1_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe1_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe1_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe1_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe1_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe1_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe1_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe1_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe1_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe1_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe1_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe1_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe1_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe1_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe1_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe1_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe1_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe1_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe1_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe1_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe1_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe1_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe1_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe1_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe1_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe1_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe1_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe1_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe1_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe1_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe1_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe1_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe1_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe1_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe1_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe1_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe1_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe1_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe1_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe1_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe1_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe1_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe1_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe1_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe1_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe1_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe1_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe1_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe1_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe1_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe1_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe1_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe1_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe1_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe1_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe1_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe1_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe1_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe1_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe1_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe1_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe1_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe1_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe1_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe1_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe1_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe1_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe1_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe1_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe1_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe1_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe1_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe1_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe1_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe1_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe1_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe1_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe1_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe1_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe1_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe1_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe1_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe1_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe1_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe1_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe1_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe1_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe1_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe1_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe1_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe1_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe1_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe1_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe1_io_pipe_phv_out_is_valid_processor),
    .io_hit(pipe1_io_hit),
    .io_match_value(pipe1_io_match_value),
    .io_args_out_0(pipe1_io_args_out_0),
    .io_args_out_1(pipe1_io_args_out_1),
    .io_args_out_2(pipe1_io_args_out_2),
    .io_args_out_3(pipe1_io_args_out_3),
    .io_args_out_4(pipe1_io_args_out_4),
    .io_args_out_5(pipe1_io_args_out_5),
    .io_args_out_6(pipe1_io_args_out_6),
    .io_vliw_out_0(pipe1_io_vliw_out_0),
    .io_vliw_out_1(pipe1_io_vliw_out_1),
    .io_vliw_out_2(pipe1_io_vliw_out_2),
    .io_vliw_out_3(pipe1_io_vliw_out_3),
    .io_action_mod_en_0(pipe1_io_action_mod_en_0),
    .io_action_mod_en_1(pipe1_io_action_mod_en_1),
    .io_action_mod_addr(pipe1_io_action_mod_addr),
    .io_action_mod_data_0(pipe1_io_action_mod_data_0),
    .io_action_mod_data_1(pipe1_io_action_mod_data_1)
  );
  PrimitiveGetOffset pipe2 ( // @[executor.scala 490:23]
    .clock(pipe2_clock),
    .io_pipe_phv_in_data_0(pipe2_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe2_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe2_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe2_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe2_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe2_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe2_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe2_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe2_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe2_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe2_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe2_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe2_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe2_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe2_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe2_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe2_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe2_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe2_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe2_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe2_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe2_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe2_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe2_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe2_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe2_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe2_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe2_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe2_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe2_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe2_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe2_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe2_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe2_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe2_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe2_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe2_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe2_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe2_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe2_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe2_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe2_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe2_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe2_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe2_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe2_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe2_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe2_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe2_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe2_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe2_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe2_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe2_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe2_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe2_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe2_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe2_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe2_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe2_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe2_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe2_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe2_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe2_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe2_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe2_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe2_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe2_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe2_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe2_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe2_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe2_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe2_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe2_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe2_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe2_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe2_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe2_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe2_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe2_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe2_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe2_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe2_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe2_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe2_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe2_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe2_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe2_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe2_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe2_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe2_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe2_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe2_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe2_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe2_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe2_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe2_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe2_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe2_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe2_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe2_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe2_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe2_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe2_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe2_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe2_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe2_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe2_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe2_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe2_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe2_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe2_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe2_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe2_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe2_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe2_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe2_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe2_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe2_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe2_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe2_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe2_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe2_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe2_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe2_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe2_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe2_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe2_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe2_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe2_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe2_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe2_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe2_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe2_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe2_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe2_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe2_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe2_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe2_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe2_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe2_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe2_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe2_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe2_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe2_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe2_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe2_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe2_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe2_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe2_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe2_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe2_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe2_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe2_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe2_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe2_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe2_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe2_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe2_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe2_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe2_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe2_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe2_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe2_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe2_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe2_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe2_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe2_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe2_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe2_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe2_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe2_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe2_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe2_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe2_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe2_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe2_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe2_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe2_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe2_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe2_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe2_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe2_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe2_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe2_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe2_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe2_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe2_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe2_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe2_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe2_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe2_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe2_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe2_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe2_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe2_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe2_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe2_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe2_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe2_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe2_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe2_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe2_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe2_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe2_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe2_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe2_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe2_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe2_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe2_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe2_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe2_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe2_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe2_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe2_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe2_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe2_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe2_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe2_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe2_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe2_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe2_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe2_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe2_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe2_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe2_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe2_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe2_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe2_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe2_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe2_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe2_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe2_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe2_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe2_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe2_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe2_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe2_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe2_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe2_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe2_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe2_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe2_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe2_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe2_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe2_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe2_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe2_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe2_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe2_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe2_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe2_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe2_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe2_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe2_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe2_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe2_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe2_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe2_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe2_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe2_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe2_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe2_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe2_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe2_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe2_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe2_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe2_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe2_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe2_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe2_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe2_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe2_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe2_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe2_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe2_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe2_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe2_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe2_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe2_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe2_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe2_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe2_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe2_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe2_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe2_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe2_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe2_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe2_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe2_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe2_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe2_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe2_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe2_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe2_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe2_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe2_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe2_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe2_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe2_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe2_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe2_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe2_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe2_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe2_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe2_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe2_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe2_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe2_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe2_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe2_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe2_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe2_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe2_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe2_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe2_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe2_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe2_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe2_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe2_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe2_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe2_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe2_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe2_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe2_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe2_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe2_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe2_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe2_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe2_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe2_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe2_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe2_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe2_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe2_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe2_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe2_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe2_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe2_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe2_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe2_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe2_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe2_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe2_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe2_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe2_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe2_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe2_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe2_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe2_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe2_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe2_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe2_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe2_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe2_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe2_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe2_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe2_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe2_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe2_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe2_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe2_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe2_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe2_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe2_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe2_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe2_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe2_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe2_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe2_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe2_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe2_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe2_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe2_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe2_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe2_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe2_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe2_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe2_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe2_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe2_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe2_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe2_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe2_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe2_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe2_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe2_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe2_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe2_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe2_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe2_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe2_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe2_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe2_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe2_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe2_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe2_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe2_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe2_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe2_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe2_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe2_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe2_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe2_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe2_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe2_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe2_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe2_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe2_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe2_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe2_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe2_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe2_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe2_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe2_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe2_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe2_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe2_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe2_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe2_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe2_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe2_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe2_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe2_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe2_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe2_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe2_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe2_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe2_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe2_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe2_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe2_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe2_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe2_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe2_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe2_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe2_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe2_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe2_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe2_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe2_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe2_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe2_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe2_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe2_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe2_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe2_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe2_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe2_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe2_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe2_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe2_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe2_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe2_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe2_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe2_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe2_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe2_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe2_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe2_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe2_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe2_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe2_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe2_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe2_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe2_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe2_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe2_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe2_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe2_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe2_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe2_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe2_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe2_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe2_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe2_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe2_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe2_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe2_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe2_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe2_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe2_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe2_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe2_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe2_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe2_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe2_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe2_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe2_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe2_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe2_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe2_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe2_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe2_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe2_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe2_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe2_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe2_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe2_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe2_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe2_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe2_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe2_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe2_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe2_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe2_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe2_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe2_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe2_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe2_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe2_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe2_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe2_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe2_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe2_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe2_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe2_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe2_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe2_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe2_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe2_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe2_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe2_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe2_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe2_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe2_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe2_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe2_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe2_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe2_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe2_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe2_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe2_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe2_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe2_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe2_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe2_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe2_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe2_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe2_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe2_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe2_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe2_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe2_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe2_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe2_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe2_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe2_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe2_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe2_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe2_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe2_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe2_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe2_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe2_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe2_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe2_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe2_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe2_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe2_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe2_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe2_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe2_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe2_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe2_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe2_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe2_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe2_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe2_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe2_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe2_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe2_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe2_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe2_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe2_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe2_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe2_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe2_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe2_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe2_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe2_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe2_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe2_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe2_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe2_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe2_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe2_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe2_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe2_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe2_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe2_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe2_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe2_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe2_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe2_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe2_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe2_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe2_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe2_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe2_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe2_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe2_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe2_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe2_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe2_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe2_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe2_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe2_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe2_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe2_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe2_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe2_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe2_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe2_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe2_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe2_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe2_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe2_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe2_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe2_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe2_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe2_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe2_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe2_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe2_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe2_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe2_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe2_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe2_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe2_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe2_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe2_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe2_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe2_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe2_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe2_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe2_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe2_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe2_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe2_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe2_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe2_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe2_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe2_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe2_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe2_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe2_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe2_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe2_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe2_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe2_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe2_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe2_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe2_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe2_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe2_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe2_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe2_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe2_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe2_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe2_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe2_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe2_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe2_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe2_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe2_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe2_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe2_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe2_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe2_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe2_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe2_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe2_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe2_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe2_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe2_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe2_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe2_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe2_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe2_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe2_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe2_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe2_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe2_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe2_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe2_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe2_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe2_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe2_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe2_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe2_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe2_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe2_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe2_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe2_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe2_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe2_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe2_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe2_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe2_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe2_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe2_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe2_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe2_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe2_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe2_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe2_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe2_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe2_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe2_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe2_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe2_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe2_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe2_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe2_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe2_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe2_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe2_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe2_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe2_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe2_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe2_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe2_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe2_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe2_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe2_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe2_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe2_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe2_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe2_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe2_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe2_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe2_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe2_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe2_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe2_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe2_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe2_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe2_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe2_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe2_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe2_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe2_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe2_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe2_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe2_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe2_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe2_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe2_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe2_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe2_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe2_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe2_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe2_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe2_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe2_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe2_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe2_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe2_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe2_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe2_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe2_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe2_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe2_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe2_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe2_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe2_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe2_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe2_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe2_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe2_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe2_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe2_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe2_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe2_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe2_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe2_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe2_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe2_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe2_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe2_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe2_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe2_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe2_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe2_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe2_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe2_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe2_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe2_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe2_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe2_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe2_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe2_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe2_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe2_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe2_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe2_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe2_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe2_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe2_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe2_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe2_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe2_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe2_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe2_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe2_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe2_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe2_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe2_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe2_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe2_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe2_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe2_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe2_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe2_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe2_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe2_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe2_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe2_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe2_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe2_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe2_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe2_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe2_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe2_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe2_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe2_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe2_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe2_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe2_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe2_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe2_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe2_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe2_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe2_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe2_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe2_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe2_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe2_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe2_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe2_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe2_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe2_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe2_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe2_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe2_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe2_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe2_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe2_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe2_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe2_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe2_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe2_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe2_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe2_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe2_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe2_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe2_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe2_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe2_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe2_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe2_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe2_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe2_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe2_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe2_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe2_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe2_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe2_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe2_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe2_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe2_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe2_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe2_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe2_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe2_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe2_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe2_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe2_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe2_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe2_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe2_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe2_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe2_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe2_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe2_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe2_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe2_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe2_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe2_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe2_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe2_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe2_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe2_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe2_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe2_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe2_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe2_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe2_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe2_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe2_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe2_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe2_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe2_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe2_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe2_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe2_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe2_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe2_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe2_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe2_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe2_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe2_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe2_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe2_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe2_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe2_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe2_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe2_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe2_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe2_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe2_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe2_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe2_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe2_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe2_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe2_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe2_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe2_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe2_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe2_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe2_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe2_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe2_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe2_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe2_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe2_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe2_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe2_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe2_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe2_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe2_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe2_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe2_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe2_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe2_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe2_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe2_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe2_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe2_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe2_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe2_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe2_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe2_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe2_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe2_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe2_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe2_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe2_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe2_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe2_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe2_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe2_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe2_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe2_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe2_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe2_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe2_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe2_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe2_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe2_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe2_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe2_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe2_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe2_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe2_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe2_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe2_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe2_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe2_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe2_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe2_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe2_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe2_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe2_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe2_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe2_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe2_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe2_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe2_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe2_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe2_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe2_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe2_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe2_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe2_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe2_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe2_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe2_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe2_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe2_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe2_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe2_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe2_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe2_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe2_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe2_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe2_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe2_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe2_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe2_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe2_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe2_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe2_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe2_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe2_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe2_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe2_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe2_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe2_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe2_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe2_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe2_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe2_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe2_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe2_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe2_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe2_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe2_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe2_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe2_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe2_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe2_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe2_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe2_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe2_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe2_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe2_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe2_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe2_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe2_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe2_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe2_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe2_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe2_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe2_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe2_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe2_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe2_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe2_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe2_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe2_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe2_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe2_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe2_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe2_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe2_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe2_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe2_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe2_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe2_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe2_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe2_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe2_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe2_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe2_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe2_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe2_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe2_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe2_io_args_in_0),
    .io_args_in_1(pipe2_io_args_in_1),
    .io_args_in_2(pipe2_io_args_in_2),
    .io_args_in_3(pipe2_io_args_in_3),
    .io_args_in_4(pipe2_io_args_in_4),
    .io_args_in_5(pipe2_io_args_in_5),
    .io_args_in_6(pipe2_io_args_in_6),
    .io_vliw_in_0(pipe2_io_vliw_in_0),
    .io_vliw_in_1(pipe2_io_vliw_in_1),
    .io_vliw_in_2(pipe2_io_vliw_in_2),
    .io_vliw_in_3(pipe2_io_vliw_in_3),
    .io_args_out_0(pipe2_io_args_out_0),
    .io_args_out_1(pipe2_io_args_out_1),
    .io_args_out_2(pipe2_io_args_out_2),
    .io_args_out_3(pipe2_io_args_out_3),
    .io_args_out_4(pipe2_io_args_out_4),
    .io_args_out_5(pipe2_io_args_out_5),
    .io_args_out_6(pipe2_io_args_out_6),
    .io_vliw_out_0(pipe2_io_vliw_out_0),
    .io_vliw_out_1(pipe2_io_vliw_out_1),
    .io_vliw_out_2(pipe2_io_vliw_out_2),
    .io_vliw_out_3(pipe2_io_vliw_out_3),
    .io_offset_out_0(pipe2_io_offset_out_0),
    .io_offset_out_1(pipe2_io_offset_out_1),
    .io_offset_out_2(pipe2_io_offset_out_2),
    .io_offset_out_3(pipe2_io_offset_out_3),
    .io_length_out_0(pipe2_io_length_out_0),
    .io_length_out_1(pipe2_io_length_out_1),
    .io_length_out_2(pipe2_io_length_out_2),
    .io_length_out_3(pipe2_io_length_out_3)
  );
  PrimitiveGetSource pipe3 ( // @[executor.scala 491:23]
    .clock(pipe3_clock),
    .io_pipe_phv_in_data_0(pipe3_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe3_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe3_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe3_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe3_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe3_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe3_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe3_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe3_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe3_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe3_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe3_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe3_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe3_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe3_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe3_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe3_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe3_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe3_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe3_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe3_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe3_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe3_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe3_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe3_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe3_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe3_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe3_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe3_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe3_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe3_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe3_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe3_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe3_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe3_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe3_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe3_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe3_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe3_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe3_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe3_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe3_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe3_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe3_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe3_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe3_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe3_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe3_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe3_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe3_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe3_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe3_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe3_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe3_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe3_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe3_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe3_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe3_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe3_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe3_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe3_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe3_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe3_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe3_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe3_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe3_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe3_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe3_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe3_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe3_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe3_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe3_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe3_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe3_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe3_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe3_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe3_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe3_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe3_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe3_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe3_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe3_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe3_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe3_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe3_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe3_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe3_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe3_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe3_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe3_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe3_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe3_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe3_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe3_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe3_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe3_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe3_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe3_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe3_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe3_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe3_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe3_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe3_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe3_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe3_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe3_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe3_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe3_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe3_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe3_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe3_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe3_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe3_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe3_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe3_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe3_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe3_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe3_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe3_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe3_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe3_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe3_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe3_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe3_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe3_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe3_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe3_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe3_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe3_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe3_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe3_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe3_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe3_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe3_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe3_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe3_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe3_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe3_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe3_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe3_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe3_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe3_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe3_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe3_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe3_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe3_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe3_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe3_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe3_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe3_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe3_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe3_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe3_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe3_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe3_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe3_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe3_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe3_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe3_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe3_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe3_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe3_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe3_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe3_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe3_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe3_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe3_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe3_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe3_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe3_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe3_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe3_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe3_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe3_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe3_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe3_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe3_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe3_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe3_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe3_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe3_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe3_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe3_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe3_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe3_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe3_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe3_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe3_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe3_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe3_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe3_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe3_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe3_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe3_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe3_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe3_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe3_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe3_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe3_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe3_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe3_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe3_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe3_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe3_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe3_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe3_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe3_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe3_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe3_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe3_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe3_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe3_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe3_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe3_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe3_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe3_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe3_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe3_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe3_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe3_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe3_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe3_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe3_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe3_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe3_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe3_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe3_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe3_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe3_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe3_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe3_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe3_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe3_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe3_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe3_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe3_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe3_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe3_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe3_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe3_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe3_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe3_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe3_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe3_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe3_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe3_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe3_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe3_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe3_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe3_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe3_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe3_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe3_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe3_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe3_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe3_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe3_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe3_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe3_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe3_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe3_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe3_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe3_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe3_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe3_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe3_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe3_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe3_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe3_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe3_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe3_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe3_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe3_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe3_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe3_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe3_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe3_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe3_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe3_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe3_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe3_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe3_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe3_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe3_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe3_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe3_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe3_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe3_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe3_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe3_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe3_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe3_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe3_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe3_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe3_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe3_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe3_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe3_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe3_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe3_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe3_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe3_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe3_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe3_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe3_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe3_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe3_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe3_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe3_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe3_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe3_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe3_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe3_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe3_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe3_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe3_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe3_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe3_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe3_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe3_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe3_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe3_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe3_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe3_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe3_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe3_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe3_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe3_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe3_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe3_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe3_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe3_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe3_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe3_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe3_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe3_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe3_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe3_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe3_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe3_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe3_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe3_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe3_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe3_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe3_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe3_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe3_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe3_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe3_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe3_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe3_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe3_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe3_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe3_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe3_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe3_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe3_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe3_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe3_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe3_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe3_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe3_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe3_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe3_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe3_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe3_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe3_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe3_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe3_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe3_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe3_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe3_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe3_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe3_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe3_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe3_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe3_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe3_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe3_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe3_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe3_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe3_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe3_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe3_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe3_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe3_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe3_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe3_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe3_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe3_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe3_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe3_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe3_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe3_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe3_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe3_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe3_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe3_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe3_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe3_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe3_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe3_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe3_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe3_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe3_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe3_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe3_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe3_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe3_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe3_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe3_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe3_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe3_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe3_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe3_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe3_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe3_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe3_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe3_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe3_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe3_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe3_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe3_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe3_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe3_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe3_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe3_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe3_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe3_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe3_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe3_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe3_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe3_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe3_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe3_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe3_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe3_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe3_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe3_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe3_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe3_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe3_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe3_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe3_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe3_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe3_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe3_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe3_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe3_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe3_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe3_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe3_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe3_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe3_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe3_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe3_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe3_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe3_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe3_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe3_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe3_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe3_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe3_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe3_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe3_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe3_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe3_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe3_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe3_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe3_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe3_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe3_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe3_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe3_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe3_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe3_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe3_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe3_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe3_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe3_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe3_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe3_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe3_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe3_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe3_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe3_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe3_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe3_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe3_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe3_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe3_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe3_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe3_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe3_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe3_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe3_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe3_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe3_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe3_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe3_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe3_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe3_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe3_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe3_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe3_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe3_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe3_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe3_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe3_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe3_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe3_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe3_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe3_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe3_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe3_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe3_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe3_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe3_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe3_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe3_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe3_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe3_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe3_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe3_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe3_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe3_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe3_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe3_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe3_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe3_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe3_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe3_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe3_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe3_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe3_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe3_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe3_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe3_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe3_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe3_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe3_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe3_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe3_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe3_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe3_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe3_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe3_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe3_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe3_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe3_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe3_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe3_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe3_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe3_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe3_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe3_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe3_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe3_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe3_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe3_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe3_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe3_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe3_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe3_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe3_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe3_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe3_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe3_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe3_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe3_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe3_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe3_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe3_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe3_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe3_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe3_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe3_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe3_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe3_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe3_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe3_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe3_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe3_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe3_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe3_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe3_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe3_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe3_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe3_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe3_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe3_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe3_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe3_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe3_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe3_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe3_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe3_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe3_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe3_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe3_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe3_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe3_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe3_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe3_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe3_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe3_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe3_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe3_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe3_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe3_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe3_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe3_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe3_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe3_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe3_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe3_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe3_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe3_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe3_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe3_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe3_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe3_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe3_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe3_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe3_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe3_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe3_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe3_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe3_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe3_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe3_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe3_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe3_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe3_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe3_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe3_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe3_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe3_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe3_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe3_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe3_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe3_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe3_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe3_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe3_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe3_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe3_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe3_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe3_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe3_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe3_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe3_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe3_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe3_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe3_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe3_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe3_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe3_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe3_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe3_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe3_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe3_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe3_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe3_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe3_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe3_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe3_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe3_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe3_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe3_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe3_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe3_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe3_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe3_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe3_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe3_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe3_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe3_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe3_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe3_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe3_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe3_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe3_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe3_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe3_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe3_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe3_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe3_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe3_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe3_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe3_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe3_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe3_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe3_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe3_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe3_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe3_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe3_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe3_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe3_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe3_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe3_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe3_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe3_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe3_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe3_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe3_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe3_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe3_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe3_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe3_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe3_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe3_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe3_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe3_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe3_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe3_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe3_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe3_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe3_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe3_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe3_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe3_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe3_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe3_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe3_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe3_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe3_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe3_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe3_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe3_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe3_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe3_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe3_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe3_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe3_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe3_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe3_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe3_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe3_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe3_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe3_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe3_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe3_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe3_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe3_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe3_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe3_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe3_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe3_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe3_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe3_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe3_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe3_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe3_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe3_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe3_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe3_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe3_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe3_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe3_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe3_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe3_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe3_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe3_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe3_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe3_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe3_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe3_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe3_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe3_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe3_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe3_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe3_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe3_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe3_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe3_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe3_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe3_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe3_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe3_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe3_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe3_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe3_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe3_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe3_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe3_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe3_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe3_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe3_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe3_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe3_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe3_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe3_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe3_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe3_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe3_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe3_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe3_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe3_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe3_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe3_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe3_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe3_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe3_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe3_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe3_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe3_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe3_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe3_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe3_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe3_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe3_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe3_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe3_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe3_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe3_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe3_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe3_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe3_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe3_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe3_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe3_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe3_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe3_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe3_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe3_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe3_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe3_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe3_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe3_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe3_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe3_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe3_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe3_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe3_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe3_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe3_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe3_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe3_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe3_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe3_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe3_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe3_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe3_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe3_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe3_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe3_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe3_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe3_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe3_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe3_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe3_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe3_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe3_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe3_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe3_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe3_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe3_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe3_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe3_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe3_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe3_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe3_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe3_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe3_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe3_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe3_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe3_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe3_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe3_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe3_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe3_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe3_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe3_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe3_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe3_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe3_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe3_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe3_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe3_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe3_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe3_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe3_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe3_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe3_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe3_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe3_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe3_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe3_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe3_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe3_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe3_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe3_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe3_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe3_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe3_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe3_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe3_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe3_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe3_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe3_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe3_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe3_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe3_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe3_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe3_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe3_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe3_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe3_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe3_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe3_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe3_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe3_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe3_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe3_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe3_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe3_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe3_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe3_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe3_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe3_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe3_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe3_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe3_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe3_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe3_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe3_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe3_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe3_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe3_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe3_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe3_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe3_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe3_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe3_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe3_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe3_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe3_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe3_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe3_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe3_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe3_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe3_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe3_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe3_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe3_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe3_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe3_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe3_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe3_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe3_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe3_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe3_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe3_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe3_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe3_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe3_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe3_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe3_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe3_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe3_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe3_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe3_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe3_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe3_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe3_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe3_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe3_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe3_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe3_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe3_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe3_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe3_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe3_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe3_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe3_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe3_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe3_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe3_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe3_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe3_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe3_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe3_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe3_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe3_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe3_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe3_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe3_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe3_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe3_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe3_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe3_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe3_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe3_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe3_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe3_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe3_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe3_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe3_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe3_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe3_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe3_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe3_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe3_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe3_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe3_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe3_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe3_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe3_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe3_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe3_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe3_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe3_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe3_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe3_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe3_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe3_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe3_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe3_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe3_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe3_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe3_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe3_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe3_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe3_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe3_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe3_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe3_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe3_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe3_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe3_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe3_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe3_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe3_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe3_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe3_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe3_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe3_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe3_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe3_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe3_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe3_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe3_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe3_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe3_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe3_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe3_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe3_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe3_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe3_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe3_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe3_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe3_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe3_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe3_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe3_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe3_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe3_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe3_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe3_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe3_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe3_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe3_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe3_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe3_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe3_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe3_io_pipe_phv_out_is_valid_processor),
    .io_args_in_0(pipe3_io_args_in_0),
    .io_args_in_1(pipe3_io_args_in_1),
    .io_args_in_2(pipe3_io_args_in_2),
    .io_args_in_3(pipe3_io_args_in_3),
    .io_args_in_4(pipe3_io_args_in_4),
    .io_args_in_5(pipe3_io_args_in_5),
    .io_args_in_6(pipe3_io_args_in_6),
    .io_vliw_in_0(pipe3_io_vliw_in_0),
    .io_vliw_in_1(pipe3_io_vliw_in_1),
    .io_vliw_in_2(pipe3_io_vliw_in_2),
    .io_vliw_in_3(pipe3_io_vliw_in_3),
    .io_offset_in_0(pipe3_io_offset_in_0),
    .io_offset_in_1(pipe3_io_offset_in_1),
    .io_offset_in_2(pipe3_io_offset_in_2),
    .io_offset_in_3(pipe3_io_offset_in_3),
    .io_length_in_0(pipe3_io_length_in_0),
    .io_length_in_1(pipe3_io_length_in_1),
    .io_length_in_2(pipe3_io_length_in_2),
    .io_length_in_3(pipe3_io_length_in_3),
    .io_vliw_out_0(pipe3_io_vliw_out_0),
    .io_vliw_out_1(pipe3_io_vliw_out_1),
    .io_vliw_out_2(pipe3_io_vliw_out_2),
    .io_vliw_out_3(pipe3_io_vliw_out_3),
    .io_field_out_0(pipe3_io_field_out_0),
    .io_field_out_1(pipe3_io_field_out_1),
    .io_field_out_2(pipe3_io_field_out_2),
    .io_field_out_3(pipe3_io_field_out_3),
    .io_mask_out_0(pipe3_io_mask_out_0),
    .io_mask_out_1(pipe3_io_mask_out_1),
    .io_mask_out_2(pipe3_io_mask_out_2),
    .io_mask_out_3(pipe3_io_mask_out_3),
    .io_bias_out_0(pipe3_io_bias_out_0),
    .io_bias_out_1(pipe3_io_bias_out_1),
    .io_bias_out_2(pipe3_io_bias_out_2),
    .io_bias_out_3(pipe3_io_bias_out_3)
  );
  PrimitiveShiftSource pipe4 ( // @[executor.scala 492:23]
    .clock(pipe4_clock),
    .io_pipe_phv_in_data_0(pipe4_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe4_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe4_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe4_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe4_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe4_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe4_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe4_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe4_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe4_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe4_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe4_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe4_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe4_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe4_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe4_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe4_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe4_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe4_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe4_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe4_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe4_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe4_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe4_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe4_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe4_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe4_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe4_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe4_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe4_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe4_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe4_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe4_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe4_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe4_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe4_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe4_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe4_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe4_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe4_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe4_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe4_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe4_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe4_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe4_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe4_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe4_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe4_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe4_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe4_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe4_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe4_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe4_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe4_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe4_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe4_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe4_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe4_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe4_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe4_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe4_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe4_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe4_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe4_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe4_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe4_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe4_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe4_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe4_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe4_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe4_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe4_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe4_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe4_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe4_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe4_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe4_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe4_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe4_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe4_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe4_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe4_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe4_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe4_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe4_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe4_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe4_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe4_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe4_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe4_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe4_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe4_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe4_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe4_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe4_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe4_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe4_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe4_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe4_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe4_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe4_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe4_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe4_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe4_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe4_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe4_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe4_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe4_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe4_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe4_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe4_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe4_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe4_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe4_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe4_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe4_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe4_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe4_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe4_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe4_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe4_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe4_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe4_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe4_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe4_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe4_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe4_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe4_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe4_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe4_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe4_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe4_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe4_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe4_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe4_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe4_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe4_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe4_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe4_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe4_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe4_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe4_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe4_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe4_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe4_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe4_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe4_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe4_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe4_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe4_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe4_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe4_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe4_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe4_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe4_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe4_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe4_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe4_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe4_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe4_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe4_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe4_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe4_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe4_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe4_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe4_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe4_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe4_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe4_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe4_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe4_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe4_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe4_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe4_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe4_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe4_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe4_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe4_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe4_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe4_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe4_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe4_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe4_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe4_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe4_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe4_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe4_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe4_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe4_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe4_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe4_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe4_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe4_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe4_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe4_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe4_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe4_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe4_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe4_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe4_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe4_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe4_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe4_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe4_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe4_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe4_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe4_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe4_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe4_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe4_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe4_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe4_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe4_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe4_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe4_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe4_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe4_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe4_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe4_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe4_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe4_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe4_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe4_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe4_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe4_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe4_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe4_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe4_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe4_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe4_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe4_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe4_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe4_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe4_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe4_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe4_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe4_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe4_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe4_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe4_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe4_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe4_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe4_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe4_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe4_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe4_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe4_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe4_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe4_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe4_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe4_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe4_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe4_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe4_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe4_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe4_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe4_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe4_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe4_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe4_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe4_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe4_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe4_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe4_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe4_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe4_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe4_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe4_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe4_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe4_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe4_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe4_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe4_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe4_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe4_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe4_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe4_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe4_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe4_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe4_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe4_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe4_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe4_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe4_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe4_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe4_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe4_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe4_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe4_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe4_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe4_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe4_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe4_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe4_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe4_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe4_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe4_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe4_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe4_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe4_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe4_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe4_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe4_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe4_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe4_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe4_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe4_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe4_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe4_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe4_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe4_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe4_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe4_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe4_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe4_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe4_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe4_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe4_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe4_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe4_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe4_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe4_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe4_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe4_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe4_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe4_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe4_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe4_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe4_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe4_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe4_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe4_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe4_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe4_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe4_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe4_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe4_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe4_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe4_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe4_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe4_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe4_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe4_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe4_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe4_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe4_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe4_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe4_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe4_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe4_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe4_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe4_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe4_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe4_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe4_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe4_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe4_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe4_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe4_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe4_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe4_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe4_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe4_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe4_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe4_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe4_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe4_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe4_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe4_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe4_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe4_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe4_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe4_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe4_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe4_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe4_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe4_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe4_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe4_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe4_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe4_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe4_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe4_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe4_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe4_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe4_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe4_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe4_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe4_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe4_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe4_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe4_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe4_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe4_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe4_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe4_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe4_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe4_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe4_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe4_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe4_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe4_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe4_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe4_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe4_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe4_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe4_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe4_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe4_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe4_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe4_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe4_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe4_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe4_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe4_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe4_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe4_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe4_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe4_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe4_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe4_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe4_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe4_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe4_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe4_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe4_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe4_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe4_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe4_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe4_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe4_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe4_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe4_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe4_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe4_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe4_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe4_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe4_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe4_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe4_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe4_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe4_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe4_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe4_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe4_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe4_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe4_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe4_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe4_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe4_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe4_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe4_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe4_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe4_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe4_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe4_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe4_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe4_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe4_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe4_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe4_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe4_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe4_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe4_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe4_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe4_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe4_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe4_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe4_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe4_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe4_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe4_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe4_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe4_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe4_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe4_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe4_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe4_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe4_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe4_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe4_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe4_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe4_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe4_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe4_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe4_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe4_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe4_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe4_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe4_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe4_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe4_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe4_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe4_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe4_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe4_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe4_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe4_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe4_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe4_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe4_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe4_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe4_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe4_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe4_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe4_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe4_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe4_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe4_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe4_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe4_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe4_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe4_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe4_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe4_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe4_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe4_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe4_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe4_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe4_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe4_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe4_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe4_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe4_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe4_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe4_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe4_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe4_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe4_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe4_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe4_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe4_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe4_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe4_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe4_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe4_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe4_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe4_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe4_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe4_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe4_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe4_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe4_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe4_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe4_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe4_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe4_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe4_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe4_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe4_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe4_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe4_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe4_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe4_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe4_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe4_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe4_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe4_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe4_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe4_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe4_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe4_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe4_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe4_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe4_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe4_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe4_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe4_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe4_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe4_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe4_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe4_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe4_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe4_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe4_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe4_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe4_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe4_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe4_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe4_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe4_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe4_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe4_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe4_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe4_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe4_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe4_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe4_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe4_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe4_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe4_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe4_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe4_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe4_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe4_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe4_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe4_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe4_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe4_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe4_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe4_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe4_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe4_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe4_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe4_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe4_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe4_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe4_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe4_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe4_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe4_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe4_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe4_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe4_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe4_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe4_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe4_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe4_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe4_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe4_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe4_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe4_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe4_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe4_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe4_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe4_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe4_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe4_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe4_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe4_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe4_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe4_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe4_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe4_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe4_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe4_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe4_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe4_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe4_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe4_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe4_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe4_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe4_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe4_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe4_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe4_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe4_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe4_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe4_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe4_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe4_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe4_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe4_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe4_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe4_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe4_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe4_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe4_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe4_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe4_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe4_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe4_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe4_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe4_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe4_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe4_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe4_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe4_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe4_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe4_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe4_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe4_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe4_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe4_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe4_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe4_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe4_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe4_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe4_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe4_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe4_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe4_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe4_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe4_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe4_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe4_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe4_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe4_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe4_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe4_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe4_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe4_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe4_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe4_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe4_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe4_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe4_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe4_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe4_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe4_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe4_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe4_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe4_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe4_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe4_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe4_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe4_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe4_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe4_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe4_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe4_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe4_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe4_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe4_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe4_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe4_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe4_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe4_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe4_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe4_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe4_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe4_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe4_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe4_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe4_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe4_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe4_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe4_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe4_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe4_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe4_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe4_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe4_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe4_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe4_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe4_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe4_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe4_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe4_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe4_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe4_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe4_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe4_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe4_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe4_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe4_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe4_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe4_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe4_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe4_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe4_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe4_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe4_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe4_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe4_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe4_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe4_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe4_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe4_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe4_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe4_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe4_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe4_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe4_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe4_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe4_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe4_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe4_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe4_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe4_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe4_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe4_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe4_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe4_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe4_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe4_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe4_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe4_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe4_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe4_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe4_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe4_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe4_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe4_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe4_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe4_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe4_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe4_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe4_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe4_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe4_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe4_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe4_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe4_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe4_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe4_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe4_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe4_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe4_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe4_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe4_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe4_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe4_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe4_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe4_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe4_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe4_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe4_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe4_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe4_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe4_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe4_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe4_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe4_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe4_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe4_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe4_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe4_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe4_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe4_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe4_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe4_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe4_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe4_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe4_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe4_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe4_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe4_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe4_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe4_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe4_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe4_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe4_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe4_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe4_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe4_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe4_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe4_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe4_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe4_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe4_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe4_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe4_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe4_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe4_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe4_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe4_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe4_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe4_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe4_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe4_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe4_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe4_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe4_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe4_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe4_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe4_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe4_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe4_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe4_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe4_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe4_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe4_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe4_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe4_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe4_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe4_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe4_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe4_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe4_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe4_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe4_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe4_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe4_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe4_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe4_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe4_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe4_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe4_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe4_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe4_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe4_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe4_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe4_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe4_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe4_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe4_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe4_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe4_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe4_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe4_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe4_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe4_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe4_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe4_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe4_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe4_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe4_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe4_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe4_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe4_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe4_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe4_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe4_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe4_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe4_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe4_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe4_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe4_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe4_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe4_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe4_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe4_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe4_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe4_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe4_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe4_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe4_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe4_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe4_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe4_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe4_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe4_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe4_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe4_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe4_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe4_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe4_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe4_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe4_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe4_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe4_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe4_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe4_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe4_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe4_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe4_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe4_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe4_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe4_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe4_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe4_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe4_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe4_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe4_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe4_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe4_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe4_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe4_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe4_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe4_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe4_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe4_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe4_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe4_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe4_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe4_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe4_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe4_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe4_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe4_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe4_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe4_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe4_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe4_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe4_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe4_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe4_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe4_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe4_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe4_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe4_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe4_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe4_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe4_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe4_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe4_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe4_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe4_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe4_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe4_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe4_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe4_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe4_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe4_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe4_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe4_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe4_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe4_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe4_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe4_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe4_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe4_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe4_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe4_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe4_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe4_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe4_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe4_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe4_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe4_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe4_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe4_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe4_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe4_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe4_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe4_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe4_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe4_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe4_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe4_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe4_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe4_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe4_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe4_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe4_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe4_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe4_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe4_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe4_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe4_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe4_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe4_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe4_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe4_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe4_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe4_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe4_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe4_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe4_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe4_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe4_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe4_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe4_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe4_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe4_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe4_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe4_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe4_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe4_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe4_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe4_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe4_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe4_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe4_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe4_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe4_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe4_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe4_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe4_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe4_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe4_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe4_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe4_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe4_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe4_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe4_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe4_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe4_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe4_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe4_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe4_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe4_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe4_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe4_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe4_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe4_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe4_io_pipe_phv_out_is_valid_processor),
    .io_vliw_in_0(pipe4_io_vliw_in_0),
    .io_vliw_in_1(pipe4_io_vliw_in_1),
    .io_vliw_in_2(pipe4_io_vliw_in_2),
    .io_vliw_in_3(pipe4_io_vliw_in_3),
    .io_field_in_0(pipe4_io_field_in_0),
    .io_field_in_1(pipe4_io_field_in_1),
    .io_field_in_2(pipe4_io_field_in_2),
    .io_field_in_3(pipe4_io_field_in_3),
    .io_mask_in_0(pipe4_io_mask_in_0),
    .io_mask_in_1(pipe4_io_mask_in_1),
    .io_mask_in_2(pipe4_io_mask_in_2),
    .io_mask_in_3(pipe4_io_mask_in_3),
    .io_bias_in_0(pipe4_io_bias_in_0),
    .io_bias_in_1(pipe4_io_bias_in_1),
    .io_bias_in_2(pipe4_io_bias_in_2),
    .io_bias_in_3(pipe4_io_bias_in_3),
    .io_vliw_out_0(pipe4_io_vliw_out_0),
    .io_vliw_out_1(pipe4_io_vliw_out_1),
    .io_vliw_out_2(pipe4_io_vliw_out_2),
    .io_vliw_out_3(pipe4_io_vliw_out_3),
    .io_field_out_0(pipe4_io_field_out_0),
    .io_field_out_1(pipe4_io_field_out_1),
    .io_field_out_2(pipe4_io_field_out_2),
    .io_field_out_3(pipe4_io_field_out_3),
    .io_mask_out_0(pipe4_io_mask_out_0),
    .io_mask_out_1(pipe4_io_mask_out_1),
    .io_mask_out_2(pipe4_io_mask_out_2),
    .io_mask_out_3(pipe4_io_mask_out_3),
    .io_bias_out_0(pipe4_io_bias_out_0),
    .io_bias_out_1(pipe4_io_bias_out_1),
    .io_bias_out_2(pipe4_io_bias_out_2),
    .io_bias_out_3(pipe4_io_bias_out_3),
    .io_dst_offset_out_0(pipe4_io_dst_offset_out_0),
    .io_dst_offset_out_1(pipe4_io_dst_offset_out_1),
    .io_dst_offset_out_2(pipe4_io_dst_offset_out_2),
    .io_dst_offset_out_3(pipe4_io_dst_offset_out_3)
  );
  PrimitiveALU pipe5 ( // @[executor.scala 493:23]
    .clock(pipe5_clock),
    .io_pipe_phv_in_data_0(pipe5_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe5_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe5_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe5_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe5_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe5_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe5_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe5_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe5_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe5_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe5_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe5_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe5_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe5_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe5_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe5_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe5_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe5_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe5_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe5_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe5_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe5_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe5_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe5_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe5_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe5_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe5_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe5_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe5_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe5_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe5_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe5_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe5_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe5_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe5_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe5_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe5_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe5_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe5_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe5_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe5_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe5_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe5_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe5_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe5_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe5_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe5_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe5_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe5_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe5_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe5_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe5_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe5_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe5_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe5_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe5_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe5_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe5_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe5_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe5_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe5_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe5_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe5_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe5_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe5_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe5_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe5_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe5_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe5_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe5_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe5_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe5_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe5_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe5_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe5_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe5_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe5_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe5_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe5_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe5_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe5_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe5_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe5_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe5_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe5_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe5_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe5_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe5_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe5_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe5_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe5_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe5_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe5_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe5_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe5_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe5_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe5_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe5_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe5_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe5_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe5_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe5_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe5_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe5_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe5_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe5_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe5_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe5_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe5_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe5_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe5_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe5_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe5_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe5_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe5_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe5_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe5_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe5_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe5_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe5_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe5_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe5_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe5_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe5_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe5_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe5_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe5_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe5_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe5_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe5_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe5_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe5_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe5_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe5_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe5_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe5_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe5_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe5_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe5_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe5_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe5_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe5_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe5_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe5_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe5_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe5_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe5_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe5_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe5_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe5_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe5_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe5_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe5_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe5_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe5_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe5_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe5_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe5_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe5_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe5_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe5_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe5_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe5_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe5_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe5_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe5_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe5_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe5_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe5_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe5_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe5_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe5_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe5_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe5_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe5_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe5_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe5_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe5_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe5_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe5_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe5_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe5_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe5_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe5_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe5_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe5_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe5_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe5_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe5_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe5_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe5_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe5_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe5_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe5_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe5_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe5_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe5_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe5_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe5_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe5_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe5_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe5_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe5_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe5_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe5_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe5_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe5_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe5_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe5_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe5_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe5_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe5_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe5_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe5_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe5_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe5_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe5_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe5_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe5_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe5_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe5_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe5_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe5_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe5_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe5_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe5_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe5_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe5_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe5_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe5_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe5_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe5_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe5_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe5_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe5_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe5_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe5_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe5_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe5_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe5_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe5_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe5_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe5_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe5_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe5_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe5_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe5_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe5_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe5_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe5_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe5_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe5_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe5_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe5_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe5_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe5_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe5_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe5_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe5_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe5_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe5_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe5_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe5_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe5_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe5_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe5_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe5_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe5_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe5_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe5_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe5_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe5_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe5_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe5_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe5_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe5_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe5_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe5_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe5_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe5_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe5_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe5_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe5_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe5_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe5_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe5_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe5_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe5_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe5_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe5_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe5_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe5_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe5_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe5_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe5_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe5_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe5_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe5_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe5_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe5_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe5_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe5_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe5_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe5_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe5_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe5_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe5_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe5_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe5_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe5_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe5_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe5_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe5_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe5_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe5_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe5_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe5_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe5_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe5_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe5_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe5_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe5_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe5_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe5_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe5_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe5_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe5_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe5_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe5_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe5_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe5_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe5_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe5_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe5_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe5_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe5_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe5_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe5_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe5_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe5_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe5_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe5_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe5_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe5_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe5_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe5_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe5_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe5_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe5_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe5_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe5_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe5_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe5_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe5_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe5_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe5_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe5_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe5_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe5_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe5_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe5_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe5_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe5_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe5_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe5_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe5_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe5_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe5_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe5_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe5_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe5_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe5_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe5_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe5_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe5_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe5_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe5_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe5_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe5_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe5_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe5_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe5_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe5_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe5_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe5_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe5_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe5_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe5_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe5_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe5_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe5_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe5_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe5_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe5_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe5_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe5_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe5_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe5_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe5_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe5_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe5_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe5_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe5_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe5_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe5_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe5_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe5_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe5_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe5_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe5_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe5_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe5_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe5_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe5_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe5_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe5_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe5_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe5_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe5_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe5_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe5_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe5_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe5_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe5_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe5_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe5_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe5_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe5_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe5_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe5_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe5_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe5_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe5_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe5_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe5_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe5_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe5_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe5_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe5_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe5_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe5_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe5_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe5_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe5_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe5_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe5_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe5_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe5_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe5_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe5_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe5_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe5_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe5_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe5_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe5_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe5_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe5_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe5_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe5_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe5_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe5_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe5_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe5_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe5_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe5_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe5_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe5_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe5_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe5_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe5_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe5_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe5_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe5_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe5_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe5_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe5_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe5_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe5_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe5_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe5_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe5_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe5_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe5_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe5_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe5_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe5_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe5_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe5_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe5_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe5_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe5_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe5_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe5_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe5_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe5_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe5_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe5_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe5_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe5_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe5_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe5_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe5_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe5_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe5_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe5_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe5_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe5_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe5_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe5_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe5_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe5_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe5_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe5_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe5_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe5_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe5_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe5_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe5_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe5_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe5_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe5_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe5_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe5_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe5_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe5_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe5_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe5_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe5_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe5_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe5_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe5_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe5_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe5_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe5_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe5_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe5_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe5_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe5_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe5_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe5_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe5_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe5_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe5_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe5_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe5_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe5_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe5_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe5_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe5_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe5_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe5_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe5_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe5_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe5_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe5_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe5_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe5_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe5_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe5_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe5_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe5_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe5_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe5_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe5_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe5_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe5_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe5_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe5_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe5_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe5_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe5_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe5_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe5_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe5_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe5_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe5_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe5_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe5_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe5_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe5_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe5_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe5_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe5_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe5_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe5_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe5_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe5_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe5_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe5_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe5_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe5_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe5_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe5_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe5_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe5_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe5_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe5_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe5_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe5_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe5_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe5_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe5_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe5_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe5_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe5_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe5_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe5_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe5_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe5_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe5_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe5_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe5_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe5_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe5_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe5_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe5_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe5_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe5_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe5_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe5_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe5_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe5_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe5_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe5_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe5_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe5_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe5_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe5_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe5_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe5_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe5_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe5_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe5_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe5_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe5_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe5_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe5_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe5_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe5_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe5_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe5_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe5_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe5_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe5_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe5_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe5_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe5_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe5_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe5_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe5_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe5_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe5_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe5_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe5_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe5_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe5_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe5_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe5_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe5_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe5_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe5_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe5_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe5_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe5_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe5_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe5_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe5_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe5_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe5_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe5_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe5_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe5_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe5_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe5_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe5_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe5_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe5_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe5_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe5_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe5_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe5_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe5_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe5_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe5_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe5_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe5_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe5_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe5_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe5_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe5_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe5_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe5_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe5_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe5_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe5_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe5_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe5_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe5_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe5_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe5_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe5_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe5_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe5_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe5_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe5_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe5_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe5_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe5_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe5_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe5_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe5_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe5_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe5_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe5_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe5_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe5_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe5_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe5_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe5_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe5_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe5_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe5_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe5_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe5_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe5_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe5_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe5_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe5_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe5_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe5_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe5_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe5_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe5_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe5_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe5_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe5_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe5_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe5_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe5_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe5_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe5_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe5_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe5_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe5_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe5_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe5_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe5_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe5_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe5_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe5_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe5_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe5_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe5_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe5_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe5_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe5_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe5_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe5_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe5_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe5_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe5_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe5_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe5_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe5_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe5_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe5_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe5_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe5_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe5_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe5_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe5_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe5_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe5_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe5_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe5_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe5_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe5_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe5_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe5_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe5_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe5_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe5_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe5_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe5_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe5_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe5_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe5_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe5_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe5_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe5_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe5_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe5_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe5_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe5_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe5_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe5_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe5_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe5_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe5_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe5_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe5_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe5_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe5_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe5_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe5_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe5_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe5_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe5_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe5_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe5_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe5_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe5_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe5_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe5_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe5_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe5_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe5_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe5_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe5_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe5_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe5_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe5_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe5_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe5_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe5_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe5_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe5_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe5_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe5_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe5_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe5_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe5_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe5_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe5_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe5_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe5_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe5_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe5_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe5_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe5_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe5_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe5_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe5_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe5_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe5_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe5_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe5_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe5_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe5_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe5_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe5_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe5_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe5_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe5_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe5_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe5_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe5_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe5_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe5_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe5_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe5_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe5_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe5_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe5_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe5_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe5_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe5_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe5_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe5_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe5_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe5_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe5_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe5_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe5_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe5_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe5_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe5_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe5_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe5_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe5_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe5_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe5_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe5_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe5_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe5_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe5_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe5_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe5_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe5_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe5_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe5_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe5_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe5_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe5_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe5_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe5_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe5_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe5_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe5_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe5_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe5_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe5_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe5_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe5_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe5_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe5_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe5_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe5_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe5_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe5_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe5_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe5_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe5_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe5_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe5_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe5_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe5_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe5_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe5_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe5_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe5_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe5_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe5_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe5_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe5_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe5_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe5_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe5_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe5_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe5_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe5_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe5_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe5_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe5_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe5_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe5_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe5_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe5_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe5_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe5_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe5_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe5_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe5_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe5_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe5_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe5_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe5_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe5_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe5_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe5_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe5_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe5_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe5_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe5_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe5_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe5_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe5_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe5_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe5_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe5_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe5_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe5_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe5_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe5_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe5_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe5_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe5_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe5_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe5_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe5_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe5_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe5_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe5_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe5_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe5_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe5_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe5_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe5_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe5_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe5_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe5_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe5_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe5_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe5_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe5_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe5_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe5_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe5_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe5_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe5_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe5_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe5_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe5_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe5_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe5_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe5_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe5_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe5_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe5_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe5_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe5_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe5_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe5_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe5_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe5_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe5_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe5_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe5_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe5_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe5_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe5_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe5_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe5_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe5_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe5_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe5_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe5_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe5_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe5_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe5_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe5_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe5_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe5_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe5_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe5_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe5_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe5_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe5_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe5_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe5_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe5_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe5_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe5_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe5_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe5_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe5_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe5_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe5_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe5_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe5_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe5_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe5_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe5_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe5_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe5_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe5_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe5_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe5_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe5_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe5_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe5_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe5_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe5_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe5_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe5_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe5_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe5_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe5_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe5_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe5_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe5_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe5_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe5_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe5_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe5_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe5_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe5_io_pipe_phv_out_next_config_id),
    .io_pipe_phv_out_is_valid_processor(pipe5_io_pipe_phv_out_is_valid_processor),
    .io_vliw_in_0(pipe5_io_vliw_in_0),
    .io_vliw_in_1(pipe5_io_vliw_in_1),
    .io_vliw_in_2(pipe5_io_vliw_in_2),
    .io_vliw_in_3(pipe5_io_vliw_in_3),
    .io_field_in_0(pipe5_io_field_in_0),
    .io_field_in_1(pipe5_io_field_in_1),
    .io_field_in_2(pipe5_io_field_in_2),
    .io_field_in_3(pipe5_io_field_in_3),
    .io_mask_in_0(pipe5_io_mask_in_0),
    .io_mask_in_1(pipe5_io_mask_in_1),
    .io_mask_in_2(pipe5_io_mask_in_2),
    .io_mask_in_3(pipe5_io_mask_in_3),
    .io_bias_in_0(pipe5_io_bias_in_0),
    .io_bias_in_1(pipe5_io_bias_in_1),
    .io_bias_in_2(pipe5_io_bias_in_2),
    .io_bias_in_3(pipe5_io_bias_in_3),
    .io_dst_offset_in_0(pipe5_io_dst_offset_in_0),
    .io_dst_offset_in_1(pipe5_io_dst_offset_in_1),
    .io_dst_offset_in_2(pipe5_io_dst_offset_in_2),
    .io_dst_offset_in_3(pipe5_io_dst_offset_in_3),
    .io_vliw_out_0(pipe5_io_vliw_out_0),
    .io_vliw_out_1(pipe5_io_vliw_out_1),
    .io_vliw_out_2(pipe5_io_vliw_out_2),
    .io_vliw_out_3(pipe5_io_vliw_out_3),
    .io_field_out_0(pipe5_io_field_out_0),
    .io_field_out_1(pipe5_io_field_out_1),
    .io_field_out_2(pipe5_io_field_out_2),
    .io_field_out_3(pipe5_io_field_out_3),
    .io_mask_out_0(pipe5_io_mask_out_0),
    .io_mask_out_1(pipe5_io_mask_out_1),
    .io_mask_out_2(pipe5_io_mask_out_2),
    .io_mask_out_3(pipe5_io_mask_out_3),
    .io_dst_offset_out_0(pipe5_io_dst_offset_out_0),
    .io_dst_offset_out_1(pipe5_io_dst_offset_out_1),
    .io_dst_offset_out_2(pipe5_io_dst_offset_out_2),
    .io_dst_offset_out_3(pipe5_io_dst_offset_out_3)
  );
  PrimitiveWriteBack pipe6 ( // @[executor.scala 494:23]
    .clock(pipe6_clock),
    .io_pipe_phv_in_data_0(pipe6_io_pipe_phv_in_data_0),
    .io_pipe_phv_in_data_1(pipe6_io_pipe_phv_in_data_1),
    .io_pipe_phv_in_data_2(pipe6_io_pipe_phv_in_data_2),
    .io_pipe_phv_in_data_3(pipe6_io_pipe_phv_in_data_3),
    .io_pipe_phv_in_data_4(pipe6_io_pipe_phv_in_data_4),
    .io_pipe_phv_in_data_5(pipe6_io_pipe_phv_in_data_5),
    .io_pipe_phv_in_data_6(pipe6_io_pipe_phv_in_data_6),
    .io_pipe_phv_in_data_7(pipe6_io_pipe_phv_in_data_7),
    .io_pipe_phv_in_data_8(pipe6_io_pipe_phv_in_data_8),
    .io_pipe_phv_in_data_9(pipe6_io_pipe_phv_in_data_9),
    .io_pipe_phv_in_data_10(pipe6_io_pipe_phv_in_data_10),
    .io_pipe_phv_in_data_11(pipe6_io_pipe_phv_in_data_11),
    .io_pipe_phv_in_data_12(pipe6_io_pipe_phv_in_data_12),
    .io_pipe_phv_in_data_13(pipe6_io_pipe_phv_in_data_13),
    .io_pipe_phv_in_data_14(pipe6_io_pipe_phv_in_data_14),
    .io_pipe_phv_in_data_15(pipe6_io_pipe_phv_in_data_15),
    .io_pipe_phv_in_data_16(pipe6_io_pipe_phv_in_data_16),
    .io_pipe_phv_in_data_17(pipe6_io_pipe_phv_in_data_17),
    .io_pipe_phv_in_data_18(pipe6_io_pipe_phv_in_data_18),
    .io_pipe_phv_in_data_19(pipe6_io_pipe_phv_in_data_19),
    .io_pipe_phv_in_data_20(pipe6_io_pipe_phv_in_data_20),
    .io_pipe_phv_in_data_21(pipe6_io_pipe_phv_in_data_21),
    .io_pipe_phv_in_data_22(pipe6_io_pipe_phv_in_data_22),
    .io_pipe_phv_in_data_23(pipe6_io_pipe_phv_in_data_23),
    .io_pipe_phv_in_data_24(pipe6_io_pipe_phv_in_data_24),
    .io_pipe_phv_in_data_25(pipe6_io_pipe_phv_in_data_25),
    .io_pipe_phv_in_data_26(pipe6_io_pipe_phv_in_data_26),
    .io_pipe_phv_in_data_27(pipe6_io_pipe_phv_in_data_27),
    .io_pipe_phv_in_data_28(pipe6_io_pipe_phv_in_data_28),
    .io_pipe_phv_in_data_29(pipe6_io_pipe_phv_in_data_29),
    .io_pipe_phv_in_data_30(pipe6_io_pipe_phv_in_data_30),
    .io_pipe_phv_in_data_31(pipe6_io_pipe_phv_in_data_31),
    .io_pipe_phv_in_data_32(pipe6_io_pipe_phv_in_data_32),
    .io_pipe_phv_in_data_33(pipe6_io_pipe_phv_in_data_33),
    .io_pipe_phv_in_data_34(pipe6_io_pipe_phv_in_data_34),
    .io_pipe_phv_in_data_35(pipe6_io_pipe_phv_in_data_35),
    .io_pipe_phv_in_data_36(pipe6_io_pipe_phv_in_data_36),
    .io_pipe_phv_in_data_37(pipe6_io_pipe_phv_in_data_37),
    .io_pipe_phv_in_data_38(pipe6_io_pipe_phv_in_data_38),
    .io_pipe_phv_in_data_39(pipe6_io_pipe_phv_in_data_39),
    .io_pipe_phv_in_data_40(pipe6_io_pipe_phv_in_data_40),
    .io_pipe_phv_in_data_41(pipe6_io_pipe_phv_in_data_41),
    .io_pipe_phv_in_data_42(pipe6_io_pipe_phv_in_data_42),
    .io_pipe_phv_in_data_43(pipe6_io_pipe_phv_in_data_43),
    .io_pipe_phv_in_data_44(pipe6_io_pipe_phv_in_data_44),
    .io_pipe_phv_in_data_45(pipe6_io_pipe_phv_in_data_45),
    .io_pipe_phv_in_data_46(pipe6_io_pipe_phv_in_data_46),
    .io_pipe_phv_in_data_47(pipe6_io_pipe_phv_in_data_47),
    .io_pipe_phv_in_data_48(pipe6_io_pipe_phv_in_data_48),
    .io_pipe_phv_in_data_49(pipe6_io_pipe_phv_in_data_49),
    .io_pipe_phv_in_data_50(pipe6_io_pipe_phv_in_data_50),
    .io_pipe_phv_in_data_51(pipe6_io_pipe_phv_in_data_51),
    .io_pipe_phv_in_data_52(pipe6_io_pipe_phv_in_data_52),
    .io_pipe_phv_in_data_53(pipe6_io_pipe_phv_in_data_53),
    .io_pipe_phv_in_data_54(pipe6_io_pipe_phv_in_data_54),
    .io_pipe_phv_in_data_55(pipe6_io_pipe_phv_in_data_55),
    .io_pipe_phv_in_data_56(pipe6_io_pipe_phv_in_data_56),
    .io_pipe_phv_in_data_57(pipe6_io_pipe_phv_in_data_57),
    .io_pipe_phv_in_data_58(pipe6_io_pipe_phv_in_data_58),
    .io_pipe_phv_in_data_59(pipe6_io_pipe_phv_in_data_59),
    .io_pipe_phv_in_data_60(pipe6_io_pipe_phv_in_data_60),
    .io_pipe_phv_in_data_61(pipe6_io_pipe_phv_in_data_61),
    .io_pipe_phv_in_data_62(pipe6_io_pipe_phv_in_data_62),
    .io_pipe_phv_in_data_63(pipe6_io_pipe_phv_in_data_63),
    .io_pipe_phv_in_data_64(pipe6_io_pipe_phv_in_data_64),
    .io_pipe_phv_in_data_65(pipe6_io_pipe_phv_in_data_65),
    .io_pipe_phv_in_data_66(pipe6_io_pipe_phv_in_data_66),
    .io_pipe_phv_in_data_67(pipe6_io_pipe_phv_in_data_67),
    .io_pipe_phv_in_data_68(pipe6_io_pipe_phv_in_data_68),
    .io_pipe_phv_in_data_69(pipe6_io_pipe_phv_in_data_69),
    .io_pipe_phv_in_data_70(pipe6_io_pipe_phv_in_data_70),
    .io_pipe_phv_in_data_71(pipe6_io_pipe_phv_in_data_71),
    .io_pipe_phv_in_data_72(pipe6_io_pipe_phv_in_data_72),
    .io_pipe_phv_in_data_73(pipe6_io_pipe_phv_in_data_73),
    .io_pipe_phv_in_data_74(pipe6_io_pipe_phv_in_data_74),
    .io_pipe_phv_in_data_75(pipe6_io_pipe_phv_in_data_75),
    .io_pipe_phv_in_data_76(pipe6_io_pipe_phv_in_data_76),
    .io_pipe_phv_in_data_77(pipe6_io_pipe_phv_in_data_77),
    .io_pipe_phv_in_data_78(pipe6_io_pipe_phv_in_data_78),
    .io_pipe_phv_in_data_79(pipe6_io_pipe_phv_in_data_79),
    .io_pipe_phv_in_data_80(pipe6_io_pipe_phv_in_data_80),
    .io_pipe_phv_in_data_81(pipe6_io_pipe_phv_in_data_81),
    .io_pipe_phv_in_data_82(pipe6_io_pipe_phv_in_data_82),
    .io_pipe_phv_in_data_83(pipe6_io_pipe_phv_in_data_83),
    .io_pipe_phv_in_data_84(pipe6_io_pipe_phv_in_data_84),
    .io_pipe_phv_in_data_85(pipe6_io_pipe_phv_in_data_85),
    .io_pipe_phv_in_data_86(pipe6_io_pipe_phv_in_data_86),
    .io_pipe_phv_in_data_87(pipe6_io_pipe_phv_in_data_87),
    .io_pipe_phv_in_data_88(pipe6_io_pipe_phv_in_data_88),
    .io_pipe_phv_in_data_89(pipe6_io_pipe_phv_in_data_89),
    .io_pipe_phv_in_data_90(pipe6_io_pipe_phv_in_data_90),
    .io_pipe_phv_in_data_91(pipe6_io_pipe_phv_in_data_91),
    .io_pipe_phv_in_data_92(pipe6_io_pipe_phv_in_data_92),
    .io_pipe_phv_in_data_93(pipe6_io_pipe_phv_in_data_93),
    .io_pipe_phv_in_data_94(pipe6_io_pipe_phv_in_data_94),
    .io_pipe_phv_in_data_95(pipe6_io_pipe_phv_in_data_95),
    .io_pipe_phv_in_data_96(pipe6_io_pipe_phv_in_data_96),
    .io_pipe_phv_in_data_97(pipe6_io_pipe_phv_in_data_97),
    .io_pipe_phv_in_data_98(pipe6_io_pipe_phv_in_data_98),
    .io_pipe_phv_in_data_99(pipe6_io_pipe_phv_in_data_99),
    .io_pipe_phv_in_data_100(pipe6_io_pipe_phv_in_data_100),
    .io_pipe_phv_in_data_101(pipe6_io_pipe_phv_in_data_101),
    .io_pipe_phv_in_data_102(pipe6_io_pipe_phv_in_data_102),
    .io_pipe_phv_in_data_103(pipe6_io_pipe_phv_in_data_103),
    .io_pipe_phv_in_data_104(pipe6_io_pipe_phv_in_data_104),
    .io_pipe_phv_in_data_105(pipe6_io_pipe_phv_in_data_105),
    .io_pipe_phv_in_data_106(pipe6_io_pipe_phv_in_data_106),
    .io_pipe_phv_in_data_107(pipe6_io_pipe_phv_in_data_107),
    .io_pipe_phv_in_data_108(pipe6_io_pipe_phv_in_data_108),
    .io_pipe_phv_in_data_109(pipe6_io_pipe_phv_in_data_109),
    .io_pipe_phv_in_data_110(pipe6_io_pipe_phv_in_data_110),
    .io_pipe_phv_in_data_111(pipe6_io_pipe_phv_in_data_111),
    .io_pipe_phv_in_data_112(pipe6_io_pipe_phv_in_data_112),
    .io_pipe_phv_in_data_113(pipe6_io_pipe_phv_in_data_113),
    .io_pipe_phv_in_data_114(pipe6_io_pipe_phv_in_data_114),
    .io_pipe_phv_in_data_115(pipe6_io_pipe_phv_in_data_115),
    .io_pipe_phv_in_data_116(pipe6_io_pipe_phv_in_data_116),
    .io_pipe_phv_in_data_117(pipe6_io_pipe_phv_in_data_117),
    .io_pipe_phv_in_data_118(pipe6_io_pipe_phv_in_data_118),
    .io_pipe_phv_in_data_119(pipe6_io_pipe_phv_in_data_119),
    .io_pipe_phv_in_data_120(pipe6_io_pipe_phv_in_data_120),
    .io_pipe_phv_in_data_121(pipe6_io_pipe_phv_in_data_121),
    .io_pipe_phv_in_data_122(pipe6_io_pipe_phv_in_data_122),
    .io_pipe_phv_in_data_123(pipe6_io_pipe_phv_in_data_123),
    .io_pipe_phv_in_data_124(pipe6_io_pipe_phv_in_data_124),
    .io_pipe_phv_in_data_125(pipe6_io_pipe_phv_in_data_125),
    .io_pipe_phv_in_data_126(pipe6_io_pipe_phv_in_data_126),
    .io_pipe_phv_in_data_127(pipe6_io_pipe_phv_in_data_127),
    .io_pipe_phv_in_data_128(pipe6_io_pipe_phv_in_data_128),
    .io_pipe_phv_in_data_129(pipe6_io_pipe_phv_in_data_129),
    .io_pipe_phv_in_data_130(pipe6_io_pipe_phv_in_data_130),
    .io_pipe_phv_in_data_131(pipe6_io_pipe_phv_in_data_131),
    .io_pipe_phv_in_data_132(pipe6_io_pipe_phv_in_data_132),
    .io_pipe_phv_in_data_133(pipe6_io_pipe_phv_in_data_133),
    .io_pipe_phv_in_data_134(pipe6_io_pipe_phv_in_data_134),
    .io_pipe_phv_in_data_135(pipe6_io_pipe_phv_in_data_135),
    .io_pipe_phv_in_data_136(pipe6_io_pipe_phv_in_data_136),
    .io_pipe_phv_in_data_137(pipe6_io_pipe_phv_in_data_137),
    .io_pipe_phv_in_data_138(pipe6_io_pipe_phv_in_data_138),
    .io_pipe_phv_in_data_139(pipe6_io_pipe_phv_in_data_139),
    .io_pipe_phv_in_data_140(pipe6_io_pipe_phv_in_data_140),
    .io_pipe_phv_in_data_141(pipe6_io_pipe_phv_in_data_141),
    .io_pipe_phv_in_data_142(pipe6_io_pipe_phv_in_data_142),
    .io_pipe_phv_in_data_143(pipe6_io_pipe_phv_in_data_143),
    .io_pipe_phv_in_data_144(pipe6_io_pipe_phv_in_data_144),
    .io_pipe_phv_in_data_145(pipe6_io_pipe_phv_in_data_145),
    .io_pipe_phv_in_data_146(pipe6_io_pipe_phv_in_data_146),
    .io_pipe_phv_in_data_147(pipe6_io_pipe_phv_in_data_147),
    .io_pipe_phv_in_data_148(pipe6_io_pipe_phv_in_data_148),
    .io_pipe_phv_in_data_149(pipe6_io_pipe_phv_in_data_149),
    .io_pipe_phv_in_data_150(pipe6_io_pipe_phv_in_data_150),
    .io_pipe_phv_in_data_151(pipe6_io_pipe_phv_in_data_151),
    .io_pipe_phv_in_data_152(pipe6_io_pipe_phv_in_data_152),
    .io_pipe_phv_in_data_153(pipe6_io_pipe_phv_in_data_153),
    .io_pipe_phv_in_data_154(pipe6_io_pipe_phv_in_data_154),
    .io_pipe_phv_in_data_155(pipe6_io_pipe_phv_in_data_155),
    .io_pipe_phv_in_data_156(pipe6_io_pipe_phv_in_data_156),
    .io_pipe_phv_in_data_157(pipe6_io_pipe_phv_in_data_157),
    .io_pipe_phv_in_data_158(pipe6_io_pipe_phv_in_data_158),
    .io_pipe_phv_in_data_159(pipe6_io_pipe_phv_in_data_159),
    .io_pipe_phv_in_data_160(pipe6_io_pipe_phv_in_data_160),
    .io_pipe_phv_in_data_161(pipe6_io_pipe_phv_in_data_161),
    .io_pipe_phv_in_data_162(pipe6_io_pipe_phv_in_data_162),
    .io_pipe_phv_in_data_163(pipe6_io_pipe_phv_in_data_163),
    .io_pipe_phv_in_data_164(pipe6_io_pipe_phv_in_data_164),
    .io_pipe_phv_in_data_165(pipe6_io_pipe_phv_in_data_165),
    .io_pipe_phv_in_data_166(pipe6_io_pipe_phv_in_data_166),
    .io_pipe_phv_in_data_167(pipe6_io_pipe_phv_in_data_167),
    .io_pipe_phv_in_data_168(pipe6_io_pipe_phv_in_data_168),
    .io_pipe_phv_in_data_169(pipe6_io_pipe_phv_in_data_169),
    .io_pipe_phv_in_data_170(pipe6_io_pipe_phv_in_data_170),
    .io_pipe_phv_in_data_171(pipe6_io_pipe_phv_in_data_171),
    .io_pipe_phv_in_data_172(pipe6_io_pipe_phv_in_data_172),
    .io_pipe_phv_in_data_173(pipe6_io_pipe_phv_in_data_173),
    .io_pipe_phv_in_data_174(pipe6_io_pipe_phv_in_data_174),
    .io_pipe_phv_in_data_175(pipe6_io_pipe_phv_in_data_175),
    .io_pipe_phv_in_data_176(pipe6_io_pipe_phv_in_data_176),
    .io_pipe_phv_in_data_177(pipe6_io_pipe_phv_in_data_177),
    .io_pipe_phv_in_data_178(pipe6_io_pipe_phv_in_data_178),
    .io_pipe_phv_in_data_179(pipe6_io_pipe_phv_in_data_179),
    .io_pipe_phv_in_data_180(pipe6_io_pipe_phv_in_data_180),
    .io_pipe_phv_in_data_181(pipe6_io_pipe_phv_in_data_181),
    .io_pipe_phv_in_data_182(pipe6_io_pipe_phv_in_data_182),
    .io_pipe_phv_in_data_183(pipe6_io_pipe_phv_in_data_183),
    .io_pipe_phv_in_data_184(pipe6_io_pipe_phv_in_data_184),
    .io_pipe_phv_in_data_185(pipe6_io_pipe_phv_in_data_185),
    .io_pipe_phv_in_data_186(pipe6_io_pipe_phv_in_data_186),
    .io_pipe_phv_in_data_187(pipe6_io_pipe_phv_in_data_187),
    .io_pipe_phv_in_data_188(pipe6_io_pipe_phv_in_data_188),
    .io_pipe_phv_in_data_189(pipe6_io_pipe_phv_in_data_189),
    .io_pipe_phv_in_data_190(pipe6_io_pipe_phv_in_data_190),
    .io_pipe_phv_in_data_191(pipe6_io_pipe_phv_in_data_191),
    .io_pipe_phv_in_data_192(pipe6_io_pipe_phv_in_data_192),
    .io_pipe_phv_in_data_193(pipe6_io_pipe_phv_in_data_193),
    .io_pipe_phv_in_data_194(pipe6_io_pipe_phv_in_data_194),
    .io_pipe_phv_in_data_195(pipe6_io_pipe_phv_in_data_195),
    .io_pipe_phv_in_data_196(pipe6_io_pipe_phv_in_data_196),
    .io_pipe_phv_in_data_197(pipe6_io_pipe_phv_in_data_197),
    .io_pipe_phv_in_data_198(pipe6_io_pipe_phv_in_data_198),
    .io_pipe_phv_in_data_199(pipe6_io_pipe_phv_in_data_199),
    .io_pipe_phv_in_data_200(pipe6_io_pipe_phv_in_data_200),
    .io_pipe_phv_in_data_201(pipe6_io_pipe_phv_in_data_201),
    .io_pipe_phv_in_data_202(pipe6_io_pipe_phv_in_data_202),
    .io_pipe_phv_in_data_203(pipe6_io_pipe_phv_in_data_203),
    .io_pipe_phv_in_data_204(pipe6_io_pipe_phv_in_data_204),
    .io_pipe_phv_in_data_205(pipe6_io_pipe_phv_in_data_205),
    .io_pipe_phv_in_data_206(pipe6_io_pipe_phv_in_data_206),
    .io_pipe_phv_in_data_207(pipe6_io_pipe_phv_in_data_207),
    .io_pipe_phv_in_data_208(pipe6_io_pipe_phv_in_data_208),
    .io_pipe_phv_in_data_209(pipe6_io_pipe_phv_in_data_209),
    .io_pipe_phv_in_data_210(pipe6_io_pipe_phv_in_data_210),
    .io_pipe_phv_in_data_211(pipe6_io_pipe_phv_in_data_211),
    .io_pipe_phv_in_data_212(pipe6_io_pipe_phv_in_data_212),
    .io_pipe_phv_in_data_213(pipe6_io_pipe_phv_in_data_213),
    .io_pipe_phv_in_data_214(pipe6_io_pipe_phv_in_data_214),
    .io_pipe_phv_in_data_215(pipe6_io_pipe_phv_in_data_215),
    .io_pipe_phv_in_data_216(pipe6_io_pipe_phv_in_data_216),
    .io_pipe_phv_in_data_217(pipe6_io_pipe_phv_in_data_217),
    .io_pipe_phv_in_data_218(pipe6_io_pipe_phv_in_data_218),
    .io_pipe_phv_in_data_219(pipe6_io_pipe_phv_in_data_219),
    .io_pipe_phv_in_data_220(pipe6_io_pipe_phv_in_data_220),
    .io_pipe_phv_in_data_221(pipe6_io_pipe_phv_in_data_221),
    .io_pipe_phv_in_data_222(pipe6_io_pipe_phv_in_data_222),
    .io_pipe_phv_in_data_223(pipe6_io_pipe_phv_in_data_223),
    .io_pipe_phv_in_data_224(pipe6_io_pipe_phv_in_data_224),
    .io_pipe_phv_in_data_225(pipe6_io_pipe_phv_in_data_225),
    .io_pipe_phv_in_data_226(pipe6_io_pipe_phv_in_data_226),
    .io_pipe_phv_in_data_227(pipe6_io_pipe_phv_in_data_227),
    .io_pipe_phv_in_data_228(pipe6_io_pipe_phv_in_data_228),
    .io_pipe_phv_in_data_229(pipe6_io_pipe_phv_in_data_229),
    .io_pipe_phv_in_data_230(pipe6_io_pipe_phv_in_data_230),
    .io_pipe_phv_in_data_231(pipe6_io_pipe_phv_in_data_231),
    .io_pipe_phv_in_data_232(pipe6_io_pipe_phv_in_data_232),
    .io_pipe_phv_in_data_233(pipe6_io_pipe_phv_in_data_233),
    .io_pipe_phv_in_data_234(pipe6_io_pipe_phv_in_data_234),
    .io_pipe_phv_in_data_235(pipe6_io_pipe_phv_in_data_235),
    .io_pipe_phv_in_data_236(pipe6_io_pipe_phv_in_data_236),
    .io_pipe_phv_in_data_237(pipe6_io_pipe_phv_in_data_237),
    .io_pipe_phv_in_data_238(pipe6_io_pipe_phv_in_data_238),
    .io_pipe_phv_in_data_239(pipe6_io_pipe_phv_in_data_239),
    .io_pipe_phv_in_data_240(pipe6_io_pipe_phv_in_data_240),
    .io_pipe_phv_in_data_241(pipe6_io_pipe_phv_in_data_241),
    .io_pipe_phv_in_data_242(pipe6_io_pipe_phv_in_data_242),
    .io_pipe_phv_in_data_243(pipe6_io_pipe_phv_in_data_243),
    .io_pipe_phv_in_data_244(pipe6_io_pipe_phv_in_data_244),
    .io_pipe_phv_in_data_245(pipe6_io_pipe_phv_in_data_245),
    .io_pipe_phv_in_data_246(pipe6_io_pipe_phv_in_data_246),
    .io_pipe_phv_in_data_247(pipe6_io_pipe_phv_in_data_247),
    .io_pipe_phv_in_data_248(pipe6_io_pipe_phv_in_data_248),
    .io_pipe_phv_in_data_249(pipe6_io_pipe_phv_in_data_249),
    .io_pipe_phv_in_data_250(pipe6_io_pipe_phv_in_data_250),
    .io_pipe_phv_in_data_251(pipe6_io_pipe_phv_in_data_251),
    .io_pipe_phv_in_data_252(pipe6_io_pipe_phv_in_data_252),
    .io_pipe_phv_in_data_253(pipe6_io_pipe_phv_in_data_253),
    .io_pipe_phv_in_data_254(pipe6_io_pipe_phv_in_data_254),
    .io_pipe_phv_in_data_255(pipe6_io_pipe_phv_in_data_255),
    .io_pipe_phv_in_data_256(pipe6_io_pipe_phv_in_data_256),
    .io_pipe_phv_in_data_257(pipe6_io_pipe_phv_in_data_257),
    .io_pipe_phv_in_data_258(pipe6_io_pipe_phv_in_data_258),
    .io_pipe_phv_in_data_259(pipe6_io_pipe_phv_in_data_259),
    .io_pipe_phv_in_data_260(pipe6_io_pipe_phv_in_data_260),
    .io_pipe_phv_in_data_261(pipe6_io_pipe_phv_in_data_261),
    .io_pipe_phv_in_data_262(pipe6_io_pipe_phv_in_data_262),
    .io_pipe_phv_in_data_263(pipe6_io_pipe_phv_in_data_263),
    .io_pipe_phv_in_data_264(pipe6_io_pipe_phv_in_data_264),
    .io_pipe_phv_in_data_265(pipe6_io_pipe_phv_in_data_265),
    .io_pipe_phv_in_data_266(pipe6_io_pipe_phv_in_data_266),
    .io_pipe_phv_in_data_267(pipe6_io_pipe_phv_in_data_267),
    .io_pipe_phv_in_data_268(pipe6_io_pipe_phv_in_data_268),
    .io_pipe_phv_in_data_269(pipe6_io_pipe_phv_in_data_269),
    .io_pipe_phv_in_data_270(pipe6_io_pipe_phv_in_data_270),
    .io_pipe_phv_in_data_271(pipe6_io_pipe_phv_in_data_271),
    .io_pipe_phv_in_data_272(pipe6_io_pipe_phv_in_data_272),
    .io_pipe_phv_in_data_273(pipe6_io_pipe_phv_in_data_273),
    .io_pipe_phv_in_data_274(pipe6_io_pipe_phv_in_data_274),
    .io_pipe_phv_in_data_275(pipe6_io_pipe_phv_in_data_275),
    .io_pipe_phv_in_data_276(pipe6_io_pipe_phv_in_data_276),
    .io_pipe_phv_in_data_277(pipe6_io_pipe_phv_in_data_277),
    .io_pipe_phv_in_data_278(pipe6_io_pipe_phv_in_data_278),
    .io_pipe_phv_in_data_279(pipe6_io_pipe_phv_in_data_279),
    .io_pipe_phv_in_data_280(pipe6_io_pipe_phv_in_data_280),
    .io_pipe_phv_in_data_281(pipe6_io_pipe_phv_in_data_281),
    .io_pipe_phv_in_data_282(pipe6_io_pipe_phv_in_data_282),
    .io_pipe_phv_in_data_283(pipe6_io_pipe_phv_in_data_283),
    .io_pipe_phv_in_data_284(pipe6_io_pipe_phv_in_data_284),
    .io_pipe_phv_in_data_285(pipe6_io_pipe_phv_in_data_285),
    .io_pipe_phv_in_data_286(pipe6_io_pipe_phv_in_data_286),
    .io_pipe_phv_in_data_287(pipe6_io_pipe_phv_in_data_287),
    .io_pipe_phv_in_data_288(pipe6_io_pipe_phv_in_data_288),
    .io_pipe_phv_in_data_289(pipe6_io_pipe_phv_in_data_289),
    .io_pipe_phv_in_data_290(pipe6_io_pipe_phv_in_data_290),
    .io_pipe_phv_in_data_291(pipe6_io_pipe_phv_in_data_291),
    .io_pipe_phv_in_data_292(pipe6_io_pipe_phv_in_data_292),
    .io_pipe_phv_in_data_293(pipe6_io_pipe_phv_in_data_293),
    .io_pipe_phv_in_data_294(pipe6_io_pipe_phv_in_data_294),
    .io_pipe_phv_in_data_295(pipe6_io_pipe_phv_in_data_295),
    .io_pipe_phv_in_data_296(pipe6_io_pipe_phv_in_data_296),
    .io_pipe_phv_in_data_297(pipe6_io_pipe_phv_in_data_297),
    .io_pipe_phv_in_data_298(pipe6_io_pipe_phv_in_data_298),
    .io_pipe_phv_in_data_299(pipe6_io_pipe_phv_in_data_299),
    .io_pipe_phv_in_data_300(pipe6_io_pipe_phv_in_data_300),
    .io_pipe_phv_in_data_301(pipe6_io_pipe_phv_in_data_301),
    .io_pipe_phv_in_data_302(pipe6_io_pipe_phv_in_data_302),
    .io_pipe_phv_in_data_303(pipe6_io_pipe_phv_in_data_303),
    .io_pipe_phv_in_data_304(pipe6_io_pipe_phv_in_data_304),
    .io_pipe_phv_in_data_305(pipe6_io_pipe_phv_in_data_305),
    .io_pipe_phv_in_data_306(pipe6_io_pipe_phv_in_data_306),
    .io_pipe_phv_in_data_307(pipe6_io_pipe_phv_in_data_307),
    .io_pipe_phv_in_data_308(pipe6_io_pipe_phv_in_data_308),
    .io_pipe_phv_in_data_309(pipe6_io_pipe_phv_in_data_309),
    .io_pipe_phv_in_data_310(pipe6_io_pipe_phv_in_data_310),
    .io_pipe_phv_in_data_311(pipe6_io_pipe_phv_in_data_311),
    .io_pipe_phv_in_data_312(pipe6_io_pipe_phv_in_data_312),
    .io_pipe_phv_in_data_313(pipe6_io_pipe_phv_in_data_313),
    .io_pipe_phv_in_data_314(pipe6_io_pipe_phv_in_data_314),
    .io_pipe_phv_in_data_315(pipe6_io_pipe_phv_in_data_315),
    .io_pipe_phv_in_data_316(pipe6_io_pipe_phv_in_data_316),
    .io_pipe_phv_in_data_317(pipe6_io_pipe_phv_in_data_317),
    .io_pipe_phv_in_data_318(pipe6_io_pipe_phv_in_data_318),
    .io_pipe_phv_in_data_319(pipe6_io_pipe_phv_in_data_319),
    .io_pipe_phv_in_data_320(pipe6_io_pipe_phv_in_data_320),
    .io_pipe_phv_in_data_321(pipe6_io_pipe_phv_in_data_321),
    .io_pipe_phv_in_data_322(pipe6_io_pipe_phv_in_data_322),
    .io_pipe_phv_in_data_323(pipe6_io_pipe_phv_in_data_323),
    .io_pipe_phv_in_data_324(pipe6_io_pipe_phv_in_data_324),
    .io_pipe_phv_in_data_325(pipe6_io_pipe_phv_in_data_325),
    .io_pipe_phv_in_data_326(pipe6_io_pipe_phv_in_data_326),
    .io_pipe_phv_in_data_327(pipe6_io_pipe_phv_in_data_327),
    .io_pipe_phv_in_data_328(pipe6_io_pipe_phv_in_data_328),
    .io_pipe_phv_in_data_329(pipe6_io_pipe_phv_in_data_329),
    .io_pipe_phv_in_data_330(pipe6_io_pipe_phv_in_data_330),
    .io_pipe_phv_in_data_331(pipe6_io_pipe_phv_in_data_331),
    .io_pipe_phv_in_data_332(pipe6_io_pipe_phv_in_data_332),
    .io_pipe_phv_in_data_333(pipe6_io_pipe_phv_in_data_333),
    .io_pipe_phv_in_data_334(pipe6_io_pipe_phv_in_data_334),
    .io_pipe_phv_in_data_335(pipe6_io_pipe_phv_in_data_335),
    .io_pipe_phv_in_data_336(pipe6_io_pipe_phv_in_data_336),
    .io_pipe_phv_in_data_337(pipe6_io_pipe_phv_in_data_337),
    .io_pipe_phv_in_data_338(pipe6_io_pipe_phv_in_data_338),
    .io_pipe_phv_in_data_339(pipe6_io_pipe_phv_in_data_339),
    .io_pipe_phv_in_data_340(pipe6_io_pipe_phv_in_data_340),
    .io_pipe_phv_in_data_341(pipe6_io_pipe_phv_in_data_341),
    .io_pipe_phv_in_data_342(pipe6_io_pipe_phv_in_data_342),
    .io_pipe_phv_in_data_343(pipe6_io_pipe_phv_in_data_343),
    .io_pipe_phv_in_data_344(pipe6_io_pipe_phv_in_data_344),
    .io_pipe_phv_in_data_345(pipe6_io_pipe_phv_in_data_345),
    .io_pipe_phv_in_data_346(pipe6_io_pipe_phv_in_data_346),
    .io_pipe_phv_in_data_347(pipe6_io_pipe_phv_in_data_347),
    .io_pipe_phv_in_data_348(pipe6_io_pipe_phv_in_data_348),
    .io_pipe_phv_in_data_349(pipe6_io_pipe_phv_in_data_349),
    .io_pipe_phv_in_data_350(pipe6_io_pipe_phv_in_data_350),
    .io_pipe_phv_in_data_351(pipe6_io_pipe_phv_in_data_351),
    .io_pipe_phv_in_data_352(pipe6_io_pipe_phv_in_data_352),
    .io_pipe_phv_in_data_353(pipe6_io_pipe_phv_in_data_353),
    .io_pipe_phv_in_data_354(pipe6_io_pipe_phv_in_data_354),
    .io_pipe_phv_in_data_355(pipe6_io_pipe_phv_in_data_355),
    .io_pipe_phv_in_data_356(pipe6_io_pipe_phv_in_data_356),
    .io_pipe_phv_in_data_357(pipe6_io_pipe_phv_in_data_357),
    .io_pipe_phv_in_data_358(pipe6_io_pipe_phv_in_data_358),
    .io_pipe_phv_in_data_359(pipe6_io_pipe_phv_in_data_359),
    .io_pipe_phv_in_data_360(pipe6_io_pipe_phv_in_data_360),
    .io_pipe_phv_in_data_361(pipe6_io_pipe_phv_in_data_361),
    .io_pipe_phv_in_data_362(pipe6_io_pipe_phv_in_data_362),
    .io_pipe_phv_in_data_363(pipe6_io_pipe_phv_in_data_363),
    .io_pipe_phv_in_data_364(pipe6_io_pipe_phv_in_data_364),
    .io_pipe_phv_in_data_365(pipe6_io_pipe_phv_in_data_365),
    .io_pipe_phv_in_data_366(pipe6_io_pipe_phv_in_data_366),
    .io_pipe_phv_in_data_367(pipe6_io_pipe_phv_in_data_367),
    .io_pipe_phv_in_data_368(pipe6_io_pipe_phv_in_data_368),
    .io_pipe_phv_in_data_369(pipe6_io_pipe_phv_in_data_369),
    .io_pipe_phv_in_data_370(pipe6_io_pipe_phv_in_data_370),
    .io_pipe_phv_in_data_371(pipe6_io_pipe_phv_in_data_371),
    .io_pipe_phv_in_data_372(pipe6_io_pipe_phv_in_data_372),
    .io_pipe_phv_in_data_373(pipe6_io_pipe_phv_in_data_373),
    .io_pipe_phv_in_data_374(pipe6_io_pipe_phv_in_data_374),
    .io_pipe_phv_in_data_375(pipe6_io_pipe_phv_in_data_375),
    .io_pipe_phv_in_data_376(pipe6_io_pipe_phv_in_data_376),
    .io_pipe_phv_in_data_377(pipe6_io_pipe_phv_in_data_377),
    .io_pipe_phv_in_data_378(pipe6_io_pipe_phv_in_data_378),
    .io_pipe_phv_in_data_379(pipe6_io_pipe_phv_in_data_379),
    .io_pipe_phv_in_data_380(pipe6_io_pipe_phv_in_data_380),
    .io_pipe_phv_in_data_381(pipe6_io_pipe_phv_in_data_381),
    .io_pipe_phv_in_data_382(pipe6_io_pipe_phv_in_data_382),
    .io_pipe_phv_in_data_383(pipe6_io_pipe_phv_in_data_383),
    .io_pipe_phv_in_data_384(pipe6_io_pipe_phv_in_data_384),
    .io_pipe_phv_in_data_385(pipe6_io_pipe_phv_in_data_385),
    .io_pipe_phv_in_data_386(pipe6_io_pipe_phv_in_data_386),
    .io_pipe_phv_in_data_387(pipe6_io_pipe_phv_in_data_387),
    .io_pipe_phv_in_data_388(pipe6_io_pipe_phv_in_data_388),
    .io_pipe_phv_in_data_389(pipe6_io_pipe_phv_in_data_389),
    .io_pipe_phv_in_data_390(pipe6_io_pipe_phv_in_data_390),
    .io_pipe_phv_in_data_391(pipe6_io_pipe_phv_in_data_391),
    .io_pipe_phv_in_data_392(pipe6_io_pipe_phv_in_data_392),
    .io_pipe_phv_in_data_393(pipe6_io_pipe_phv_in_data_393),
    .io_pipe_phv_in_data_394(pipe6_io_pipe_phv_in_data_394),
    .io_pipe_phv_in_data_395(pipe6_io_pipe_phv_in_data_395),
    .io_pipe_phv_in_data_396(pipe6_io_pipe_phv_in_data_396),
    .io_pipe_phv_in_data_397(pipe6_io_pipe_phv_in_data_397),
    .io_pipe_phv_in_data_398(pipe6_io_pipe_phv_in_data_398),
    .io_pipe_phv_in_data_399(pipe6_io_pipe_phv_in_data_399),
    .io_pipe_phv_in_data_400(pipe6_io_pipe_phv_in_data_400),
    .io_pipe_phv_in_data_401(pipe6_io_pipe_phv_in_data_401),
    .io_pipe_phv_in_data_402(pipe6_io_pipe_phv_in_data_402),
    .io_pipe_phv_in_data_403(pipe6_io_pipe_phv_in_data_403),
    .io_pipe_phv_in_data_404(pipe6_io_pipe_phv_in_data_404),
    .io_pipe_phv_in_data_405(pipe6_io_pipe_phv_in_data_405),
    .io_pipe_phv_in_data_406(pipe6_io_pipe_phv_in_data_406),
    .io_pipe_phv_in_data_407(pipe6_io_pipe_phv_in_data_407),
    .io_pipe_phv_in_data_408(pipe6_io_pipe_phv_in_data_408),
    .io_pipe_phv_in_data_409(pipe6_io_pipe_phv_in_data_409),
    .io_pipe_phv_in_data_410(pipe6_io_pipe_phv_in_data_410),
    .io_pipe_phv_in_data_411(pipe6_io_pipe_phv_in_data_411),
    .io_pipe_phv_in_data_412(pipe6_io_pipe_phv_in_data_412),
    .io_pipe_phv_in_data_413(pipe6_io_pipe_phv_in_data_413),
    .io_pipe_phv_in_data_414(pipe6_io_pipe_phv_in_data_414),
    .io_pipe_phv_in_data_415(pipe6_io_pipe_phv_in_data_415),
    .io_pipe_phv_in_data_416(pipe6_io_pipe_phv_in_data_416),
    .io_pipe_phv_in_data_417(pipe6_io_pipe_phv_in_data_417),
    .io_pipe_phv_in_data_418(pipe6_io_pipe_phv_in_data_418),
    .io_pipe_phv_in_data_419(pipe6_io_pipe_phv_in_data_419),
    .io_pipe_phv_in_data_420(pipe6_io_pipe_phv_in_data_420),
    .io_pipe_phv_in_data_421(pipe6_io_pipe_phv_in_data_421),
    .io_pipe_phv_in_data_422(pipe6_io_pipe_phv_in_data_422),
    .io_pipe_phv_in_data_423(pipe6_io_pipe_phv_in_data_423),
    .io_pipe_phv_in_data_424(pipe6_io_pipe_phv_in_data_424),
    .io_pipe_phv_in_data_425(pipe6_io_pipe_phv_in_data_425),
    .io_pipe_phv_in_data_426(pipe6_io_pipe_phv_in_data_426),
    .io_pipe_phv_in_data_427(pipe6_io_pipe_phv_in_data_427),
    .io_pipe_phv_in_data_428(pipe6_io_pipe_phv_in_data_428),
    .io_pipe_phv_in_data_429(pipe6_io_pipe_phv_in_data_429),
    .io_pipe_phv_in_data_430(pipe6_io_pipe_phv_in_data_430),
    .io_pipe_phv_in_data_431(pipe6_io_pipe_phv_in_data_431),
    .io_pipe_phv_in_data_432(pipe6_io_pipe_phv_in_data_432),
    .io_pipe_phv_in_data_433(pipe6_io_pipe_phv_in_data_433),
    .io_pipe_phv_in_data_434(pipe6_io_pipe_phv_in_data_434),
    .io_pipe_phv_in_data_435(pipe6_io_pipe_phv_in_data_435),
    .io_pipe_phv_in_data_436(pipe6_io_pipe_phv_in_data_436),
    .io_pipe_phv_in_data_437(pipe6_io_pipe_phv_in_data_437),
    .io_pipe_phv_in_data_438(pipe6_io_pipe_phv_in_data_438),
    .io_pipe_phv_in_data_439(pipe6_io_pipe_phv_in_data_439),
    .io_pipe_phv_in_data_440(pipe6_io_pipe_phv_in_data_440),
    .io_pipe_phv_in_data_441(pipe6_io_pipe_phv_in_data_441),
    .io_pipe_phv_in_data_442(pipe6_io_pipe_phv_in_data_442),
    .io_pipe_phv_in_data_443(pipe6_io_pipe_phv_in_data_443),
    .io_pipe_phv_in_data_444(pipe6_io_pipe_phv_in_data_444),
    .io_pipe_phv_in_data_445(pipe6_io_pipe_phv_in_data_445),
    .io_pipe_phv_in_data_446(pipe6_io_pipe_phv_in_data_446),
    .io_pipe_phv_in_data_447(pipe6_io_pipe_phv_in_data_447),
    .io_pipe_phv_in_data_448(pipe6_io_pipe_phv_in_data_448),
    .io_pipe_phv_in_data_449(pipe6_io_pipe_phv_in_data_449),
    .io_pipe_phv_in_data_450(pipe6_io_pipe_phv_in_data_450),
    .io_pipe_phv_in_data_451(pipe6_io_pipe_phv_in_data_451),
    .io_pipe_phv_in_data_452(pipe6_io_pipe_phv_in_data_452),
    .io_pipe_phv_in_data_453(pipe6_io_pipe_phv_in_data_453),
    .io_pipe_phv_in_data_454(pipe6_io_pipe_phv_in_data_454),
    .io_pipe_phv_in_data_455(pipe6_io_pipe_phv_in_data_455),
    .io_pipe_phv_in_data_456(pipe6_io_pipe_phv_in_data_456),
    .io_pipe_phv_in_data_457(pipe6_io_pipe_phv_in_data_457),
    .io_pipe_phv_in_data_458(pipe6_io_pipe_phv_in_data_458),
    .io_pipe_phv_in_data_459(pipe6_io_pipe_phv_in_data_459),
    .io_pipe_phv_in_data_460(pipe6_io_pipe_phv_in_data_460),
    .io_pipe_phv_in_data_461(pipe6_io_pipe_phv_in_data_461),
    .io_pipe_phv_in_data_462(pipe6_io_pipe_phv_in_data_462),
    .io_pipe_phv_in_data_463(pipe6_io_pipe_phv_in_data_463),
    .io_pipe_phv_in_data_464(pipe6_io_pipe_phv_in_data_464),
    .io_pipe_phv_in_data_465(pipe6_io_pipe_phv_in_data_465),
    .io_pipe_phv_in_data_466(pipe6_io_pipe_phv_in_data_466),
    .io_pipe_phv_in_data_467(pipe6_io_pipe_phv_in_data_467),
    .io_pipe_phv_in_data_468(pipe6_io_pipe_phv_in_data_468),
    .io_pipe_phv_in_data_469(pipe6_io_pipe_phv_in_data_469),
    .io_pipe_phv_in_data_470(pipe6_io_pipe_phv_in_data_470),
    .io_pipe_phv_in_data_471(pipe6_io_pipe_phv_in_data_471),
    .io_pipe_phv_in_data_472(pipe6_io_pipe_phv_in_data_472),
    .io_pipe_phv_in_data_473(pipe6_io_pipe_phv_in_data_473),
    .io_pipe_phv_in_data_474(pipe6_io_pipe_phv_in_data_474),
    .io_pipe_phv_in_data_475(pipe6_io_pipe_phv_in_data_475),
    .io_pipe_phv_in_data_476(pipe6_io_pipe_phv_in_data_476),
    .io_pipe_phv_in_data_477(pipe6_io_pipe_phv_in_data_477),
    .io_pipe_phv_in_data_478(pipe6_io_pipe_phv_in_data_478),
    .io_pipe_phv_in_data_479(pipe6_io_pipe_phv_in_data_479),
    .io_pipe_phv_in_data_480(pipe6_io_pipe_phv_in_data_480),
    .io_pipe_phv_in_data_481(pipe6_io_pipe_phv_in_data_481),
    .io_pipe_phv_in_data_482(pipe6_io_pipe_phv_in_data_482),
    .io_pipe_phv_in_data_483(pipe6_io_pipe_phv_in_data_483),
    .io_pipe_phv_in_data_484(pipe6_io_pipe_phv_in_data_484),
    .io_pipe_phv_in_data_485(pipe6_io_pipe_phv_in_data_485),
    .io_pipe_phv_in_data_486(pipe6_io_pipe_phv_in_data_486),
    .io_pipe_phv_in_data_487(pipe6_io_pipe_phv_in_data_487),
    .io_pipe_phv_in_data_488(pipe6_io_pipe_phv_in_data_488),
    .io_pipe_phv_in_data_489(pipe6_io_pipe_phv_in_data_489),
    .io_pipe_phv_in_data_490(pipe6_io_pipe_phv_in_data_490),
    .io_pipe_phv_in_data_491(pipe6_io_pipe_phv_in_data_491),
    .io_pipe_phv_in_data_492(pipe6_io_pipe_phv_in_data_492),
    .io_pipe_phv_in_data_493(pipe6_io_pipe_phv_in_data_493),
    .io_pipe_phv_in_data_494(pipe6_io_pipe_phv_in_data_494),
    .io_pipe_phv_in_data_495(pipe6_io_pipe_phv_in_data_495),
    .io_pipe_phv_in_data_496(pipe6_io_pipe_phv_in_data_496),
    .io_pipe_phv_in_data_497(pipe6_io_pipe_phv_in_data_497),
    .io_pipe_phv_in_data_498(pipe6_io_pipe_phv_in_data_498),
    .io_pipe_phv_in_data_499(pipe6_io_pipe_phv_in_data_499),
    .io_pipe_phv_in_data_500(pipe6_io_pipe_phv_in_data_500),
    .io_pipe_phv_in_data_501(pipe6_io_pipe_phv_in_data_501),
    .io_pipe_phv_in_data_502(pipe6_io_pipe_phv_in_data_502),
    .io_pipe_phv_in_data_503(pipe6_io_pipe_phv_in_data_503),
    .io_pipe_phv_in_data_504(pipe6_io_pipe_phv_in_data_504),
    .io_pipe_phv_in_data_505(pipe6_io_pipe_phv_in_data_505),
    .io_pipe_phv_in_data_506(pipe6_io_pipe_phv_in_data_506),
    .io_pipe_phv_in_data_507(pipe6_io_pipe_phv_in_data_507),
    .io_pipe_phv_in_data_508(pipe6_io_pipe_phv_in_data_508),
    .io_pipe_phv_in_data_509(pipe6_io_pipe_phv_in_data_509),
    .io_pipe_phv_in_data_510(pipe6_io_pipe_phv_in_data_510),
    .io_pipe_phv_in_data_511(pipe6_io_pipe_phv_in_data_511),
    .io_pipe_phv_in_header_0(pipe6_io_pipe_phv_in_header_0),
    .io_pipe_phv_in_header_1(pipe6_io_pipe_phv_in_header_1),
    .io_pipe_phv_in_header_2(pipe6_io_pipe_phv_in_header_2),
    .io_pipe_phv_in_header_3(pipe6_io_pipe_phv_in_header_3),
    .io_pipe_phv_in_header_4(pipe6_io_pipe_phv_in_header_4),
    .io_pipe_phv_in_header_5(pipe6_io_pipe_phv_in_header_5),
    .io_pipe_phv_in_header_6(pipe6_io_pipe_phv_in_header_6),
    .io_pipe_phv_in_header_7(pipe6_io_pipe_phv_in_header_7),
    .io_pipe_phv_in_header_8(pipe6_io_pipe_phv_in_header_8),
    .io_pipe_phv_in_header_9(pipe6_io_pipe_phv_in_header_9),
    .io_pipe_phv_in_header_10(pipe6_io_pipe_phv_in_header_10),
    .io_pipe_phv_in_header_11(pipe6_io_pipe_phv_in_header_11),
    .io_pipe_phv_in_header_12(pipe6_io_pipe_phv_in_header_12),
    .io_pipe_phv_in_header_13(pipe6_io_pipe_phv_in_header_13),
    .io_pipe_phv_in_header_14(pipe6_io_pipe_phv_in_header_14),
    .io_pipe_phv_in_header_15(pipe6_io_pipe_phv_in_header_15),
    .io_pipe_phv_in_parse_current_state(pipe6_io_pipe_phv_in_parse_current_state),
    .io_pipe_phv_in_parse_current_offset(pipe6_io_pipe_phv_in_parse_current_offset),
    .io_pipe_phv_in_parse_transition_field(pipe6_io_pipe_phv_in_parse_transition_field),
    .io_pipe_phv_in_next_processor_id(pipe6_io_pipe_phv_in_next_processor_id),
    .io_pipe_phv_in_next_config_id(pipe6_io_pipe_phv_in_next_config_id),
    .io_pipe_phv_in_is_valid_processor(pipe6_io_pipe_phv_in_is_valid_processor),
    .io_pipe_phv_out_data_0(pipe6_io_pipe_phv_out_data_0),
    .io_pipe_phv_out_data_1(pipe6_io_pipe_phv_out_data_1),
    .io_pipe_phv_out_data_2(pipe6_io_pipe_phv_out_data_2),
    .io_pipe_phv_out_data_3(pipe6_io_pipe_phv_out_data_3),
    .io_pipe_phv_out_data_4(pipe6_io_pipe_phv_out_data_4),
    .io_pipe_phv_out_data_5(pipe6_io_pipe_phv_out_data_5),
    .io_pipe_phv_out_data_6(pipe6_io_pipe_phv_out_data_6),
    .io_pipe_phv_out_data_7(pipe6_io_pipe_phv_out_data_7),
    .io_pipe_phv_out_data_8(pipe6_io_pipe_phv_out_data_8),
    .io_pipe_phv_out_data_9(pipe6_io_pipe_phv_out_data_9),
    .io_pipe_phv_out_data_10(pipe6_io_pipe_phv_out_data_10),
    .io_pipe_phv_out_data_11(pipe6_io_pipe_phv_out_data_11),
    .io_pipe_phv_out_data_12(pipe6_io_pipe_phv_out_data_12),
    .io_pipe_phv_out_data_13(pipe6_io_pipe_phv_out_data_13),
    .io_pipe_phv_out_data_14(pipe6_io_pipe_phv_out_data_14),
    .io_pipe_phv_out_data_15(pipe6_io_pipe_phv_out_data_15),
    .io_pipe_phv_out_data_16(pipe6_io_pipe_phv_out_data_16),
    .io_pipe_phv_out_data_17(pipe6_io_pipe_phv_out_data_17),
    .io_pipe_phv_out_data_18(pipe6_io_pipe_phv_out_data_18),
    .io_pipe_phv_out_data_19(pipe6_io_pipe_phv_out_data_19),
    .io_pipe_phv_out_data_20(pipe6_io_pipe_phv_out_data_20),
    .io_pipe_phv_out_data_21(pipe6_io_pipe_phv_out_data_21),
    .io_pipe_phv_out_data_22(pipe6_io_pipe_phv_out_data_22),
    .io_pipe_phv_out_data_23(pipe6_io_pipe_phv_out_data_23),
    .io_pipe_phv_out_data_24(pipe6_io_pipe_phv_out_data_24),
    .io_pipe_phv_out_data_25(pipe6_io_pipe_phv_out_data_25),
    .io_pipe_phv_out_data_26(pipe6_io_pipe_phv_out_data_26),
    .io_pipe_phv_out_data_27(pipe6_io_pipe_phv_out_data_27),
    .io_pipe_phv_out_data_28(pipe6_io_pipe_phv_out_data_28),
    .io_pipe_phv_out_data_29(pipe6_io_pipe_phv_out_data_29),
    .io_pipe_phv_out_data_30(pipe6_io_pipe_phv_out_data_30),
    .io_pipe_phv_out_data_31(pipe6_io_pipe_phv_out_data_31),
    .io_pipe_phv_out_data_32(pipe6_io_pipe_phv_out_data_32),
    .io_pipe_phv_out_data_33(pipe6_io_pipe_phv_out_data_33),
    .io_pipe_phv_out_data_34(pipe6_io_pipe_phv_out_data_34),
    .io_pipe_phv_out_data_35(pipe6_io_pipe_phv_out_data_35),
    .io_pipe_phv_out_data_36(pipe6_io_pipe_phv_out_data_36),
    .io_pipe_phv_out_data_37(pipe6_io_pipe_phv_out_data_37),
    .io_pipe_phv_out_data_38(pipe6_io_pipe_phv_out_data_38),
    .io_pipe_phv_out_data_39(pipe6_io_pipe_phv_out_data_39),
    .io_pipe_phv_out_data_40(pipe6_io_pipe_phv_out_data_40),
    .io_pipe_phv_out_data_41(pipe6_io_pipe_phv_out_data_41),
    .io_pipe_phv_out_data_42(pipe6_io_pipe_phv_out_data_42),
    .io_pipe_phv_out_data_43(pipe6_io_pipe_phv_out_data_43),
    .io_pipe_phv_out_data_44(pipe6_io_pipe_phv_out_data_44),
    .io_pipe_phv_out_data_45(pipe6_io_pipe_phv_out_data_45),
    .io_pipe_phv_out_data_46(pipe6_io_pipe_phv_out_data_46),
    .io_pipe_phv_out_data_47(pipe6_io_pipe_phv_out_data_47),
    .io_pipe_phv_out_data_48(pipe6_io_pipe_phv_out_data_48),
    .io_pipe_phv_out_data_49(pipe6_io_pipe_phv_out_data_49),
    .io_pipe_phv_out_data_50(pipe6_io_pipe_phv_out_data_50),
    .io_pipe_phv_out_data_51(pipe6_io_pipe_phv_out_data_51),
    .io_pipe_phv_out_data_52(pipe6_io_pipe_phv_out_data_52),
    .io_pipe_phv_out_data_53(pipe6_io_pipe_phv_out_data_53),
    .io_pipe_phv_out_data_54(pipe6_io_pipe_phv_out_data_54),
    .io_pipe_phv_out_data_55(pipe6_io_pipe_phv_out_data_55),
    .io_pipe_phv_out_data_56(pipe6_io_pipe_phv_out_data_56),
    .io_pipe_phv_out_data_57(pipe6_io_pipe_phv_out_data_57),
    .io_pipe_phv_out_data_58(pipe6_io_pipe_phv_out_data_58),
    .io_pipe_phv_out_data_59(pipe6_io_pipe_phv_out_data_59),
    .io_pipe_phv_out_data_60(pipe6_io_pipe_phv_out_data_60),
    .io_pipe_phv_out_data_61(pipe6_io_pipe_phv_out_data_61),
    .io_pipe_phv_out_data_62(pipe6_io_pipe_phv_out_data_62),
    .io_pipe_phv_out_data_63(pipe6_io_pipe_phv_out_data_63),
    .io_pipe_phv_out_data_64(pipe6_io_pipe_phv_out_data_64),
    .io_pipe_phv_out_data_65(pipe6_io_pipe_phv_out_data_65),
    .io_pipe_phv_out_data_66(pipe6_io_pipe_phv_out_data_66),
    .io_pipe_phv_out_data_67(pipe6_io_pipe_phv_out_data_67),
    .io_pipe_phv_out_data_68(pipe6_io_pipe_phv_out_data_68),
    .io_pipe_phv_out_data_69(pipe6_io_pipe_phv_out_data_69),
    .io_pipe_phv_out_data_70(pipe6_io_pipe_phv_out_data_70),
    .io_pipe_phv_out_data_71(pipe6_io_pipe_phv_out_data_71),
    .io_pipe_phv_out_data_72(pipe6_io_pipe_phv_out_data_72),
    .io_pipe_phv_out_data_73(pipe6_io_pipe_phv_out_data_73),
    .io_pipe_phv_out_data_74(pipe6_io_pipe_phv_out_data_74),
    .io_pipe_phv_out_data_75(pipe6_io_pipe_phv_out_data_75),
    .io_pipe_phv_out_data_76(pipe6_io_pipe_phv_out_data_76),
    .io_pipe_phv_out_data_77(pipe6_io_pipe_phv_out_data_77),
    .io_pipe_phv_out_data_78(pipe6_io_pipe_phv_out_data_78),
    .io_pipe_phv_out_data_79(pipe6_io_pipe_phv_out_data_79),
    .io_pipe_phv_out_data_80(pipe6_io_pipe_phv_out_data_80),
    .io_pipe_phv_out_data_81(pipe6_io_pipe_phv_out_data_81),
    .io_pipe_phv_out_data_82(pipe6_io_pipe_phv_out_data_82),
    .io_pipe_phv_out_data_83(pipe6_io_pipe_phv_out_data_83),
    .io_pipe_phv_out_data_84(pipe6_io_pipe_phv_out_data_84),
    .io_pipe_phv_out_data_85(pipe6_io_pipe_phv_out_data_85),
    .io_pipe_phv_out_data_86(pipe6_io_pipe_phv_out_data_86),
    .io_pipe_phv_out_data_87(pipe6_io_pipe_phv_out_data_87),
    .io_pipe_phv_out_data_88(pipe6_io_pipe_phv_out_data_88),
    .io_pipe_phv_out_data_89(pipe6_io_pipe_phv_out_data_89),
    .io_pipe_phv_out_data_90(pipe6_io_pipe_phv_out_data_90),
    .io_pipe_phv_out_data_91(pipe6_io_pipe_phv_out_data_91),
    .io_pipe_phv_out_data_92(pipe6_io_pipe_phv_out_data_92),
    .io_pipe_phv_out_data_93(pipe6_io_pipe_phv_out_data_93),
    .io_pipe_phv_out_data_94(pipe6_io_pipe_phv_out_data_94),
    .io_pipe_phv_out_data_95(pipe6_io_pipe_phv_out_data_95),
    .io_pipe_phv_out_data_96(pipe6_io_pipe_phv_out_data_96),
    .io_pipe_phv_out_data_97(pipe6_io_pipe_phv_out_data_97),
    .io_pipe_phv_out_data_98(pipe6_io_pipe_phv_out_data_98),
    .io_pipe_phv_out_data_99(pipe6_io_pipe_phv_out_data_99),
    .io_pipe_phv_out_data_100(pipe6_io_pipe_phv_out_data_100),
    .io_pipe_phv_out_data_101(pipe6_io_pipe_phv_out_data_101),
    .io_pipe_phv_out_data_102(pipe6_io_pipe_phv_out_data_102),
    .io_pipe_phv_out_data_103(pipe6_io_pipe_phv_out_data_103),
    .io_pipe_phv_out_data_104(pipe6_io_pipe_phv_out_data_104),
    .io_pipe_phv_out_data_105(pipe6_io_pipe_phv_out_data_105),
    .io_pipe_phv_out_data_106(pipe6_io_pipe_phv_out_data_106),
    .io_pipe_phv_out_data_107(pipe6_io_pipe_phv_out_data_107),
    .io_pipe_phv_out_data_108(pipe6_io_pipe_phv_out_data_108),
    .io_pipe_phv_out_data_109(pipe6_io_pipe_phv_out_data_109),
    .io_pipe_phv_out_data_110(pipe6_io_pipe_phv_out_data_110),
    .io_pipe_phv_out_data_111(pipe6_io_pipe_phv_out_data_111),
    .io_pipe_phv_out_data_112(pipe6_io_pipe_phv_out_data_112),
    .io_pipe_phv_out_data_113(pipe6_io_pipe_phv_out_data_113),
    .io_pipe_phv_out_data_114(pipe6_io_pipe_phv_out_data_114),
    .io_pipe_phv_out_data_115(pipe6_io_pipe_phv_out_data_115),
    .io_pipe_phv_out_data_116(pipe6_io_pipe_phv_out_data_116),
    .io_pipe_phv_out_data_117(pipe6_io_pipe_phv_out_data_117),
    .io_pipe_phv_out_data_118(pipe6_io_pipe_phv_out_data_118),
    .io_pipe_phv_out_data_119(pipe6_io_pipe_phv_out_data_119),
    .io_pipe_phv_out_data_120(pipe6_io_pipe_phv_out_data_120),
    .io_pipe_phv_out_data_121(pipe6_io_pipe_phv_out_data_121),
    .io_pipe_phv_out_data_122(pipe6_io_pipe_phv_out_data_122),
    .io_pipe_phv_out_data_123(pipe6_io_pipe_phv_out_data_123),
    .io_pipe_phv_out_data_124(pipe6_io_pipe_phv_out_data_124),
    .io_pipe_phv_out_data_125(pipe6_io_pipe_phv_out_data_125),
    .io_pipe_phv_out_data_126(pipe6_io_pipe_phv_out_data_126),
    .io_pipe_phv_out_data_127(pipe6_io_pipe_phv_out_data_127),
    .io_pipe_phv_out_data_128(pipe6_io_pipe_phv_out_data_128),
    .io_pipe_phv_out_data_129(pipe6_io_pipe_phv_out_data_129),
    .io_pipe_phv_out_data_130(pipe6_io_pipe_phv_out_data_130),
    .io_pipe_phv_out_data_131(pipe6_io_pipe_phv_out_data_131),
    .io_pipe_phv_out_data_132(pipe6_io_pipe_phv_out_data_132),
    .io_pipe_phv_out_data_133(pipe6_io_pipe_phv_out_data_133),
    .io_pipe_phv_out_data_134(pipe6_io_pipe_phv_out_data_134),
    .io_pipe_phv_out_data_135(pipe6_io_pipe_phv_out_data_135),
    .io_pipe_phv_out_data_136(pipe6_io_pipe_phv_out_data_136),
    .io_pipe_phv_out_data_137(pipe6_io_pipe_phv_out_data_137),
    .io_pipe_phv_out_data_138(pipe6_io_pipe_phv_out_data_138),
    .io_pipe_phv_out_data_139(pipe6_io_pipe_phv_out_data_139),
    .io_pipe_phv_out_data_140(pipe6_io_pipe_phv_out_data_140),
    .io_pipe_phv_out_data_141(pipe6_io_pipe_phv_out_data_141),
    .io_pipe_phv_out_data_142(pipe6_io_pipe_phv_out_data_142),
    .io_pipe_phv_out_data_143(pipe6_io_pipe_phv_out_data_143),
    .io_pipe_phv_out_data_144(pipe6_io_pipe_phv_out_data_144),
    .io_pipe_phv_out_data_145(pipe6_io_pipe_phv_out_data_145),
    .io_pipe_phv_out_data_146(pipe6_io_pipe_phv_out_data_146),
    .io_pipe_phv_out_data_147(pipe6_io_pipe_phv_out_data_147),
    .io_pipe_phv_out_data_148(pipe6_io_pipe_phv_out_data_148),
    .io_pipe_phv_out_data_149(pipe6_io_pipe_phv_out_data_149),
    .io_pipe_phv_out_data_150(pipe6_io_pipe_phv_out_data_150),
    .io_pipe_phv_out_data_151(pipe6_io_pipe_phv_out_data_151),
    .io_pipe_phv_out_data_152(pipe6_io_pipe_phv_out_data_152),
    .io_pipe_phv_out_data_153(pipe6_io_pipe_phv_out_data_153),
    .io_pipe_phv_out_data_154(pipe6_io_pipe_phv_out_data_154),
    .io_pipe_phv_out_data_155(pipe6_io_pipe_phv_out_data_155),
    .io_pipe_phv_out_data_156(pipe6_io_pipe_phv_out_data_156),
    .io_pipe_phv_out_data_157(pipe6_io_pipe_phv_out_data_157),
    .io_pipe_phv_out_data_158(pipe6_io_pipe_phv_out_data_158),
    .io_pipe_phv_out_data_159(pipe6_io_pipe_phv_out_data_159),
    .io_pipe_phv_out_data_160(pipe6_io_pipe_phv_out_data_160),
    .io_pipe_phv_out_data_161(pipe6_io_pipe_phv_out_data_161),
    .io_pipe_phv_out_data_162(pipe6_io_pipe_phv_out_data_162),
    .io_pipe_phv_out_data_163(pipe6_io_pipe_phv_out_data_163),
    .io_pipe_phv_out_data_164(pipe6_io_pipe_phv_out_data_164),
    .io_pipe_phv_out_data_165(pipe6_io_pipe_phv_out_data_165),
    .io_pipe_phv_out_data_166(pipe6_io_pipe_phv_out_data_166),
    .io_pipe_phv_out_data_167(pipe6_io_pipe_phv_out_data_167),
    .io_pipe_phv_out_data_168(pipe6_io_pipe_phv_out_data_168),
    .io_pipe_phv_out_data_169(pipe6_io_pipe_phv_out_data_169),
    .io_pipe_phv_out_data_170(pipe6_io_pipe_phv_out_data_170),
    .io_pipe_phv_out_data_171(pipe6_io_pipe_phv_out_data_171),
    .io_pipe_phv_out_data_172(pipe6_io_pipe_phv_out_data_172),
    .io_pipe_phv_out_data_173(pipe6_io_pipe_phv_out_data_173),
    .io_pipe_phv_out_data_174(pipe6_io_pipe_phv_out_data_174),
    .io_pipe_phv_out_data_175(pipe6_io_pipe_phv_out_data_175),
    .io_pipe_phv_out_data_176(pipe6_io_pipe_phv_out_data_176),
    .io_pipe_phv_out_data_177(pipe6_io_pipe_phv_out_data_177),
    .io_pipe_phv_out_data_178(pipe6_io_pipe_phv_out_data_178),
    .io_pipe_phv_out_data_179(pipe6_io_pipe_phv_out_data_179),
    .io_pipe_phv_out_data_180(pipe6_io_pipe_phv_out_data_180),
    .io_pipe_phv_out_data_181(pipe6_io_pipe_phv_out_data_181),
    .io_pipe_phv_out_data_182(pipe6_io_pipe_phv_out_data_182),
    .io_pipe_phv_out_data_183(pipe6_io_pipe_phv_out_data_183),
    .io_pipe_phv_out_data_184(pipe6_io_pipe_phv_out_data_184),
    .io_pipe_phv_out_data_185(pipe6_io_pipe_phv_out_data_185),
    .io_pipe_phv_out_data_186(pipe6_io_pipe_phv_out_data_186),
    .io_pipe_phv_out_data_187(pipe6_io_pipe_phv_out_data_187),
    .io_pipe_phv_out_data_188(pipe6_io_pipe_phv_out_data_188),
    .io_pipe_phv_out_data_189(pipe6_io_pipe_phv_out_data_189),
    .io_pipe_phv_out_data_190(pipe6_io_pipe_phv_out_data_190),
    .io_pipe_phv_out_data_191(pipe6_io_pipe_phv_out_data_191),
    .io_pipe_phv_out_data_192(pipe6_io_pipe_phv_out_data_192),
    .io_pipe_phv_out_data_193(pipe6_io_pipe_phv_out_data_193),
    .io_pipe_phv_out_data_194(pipe6_io_pipe_phv_out_data_194),
    .io_pipe_phv_out_data_195(pipe6_io_pipe_phv_out_data_195),
    .io_pipe_phv_out_data_196(pipe6_io_pipe_phv_out_data_196),
    .io_pipe_phv_out_data_197(pipe6_io_pipe_phv_out_data_197),
    .io_pipe_phv_out_data_198(pipe6_io_pipe_phv_out_data_198),
    .io_pipe_phv_out_data_199(pipe6_io_pipe_phv_out_data_199),
    .io_pipe_phv_out_data_200(pipe6_io_pipe_phv_out_data_200),
    .io_pipe_phv_out_data_201(pipe6_io_pipe_phv_out_data_201),
    .io_pipe_phv_out_data_202(pipe6_io_pipe_phv_out_data_202),
    .io_pipe_phv_out_data_203(pipe6_io_pipe_phv_out_data_203),
    .io_pipe_phv_out_data_204(pipe6_io_pipe_phv_out_data_204),
    .io_pipe_phv_out_data_205(pipe6_io_pipe_phv_out_data_205),
    .io_pipe_phv_out_data_206(pipe6_io_pipe_phv_out_data_206),
    .io_pipe_phv_out_data_207(pipe6_io_pipe_phv_out_data_207),
    .io_pipe_phv_out_data_208(pipe6_io_pipe_phv_out_data_208),
    .io_pipe_phv_out_data_209(pipe6_io_pipe_phv_out_data_209),
    .io_pipe_phv_out_data_210(pipe6_io_pipe_phv_out_data_210),
    .io_pipe_phv_out_data_211(pipe6_io_pipe_phv_out_data_211),
    .io_pipe_phv_out_data_212(pipe6_io_pipe_phv_out_data_212),
    .io_pipe_phv_out_data_213(pipe6_io_pipe_phv_out_data_213),
    .io_pipe_phv_out_data_214(pipe6_io_pipe_phv_out_data_214),
    .io_pipe_phv_out_data_215(pipe6_io_pipe_phv_out_data_215),
    .io_pipe_phv_out_data_216(pipe6_io_pipe_phv_out_data_216),
    .io_pipe_phv_out_data_217(pipe6_io_pipe_phv_out_data_217),
    .io_pipe_phv_out_data_218(pipe6_io_pipe_phv_out_data_218),
    .io_pipe_phv_out_data_219(pipe6_io_pipe_phv_out_data_219),
    .io_pipe_phv_out_data_220(pipe6_io_pipe_phv_out_data_220),
    .io_pipe_phv_out_data_221(pipe6_io_pipe_phv_out_data_221),
    .io_pipe_phv_out_data_222(pipe6_io_pipe_phv_out_data_222),
    .io_pipe_phv_out_data_223(pipe6_io_pipe_phv_out_data_223),
    .io_pipe_phv_out_data_224(pipe6_io_pipe_phv_out_data_224),
    .io_pipe_phv_out_data_225(pipe6_io_pipe_phv_out_data_225),
    .io_pipe_phv_out_data_226(pipe6_io_pipe_phv_out_data_226),
    .io_pipe_phv_out_data_227(pipe6_io_pipe_phv_out_data_227),
    .io_pipe_phv_out_data_228(pipe6_io_pipe_phv_out_data_228),
    .io_pipe_phv_out_data_229(pipe6_io_pipe_phv_out_data_229),
    .io_pipe_phv_out_data_230(pipe6_io_pipe_phv_out_data_230),
    .io_pipe_phv_out_data_231(pipe6_io_pipe_phv_out_data_231),
    .io_pipe_phv_out_data_232(pipe6_io_pipe_phv_out_data_232),
    .io_pipe_phv_out_data_233(pipe6_io_pipe_phv_out_data_233),
    .io_pipe_phv_out_data_234(pipe6_io_pipe_phv_out_data_234),
    .io_pipe_phv_out_data_235(pipe6_io_pipe_phv_out_data_235),
    .io_pipe_phv_out_data_236(pipe6_io_pipe_phv_out_data_236),
    .io_pipe_phv_out_data_237(pipe6_io_pipe_phv_out_data_237),
    .io_pipe_phv_out_data_238(pipe6_io_pipe_phv_out_data_238),
    .io_pipe_phv_out_data_239(pipe6_io_pipe_phv_out_data_239),
    .io_pipe_phv_out_data_240(pipe6_io_pipe_phv_out_data_240),
    .io_pipe_phv_out_data_241(pipe6_io_pipe_phv_out_data_241),
    .io_pipe_phv_out_data_242(pipe6_io_pipe_phv_out_data_242),
    .io_pipe_phv_out_data_243(pipe6_io_pipe_phv_out_data_243),
    .io_pipe_phv_out_data_244(pipe6_io_pipe_phv_out_data_244),
    .io_pipe_phv_out_data_245(pipe6_io_pipe_phv_out_data_245),
    .io_pipe_phv_out_data_246(pipe6_io_pipe_phv_out_data_246),
    .io_pipe_phv_out_data_247(pipe6_io_pipe_phv_out_data_247),
    .io_pipe_phv_out_data_248(pipe6_io_pipe_phv_out_data_248),
    .io_pipe_phv_out_data_249(pipe6_io_pipe_phv_out_data_249),
    .io_pipe_phv_out_data_250(pipe6_io_pipe_phv_out_data_250),
    .io_pipe_phv_out_data_251(pipe6_io_pipe_phv_out_data_251),
    .io_pipe_phv_out_data_252(pipe6_io_pipe_phv_out_data_252),
    .io_pipe_phv_out_data_253(pipe6_io_pipe_phv_out_data_253),
    .io_pipe_phv_out_data_254(pipe6_io_pipe_phv_out_data_254),
    .io_pipe_phv_out_data_255(pipe6_io_pipe_phv_out_data_255),
    .io_pipe_phv_out_data_256(pipe6_io_pipe_phv_out_data_256),
    .io_pipe_phv_out_data_257(pipe6_io_pipe_phv_out_data_257),
    .io_pipe_phv_out_data_258(pipe6_io_pipe_phv_out_data_258),
    .io_pipe_phv_out_data_259(pipe6_io_pipe_phv_out_data_259),
    .io_pipe_phv_out_data_260(pipe6_io_pipe_phv_out_data_260),
    .io_pipe_phv_out_data_261(pipe6_io_pipe_phv_out_data_261),
    .io_pipe_phv_out_data_262(pipe6_io_pipe_phv_out_data_262),
    .io_pipe_phv_out_data_263(pipe6_io_pipe_phv_out_data_263),
    .io_pipe_phv_out_data_264(pipe6_io_pipe_phv_out_data_264),
    .io_pipe_phv_out_data_265(pipe6_io_pipe_phv_out_data_265),
    .io_pipe_phv_out_data_266(pipe6_io_pipe_phv_out_data_266),
    .io_pipe_phv_out_data_267(pipe6_io_pipe_phv_out_data_267),
    .io_pipe_phv_out_data_268(pipe6_io_pipe_phv_out_data_268),
    .io_pipe_phv_out_data_269(pipe6_io_pipe_phv_out_data_269),
    .io_pipe_phv_out_data_270(pipe6_io_pipe_phv_out_data_270),
    .io_pipe_phv_out_data_271(pipe6_io_pipe_phv_out_data_271),
    .io_pipe_phv_out_data_272(pipe6_io_pipe_phv_out_data_272),
    .io_pipe_phv_out_data_273(pipe6_io_pipe_phv_out_data_273),
    .io_pipe_phv_out_data_274(pipe6_io_pipe_phv_out_data_274),
    .io_pipe_phv_out_data_275(pipe6_io_pipe_phv_out_data_275),
    .io_pipe_phv_out_data_276(pipe6_io_pipe_phv_out_data_276),
    .io_pipe_phv_out_data_277(pipe6_io_pipe_phv_out_data_277),
    .io_pipe_phv_out_data_278(pipe6_io_pipe_phv_out_data_278),
    .io_pipe_phv_out_data_279(pipe6_io_pipe_phv_out_data_279),
    .io_pipe_phv_out_data_280(pipe6_io_pipe_phv_out_data_280),
    .io_pipe_phv_out_data_281(pipe6_io_pipe_phv_out_data_281),
    .io_pipe_phv_out_data_282(pipe6_io_pipe_phv_out_data_282),
    .io_pipe_phv_out_data_283(pipe6_io_pipe_phv_out_data_283),
    .io_pipe_phv_out_data_284(pipe6_io_pipe_phv_out_data_284),
    .io_pipe_phv_out_data_285(pipe6_io_pipe_phv_out_data_285),
    .io_pipe_phv_out_data_286(pipe6_io_pipe_phv_out_data_286),
    .io_pipe_phv_out_data_287(pipe6_io_pipe_phv_out_data_287),
    .io_pipe_phv_out_data_288(pipe6_io_pipe_phv_out_data_288),
    .io_pipe_phv_out_data_289(pipe6_io_pipe_phv_out_data_289),
    .io_pipe_phv_out_data_290(pipe6_io_pipe_phv_out_data_290),
    .io_pipe_phv_out_data_291(pipe6_io_pipe_phv_out_data_291),
    .io_pipe_phv_out_data_292(pipe6_io_pipe_phv_out_data_292),
    .io_pipe_phv_out_data_293(pipe6_io_pipe_phv_out_data_293),
    .io_pipe_phv_out_data_294(pipe6_io_pipe_phv_out_data_294),
    .io_pipe_phv_out_data_295(pipe6_io_pipe_phv_out_data_295),
    .io_pipe_phv_out_data_296(pipe6_io_pipe_phv_out_data_296),
    .io_pipe_phv_out_data_297(pipe6_io_pipe_phv_out_data_297),
    .io_pipe_phv_out_data_298(pipe6_io_pipe_phv_out_data_298),
    .io_pipe_phv_out_data_299(pipe6_io_pipe_phv_out_data_299),
    .io_pipe_phv_out_data_300(pipe6_io_pipe_phv_out_data_300),
    .io_pipe_phv_out_data_301(pipe6_io_pipe_phv_out_data_301),
    .io_pipe_phv_out_data_302(pipe6_io_pipe_phv_out_data_302),
    .io_pipe_phv_out_data_303(pipe6_io_pipe_phv_out_data_303),
    .io_pipe_phv_out_data_304(pipe6_io_pipe_phv_out_data_304),
    .io_pipe_phv_out_data_305(pipe6_io_pipe_phv_out_data_305),
    .io_pipe_phv_out_data_306(pipe6_io_pipe_phv_out_data_306),
    .io_pipe_phv_out_data_307(pipe6_io_pipe_phv_out_data_307),
    .io_pipe_phv_out_data_308(pipe6_io_pipe_phv_out_data_308),
    .io_pipe_phv_out_data_309(pipe6_io_pipe_phv_out_data_309),
    .io_pipe_phv_out_data_310(pipe6_io_pipe_phv_out_data_310),
    .io_pipe_phv_out_data_311(pipe6_io_pipe_phv_out_data_311),
    .io_pipe_phv_out_data_312(pipe6_io_pipe_phv_out_data_312),
    .io_pipe_phv_out_data_313(pipe6_io_pipe_phv_out_data_313),
    .io_pipe_phv_out_data_314(pipe6_io_pipe_phv_out_data_314),
    .io_pipe_phv_out_data_315(pipe6_io_pipe_phv_out_data_315),
    .io_pipe_phv_out_data_316(pipe6_io_pipe_phv_out_data_316),
    .io_pipe_phv_out_data_317(pipe6_io_pipe_phv_out_data_317),
    .io_pipe_phv_out_data_318(pipe6_io_pipe_phv_out_data_318),
    .io_pipe_phv_out_data_319(pipe6_io_pipe_phv_out_data_319),
    .io_pipe_phv_out_data_320(pipe6_io_pipe_phv_out_data_320),
    .io_pipe_phv_out_data_321(pipe6_io_pipe_phv_out_data_321),
    .io_pipe_phv_out_data_322(pipe6_io_pipe_phv_out_data_322),
    .io_pipe_phv_out_data_323(pipe6_io_pipe_phv_out_data_323),
    .io_pipe_phv_out_data_324(pipe6_io_pipe_phv_out_data_324),
    .io_pipe_phv_out_data_325(pipe6_io_pipe_phv_out_data_325),
    .io_pipe_phv_out_data_326(pipe6_io_pipe_phv_out_data_326),
    .io_pipe_phv_out_data_327(pipe6_io_pipe_phv_out_data_327),
    .io_pipe_phv_out_data_328(pipe6_io_pipe_phv_out_data_328),
    .io_pipe_phv_out_data_329(pipe6_io_pipe_phv_out_data_329),
    .io_pipe_phv_out_data_330(pipe6_io_pipe_phv_out_data_330),
    .io_pipe_phv_out_data_331(pipe6_io_pipe_phv_out_data_331),
    .io_pipe_phv_out_data_332(pipe6_io_pipe_phv_out_data_332),
    .io_pipe_phv_out_data_333(pipe6_io_pipe_phv_out_data_333),
    .io_pipe_phv_out_data_334(pipe6_io_pipe_phv_out_data_334),
    .io_pipe_phv_out_data_335(pipe6_io_pipe_phv_out_data_335),
    .io_pipe_phv_out_data_336(pipe6_io_pipe_phv_out_data_336),
    .io_pipe_phv_out_data_337(pipe6_io_pipe_phv_out_data_337),
    .io_pipe_phv_out_data_338(pipe6_io_pipe_phv_out_data_338),
    .io_pipe_phv_out_data_339(pipe6_io_pipe_phv_out_data_339),
    .io_pipe_phv_out_data_340(pipe6_io_pipe_phv_out_data_340),
    .io_pipe_phv_out_data_341(pipe6_io_pipe_phv_out_data_341),
    .io_pipe_phv_out_data_342(pipe6_io_pipe_phv_out_data_342),
    .io_pipe_phv_out_data_343(pipe6_io_pipe_phv_out_data_343),
    .io_pipe_phv_out_data_344(pipe6_io_pipe_phv_out_data_344),
    .io_pipe_phv_out_data_345(pipe6_io_pipe_phv_out_data_345),
    .io_pipe_phv_out_data_346(pipe6_io_pipe_phv_out_data_346),
    .io_pipe_phv_out_data_347(pipe6_io_pipe_phv_out_data_347),
    .io_pipe_phv_out_data_348(pipe6_io_pipe_phv_out_data_348),
    .io_pipe_phv_out_data_349(pipe6_io_pipe_phv_out_data_349),
    .io_pipe_phv_out_data_350(pipe6_io_pipe_phv_out_data_350),
    .io_pipe_phv_out_data_351(pipe6_io_pipe_phv_out_data_351),
    .io_pipe_phv_out_data_352(pipe6_io_pipe_phv_out_data_352),
    .io_pipe_phv_out_data_353(pipe6_io_pipe_phv_out_data_353),
    .io_pipe_phv_out_data_354(pipe6_io_pipe_phv_out_data_354),
    .io_pipe_phv_out_data_355(pipe6_io_pipe_phv_out_data_355),
    .io_pipe_phv_out_data_356(pipe6_io_pipe_phv_out_data_356),
    .io_pipe_phv_out_data_357(pipe6_io_pipe_phv_out_data_357),
    .io_pipe_phv_out_data_358(pipe6_io_pipe_phv_out_data_358),
    .io_pipe_phv_out_data_359(pipe6_io_pipe_phv_out_data_359),
    .io_pipe_phv_out_data_360(pipe6_io_pipe_phv_out_data_360),
    .io_pipe_phv_out_data_361(pipe6_io_pipe_phv_out_data_361),
    .io_pipe_phv_out_data_362(pipe6_io_pipe_phv_out_data_362),
    .io_pipe_phv_out_data_363(pipe6_io_pipe_phv_out_data_363),
    .io_pipe_phv_out_data_364(pipe6_io_pipe_phv_out_data_364),
    .io_pipe_phv_out_data_365(pipe6_io_pipe_phv_out_data_365),
    .io_pipe_phv_out_data_366(pipe6_io_pipe_phv_out_data_366),
    .io_pipe_phv_out_data_367(pipe6_io_pipe_phv_out_data_367),
    .io_pipe_phv_out_data_368(pipe6_io_pipe_phv_out_data_368),
    .io_pipe_phv_out_data_369(pipe6_io_pipe_phv_out_data_369),
    .io_pipe_phv_out_data_370(pipe6_io_pipe_phv_out_data_370),
    .io_pipe_phv_out_data_371(pipe6_io_pipe_phv_out_data_371),
    .io_pipe_phv_out_data_372(pipe6_io_pipe_phv_out_data_372),
    .io_pipe_phv_out_data_373(pipe6_io_pipe_phv_out_data_373),
    .io_pipe_phv_out_data_374(pipe6_io_pipe_phv_out_data_374),
    .io_pipe_phv_out_data_375(pipe6_io_pipe_phv_out_data_375),
    .io_pipe_phv_out_data_376(pipe6_io_pipe_phv_out_data_376),
    .io_pipe_phv_out_data_377(pipe6_io_pipe_phv_out_data_377),
    .io_pipe_phv_out_data_378(pipe6_io_pipe_phv_out_data_378),
    .io_pipe_phv_out_data_379(pipe6_io_pipe_phv_out_data_379),
    .io_pipe_phv_out_data_380(pipe6_io_pipe_phv_out_data_380),
    .io_pipe_phv_out_data_381(pipe6_io_pipe_phv_out_data_381),
    .io_pipe_phv_out_data_382(pipe6_io_pipe_phv_out_data_382),
    .io_pipe_phv_out_data_383(pipe6_io_pipe_phv_out_data_383),
    .io_pipe_phv_out_data_384(pipe6_io_pipe_phv_out_data_384),
    .io_pipe_phv_out_data_385(pipe6_io_pipe_phv_out_data_385),
    .io_pipe_phv_out_data_386(pipe6_io_pipe_phv_out_data_386),
    .io_pipe_phv_out_data_387(pipe6_io_pipe_phv_out_data_387),
    .io_pipe_phv_out_data_388(pipe6_io_pipe_phv_out_data_388),
    .io_pipe_phv_out_data_389(pipe6_io_pipe_phv_out_data_389),
    .io_pipe_phv_out_data_390(pipe6_io_pipe_phv_out_data_390),
    .io_pipe_phv_out_data_391(pipe6_io_pipe_phv_out_data_391),
    .io_pipe_phv_out_data_392(pipe6_io_pipe_phv_out_data_392),
    .io_pipe_phv_out_data_393(pipe6_io_pipe_phv_out_data_393),
    .io_pipe_phv_out_data_394(pipe6_io_pipe_phv_out_data_394),
    .io_pipe_phv_out_data_395(pipe6_io_pipe_phv_out_data_395),
    .io_pipe_phv_out_data_396(pipe6_io_pipe_phv_out_data_396),
    .io_pipe_phv_out_data_397(pipe6_io_pipe_phv_out_data_397),
    .io_pipe_phv_out_data_398(pipe6_io_pipe_phv_out_data_398),
    .io_pipe_phv_out_data_399(pipe6_io_pipe_phv_out_data_399),
    .io_pipe_phv_out_data_400(pipe6_io_pipe_phv_out_data_400),
    .io_pipe_phv_out_data_401(pipe6_io_pipe_phv_out_data_401),
    .io_pipe_phv_out_data_402(pipe6_io_pipe_phv_out_data_402),
    .io_pipe_phv_out_data_403(pipe6_io_pipe_phv_out_data_403),
    .io_pipe_phv_out_data_404(pipe6_io_pipe_phv_out_data_404),
    .io_pipe_phv_out_data_405(pipe6_io_pipe_phv_out_data_405),
    .io_pipe_phv_out_data_406(pipe6_io_pipe_phv_out_data_406),
    .io_pipe_phv_out_data_407(pipe6_io_pipe_phv_out_data_407),
    .io_pipe_phv_out_data_408(pipe6_io_pipe_phv_out_data_408),
    .io_pipe_phv_out_data_409(pipe6_io_pipe_phv_out_data_409),
    .io_pipe_phv_out_data_410(pipe6_io_pipe_phv_out_data_410),
    .io_pipe_phv_out_data_411(pipe6_io_pipe_phv_out_data_411),
    .io_pipe_phv_out_data_412(pipe6_io_pipe_phv_out_data_412),
    .io_pipe_phv_out_data_413(pipe6_io_pipe_phv_out_data_413),
    .io_pipe_phv_out_data_414(pipe6_io_pipe_phv_out_data_414),
    .io_pipe_phv_out_data_415(pipe6_io_pipe_phv_out_data_415),
    .io_pipe_phv_out_data_416(pipe6_io_pipe_phv_out_data_416),
    .io_pipe_phv_out_data_417(pipe6_io_pipe_phv_out_data_417),
    .io_pipe_phv_out_data_418(pipe6_io_pipe_phv_out_data_418),
    .io_pipe_phv_out_data_419(pipe6_io_pipe_phv_out_data_419),
    .io_pipe_phv_out_data_420(pipe6_io_pipe_phv_out_data_420),
    .io_pipe_phv_out_data_421(pipe6_io_pipe_phv_out_data_421),
    .io_pipe_phv_out_data_422(pipe6_io_pipe_phv_out_data_422),
    .io_pipe_phv_out_data_423(pipe6_io_pipe_phv_out_data_423),
    .io_pipe_phv_out_data_424(pipe6_io_pipe_phv_out_data_424),
    .io_pipe_phv_out_data_425(pipe6_io_pipe_phv_out_data_425),
    .io_pipe_phv_out_data_426(pipe6_io_pipe_phv_out_data_426),
    .io_pipe_phv_out_data_427(pipe6_io_pipe_phv_out_data_427),
    .io_pipe_phv_out_data_428(pipe6_io_pipe_phv_out_data_428),
    .io_pipe_phv_out_data_429(pipe6_io_pipe_phv_out_data_429),
    .io_pipe_phv_out_data_430(pipe6_io_pipe_phv_out_data_430),
    .io_pipe_phv_out_data_431(pipe6_io_pipe_phv_out_data_431),
    .io_pipe_phv_out_data_432(pipe6_io_pipe_phv_out_data_432),
    .io_pipe_phv_out_data_433(pipe6_io_pipe_phv_out_data_433),
    .io_pipe_phv_out_data_434(pipe6_io_pipe_phv_out_data_434),
    .io_pipe_phv_out_data_435(pipe6_io_pipe_phv_out_data_435),
    .io_pipe_phv_out_data_436(pipe6_io_pipe_phv_out_data_436),
    .io_pipe_phv_out_data_437(pipe6_io_pipe_phv_out_data_437),
    .io_pipe_phv_out_data_438(pipe6_io_pipe_phv_out_data_438),
    .io_pipe_phv_out_data_439(pipe6_io_pipe_phv_out_data_439),
    .io_pipe_phv_out_data_440(pipe6_io_pipe_phv_out_data_440),
    .io_pipe_phv_out_data_441(pipe6_io_pipe_phv_out_data_441),
    .io_pipe_phv_out_data_442(pipe6_io_pipe_phv_out_data_442),
    .io_pipe_phv_out_data_443(pipe6_io_pipe_phv_out_data_443),
    .io_pipe_phv_out_data_444(pipe6_io_pipe_phv_out_data_444),
    .io_pipe_phv_out_data_445(pipe6_io_pipe_phv_out_data_445),
    .io_pipe_phv_out_data_446(pipe6_io_pipe_phv_out_data_446),
    .io_pipe_phv_out_data_447(pipe6_io_pipe_phv_out_data_447),
    .io_pipe_phv_out_data_448(pipe6_io_pipe_phv_out_data_448),
    .io_pipe_phv_out_data_449(pipe6_io_pipe_phv_out_data_449),
    .io_pipe_phv_out_data_450(pipe6_io_pipe_phv_out_data_450),
    .io_pipe_phv_out_data_451(pipe6_io_pipe_phv_out_data_451),
    .io_pipe_phv_out_data_452(pipe6_io_pipe_phv_out_data_452),
    .io_pipe_phv_out_data_453(pipe6_io_pipe_phv_out_data_453),
    .io_pipe_phv_out_data_454(pipe6_io_pipe_phv_out_data_454),
    .io_pipe_phv_out_data_455(pipe6_io_pipe_phv_out_data_455),
    .io_pipe_phv_out_data_456(pipe6_io_pipe_phv_out_data_456),
    .io_pipe_phv_out_data_457(pipe6_io_pipe_phv_out_data_457),
    .io_pipe_phv_out_data_458(pipe6_io_pipe_phv_out_data_458),
    .io_pipe_phv_out_data_459(pipe6_io_pipe_phv_out_data_459),
    .io_pipe_phv_out_data_460(pipe6_io_pipe_phv_out_data_460),
    .io_pipe_phv_out_data_461(pipe6_io_pipe_phv_out_data_461),
    .io_pipe_phv_out_data_462(pipe6_io_pipe_phv_out_data_462),
    .io_pipe_phv_out_data_463(pipe6_io_pipe_phv_out_data_463),
    .io_pipe_phv_out_data_464(pipe6_io_pipe_phv_out_data_464),
    .io_pipe_phv_out_data_465(pipe6_io_pipe_phv_out_data_465),
    .io_pipe_phv_out_data_466(pipe6_io_pipe_phv_out_data_466),
    .io_pipe_phv_out_data_467(pipe6_io_pipe_phv_out_data_467),
    .io_pipe_phv_out_data_468(pipe6_io_pipe_phv_out_data_468),
    .io_pipe_phv_out_data_469(pipe6_io_pipe_phv_out_data_469),
    .io_pipe_phv_out_data_470(pipe6_io_pipe_phv_out_data_470),
    .io_pipe_phv_out_data_471(pipe6_io_pipe_phv_out_data_471),
    .io_pipe_phv_out_data_472(pipe6_io_pipe_phv_out_data_472),
    .io_pipe_phv_out_data_473(pipe6_io_pipe_phv_out_data_473),
    .io_pipe_phv_out_data_474(pipe6_io_pipe_phv_out_data_474),
    .io_pipe_phv_out_data_475(pipe6_io_pipe_phv_out_data_475),
    .io_pipe_phv_out_data_476(pipe6_io_pipe_phv_out_data_476),
    .io_pipe_phv_out_data_477(pipe6_io_pipe_phv_out_data_477),
    .io_pipe_phv_out_data_478(pipe6_io_pipe_phv_out_data_478),
    .io_pipe_phv_out_data_479(pipe6_io_pipe_phv_out_data_479),
    .io_pipe_phv_out_data_480(pipe6_io_pipe_phv_out_data_480),
    .io_pipe_phv_out_data_481(pipe6_io_pipe_phv_out_data_481),
    .io_pipe_phv_out_data_482(pipe6_io_pipe_phv_out_data_482),
    .io_pipe_phv_out_data_483(pipe6_io_pipe_phv_out_data_483),
    .io_pipe_phv_out_data_484(pipe6_io_pipe_phv_out_data_484),
    .io_pipe_phv_out_data_485(pipe6_io_pipe_phv_out_data_485),
    .io_pipe_phv_out_data_486(pipe6_io_pipe_phv_out_data_486),
    .io_pipe_phv_out_data_487(pipe6_io_pipe_phv_out_data_487),
    .io_pipe_phv_out_data_488(pipe6_io_pipe_phv_out_data_488),
    .io_pipe_phv_out_data_489(pipe6_io_pipe_phv_out_data_489),
    .io_pipe_phv_out_data_490(pipe6_io_pipe_phv_out_data_490),
    .io_pipe_phv_out_data_491(pipe6_io_pipe_phv_out_data_491),
    .io_pipe_phv_out_data_492(pipe6_io_pipe_phv_out_data_492),
    .io_pipe_phv_out_data_493(pipe6_io_pipe_phv_out_data_493),
    .io_pipe_phv_out_data_494(pipe6_io_pipe_phv_out_data_494),
    .io_pipe_phv_out_data_495(pipe6_io_pipe_phv_out_data_495),
    .io_pipe_phv_out_data_496(pipe6_io_pipe_phv_out_data_496),
    .io_pipe_phv_out_data_497(pipe6_io_pipe_phv_out_data_497),
    .io_pipe_phv_out_data_498(pipe6_io_pipe_phv_out_data_498),
    .io_pipe_phv_out_data_499(pipe6_io_pipe_phv_out_data_499),
    .io_pipe_phv_out_data_500(pipe6_io_pipe_phv_out_data_500),
    .io_pipe_phv_out_data_501(pipe6_io_pipe_phv_out_data_501),
    .io_pipe_phv_out_data_502(pipe6_io_pipe_phv_out_data_502),
    .io_pipe_phv_out_data_503(pipe6_io_pipe_phv_out_data_503),
    .io_pipe_phv_out_data_504(pipe6_io_pipe_phv_out_data_504),
    .io_pipe_phv_out_data_505(pipe6_io_pipe_phv_out_data_505),
    .io_pipe_phv_out_data_506(pipe6_io_pipe_phv_out_data_506),
    .io_pipe_phv_out_data_507(pipe6_io_pipe_phv_out_data_507),
    .io_pipe_phv_out_data_508(pipe6_io_pipe_phv_out_data_508),
    .io_pipe_phv_out_data_509(pipe6_io_pipe_phv_out_data_509),
    .io_pipe_phv_out_data_510(pipe6_io_pipe_phv_out_data_510),
    .io_pipe_phv_out_data_511(pipe6_io_pipe_phv_out_data_511),
    .io_pipe_phv_out_header_0(pipe6_io_pipe_phv_out_header_0),
    .io_pipe_phv_out_header_1(pipe6_io_pipe_phv_out_header_1),
    .io_pipe_phv_out_header_2(pipe6_io_pipe_phv_out_header_2),
    .io_pipe_phv_out_header_3(pipe6_io_pipe_phv_out_header_3),
    .io_pipe_phv_out_header_4(pipe6_io_pipe_phv_out_header_4),
    .io_pipe_phv_out_header_5(pipe6_io_pipe_phv_out_header_5),
    .io_pipe_phv_out_header_6(pipe6_io_pipe_phv_out_header_6),
    .io_pipe_phv_out_header_7(pipe6_io_pipe_phv_out_header_7),
    .io_pipe_phv_out_header_8(pipe6_io_pipe_phv_out_header_8),
    .io_pipe_phv_out_header_9(pipe6_io_pipe_phv_out_header_9),
    .io_pipe_phv_out_header_10(pipe6_io_pipe_phv_out_header_10),
    .io_pipe_phv_out_header_11(pipe6_io_pipe_phv_out_header_11),
    .io_pipe_phv_out_header_12(pipe6_io_pipe_phv_out_header_12),
    .io_pipe_phv_out_header_13(pipe6_io_pipe_phv_out_header_13),
    .io_pipe_phv_out_header_14(pipe6_io_pipe_phv_out_header_14),
    .io_pipe_phv_out_header_15(pipe6_io_pipe_phv_out_header_15),
    .io_pipe_phv_out_parse_current_state(pipe6_io_pipe_phv_out_parse_current_state),
    .io_pipe_phv_out_parse_current_offset(pipe6_io_pipe_phv_out_parse_current_offset),
    .io_pipe_phv_out_parse_transition_field(pipe6_io_pipe_phv_out_parse_transition_field),
    .io_pipe_phv_out_next_processor_id(pipe6_io_pipe_phv_out_next_processor_id),
    .io_pipe_phv_out_next_config_id(pipe6_io_pipe_phv_out_next_config_id),
    .io_vliw_in_0(pipe6_io_vliw_in_0),
    .io_vliw_in_1(pipe6_io_vliw_in_1),
    .io_vliw_in_2(pipe6_io_vliw_in_2),
    .io_vliw_in_3(pipe6_io_vliw_in_3),
    .io_field_in_0(pipe6_io_field_in_0),
    .io_field_in_1(pipe6_io_field_in_1),
    .io_field_in_2(pipe6_io_field_in_2),
    .io_field_in_3(pipe6_io_field_in_3),
    .io_mask_in_0(pipe6_io_mask_in_0),
    .io_mask_in_1(pipe6_io_mask_in_1),
    .io_mask_in_2(pipe6_io_mask_in_2),
    .io_mask_in_3(pipe6_io_mask_in_3),
    .io_dst_offset_in_0(pipe6_io_dst_offset_in_0),
    .io_dst_offset_in_1(pipe6_io_dst_offset_in_1),
    .io_dst_offset_in_2(pipe6_io_dst_offset_in_2),
    .io_dst_offset_in_3(pipe6_io_dst_offset_in_3)
  );
  assign io_pipe_phv_out_data_0 = pipe6_io_pipe_phv_out_data_0; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_1 = pipe6_io_pipe_phv_out_data_1; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_2 = pipe6_io_pipe_phv_out_data_2; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_3 = pipe6_io_pipe_phv_out_data_3; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_4 = pipe6_io_pipe_phv_out_data_4; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_5 = pipe6_io_pipe_phv_out_data_5; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_6 = pipe6_io_pipe_phv_out_data_6; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_7 = pipe6_io_pipe_phv_out_data_7; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_8 = pipe6_io_pipe_phv_out_data_8; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_9 = pipe6_io_pipe_phv_out_data_9; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_10 = pipe6_io_pipe_phv_out_data_10; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_11 = pipe6_io_pipe_phv_out_data_11; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_12 = pipe6_io_pipe_phv_out_data_12; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_13 = pipe6_io_pipe_phv_out_data_13; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_14 = pipe6_io_pipe_phv_out_data_14; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_15 = pipe6_io_pipe_phv_out_data_15; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_16 = pipe6_io_pipe_phv_out_data_16; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_17 = pipe6_io_pipe_phv_out_data_17; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_18 = pipe6_io_pipe_phv_out_data_18; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_19 = pipe6_io_pipe_phv_out_data_19; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_20 = pipe6_io_pipe_phv_out_data_20; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_21 = pipe6_io_pipe_phv_out_data_21; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_22 = pipe6_io_pipe_phv_out_data_22; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_23 = pipe6_io_pipe_phv_out_data_23; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_24 = pipe6_io_pipe_phv_out_data_24; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_25 = pipe6_io_pipe_phv_out_data_25; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_26 = pipe6_io_pipe_phv_out_data_26; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_27 = pipe6_io_pipe_phv_out_data_27; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_28 = pipe6_io_pipe_phv_out_data_28; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_29 = pipe6_io_pipe_phv_out_data_29; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_30 = pipe6_io_pipe_phv_out_data_30; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_31 = pipe6_io_pipe_phv_out_data_31; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_32 = pipe6_io_pipe_phv_out_data_32; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_33 = pipe6_io_pipe_phv_out_data_33; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_34 = pipe6_io_pipe_phv_out_data_34; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_35 = pipe6_io_pipe_phv_out_data_35; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_36 = pipe6_io_pipe_phv_out_data_36; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_37 = pipe6_io_pipe_phv_out_data_37; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_38 = pipe6_io_pipe_phv_out_data_38; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_39 = pipe6_io_pipe_phv_out_data_39; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_40 = pipe6_io_pipe_phv_out_data_40; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_41 = pipe6_io_pipe_phv_out_data_41; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_42 = pipe6_io_pipe_phv_out_data_42; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_43 = pipe6_io_pipe_phv_out_data_43; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_44 = pipe6_io_pipe_phv_out_data_44; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_45 = pipe6_io_pipe_phv_out_data_45; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_46 = pipe6_io_pipe_phv_out_data_46; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_47 = pipe6_io_pipe_phv_out_data_47; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_48 = pipe6_io_pipe_phv_out_data_48; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_49 = pipe6_io_pipe_phv_out_data_49; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_50 = pipe6_io_pipe_phv_out_data_50; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_51 = pipe6_io_pipe_phv_out_data_51; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_52 = pipe6_io_pipe_phv_out_data_52; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_53 = pipe6_io_pipe_phv_out_data_53; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_54 = pipe6_io_pipe_phv_out_data_54; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_55 = pipe6_io_pipe_phv_out_data_55; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_56 = pipe6_io_pipe_phv_out_data_56; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_57 = pipe6_io_pipe_phv_out_data_57; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_58 = pipe6_io_pipe_phv_out_data_58; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_59 = pipe6_io_pipe_phv_out_data_59; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_60 = pipe6_io_pipe_phv_out_data_60; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_61 = pipe6_io_pipe_phv_out_data_61; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_62 = pipe6_io_pipe_phv_out_data_62; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_63 = pipe6_io_pipe_phv_out_data_63; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_64 = pipe6_io_pipe_phv_out_data_64; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_65 = pipe6_io_pipe_phv_out_data_65; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_66 = pipe6_io_pipe_phv_out_data_66; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_67 = pipe6_io_pipe_phv_out_data_67; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_68 = pipe6_io_pipe_phv_out_data_68; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_69 = pipe6_io_pipe_phv_out_data_69; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_70 = pipe6_io_pipe_phv_out_data_70; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_71 = pipe6_io_pipe_phv_out_data_71; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_72 = pipe6_io_pipe_phv_out_data_72; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_73 = pipe6_io_pipe_phv_out_data_73; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_74 = pipe6_io_pipe_phv_out_data_74; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_75 = pipe6_io_pipe_phv_out_data_75; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_76 = pipe6_io_pipe_phv_out_data_76; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_77 = pipe6_io_pipe_phv_out_data_77; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_78 = pipe6_io_pipe_phv_out_data_78; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_79 = pipe6_io_pipe_phv_out_data_79; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_80 = pipe6_io_pipe_phv_out_data_80; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_81 = pipe6_io_pipe_phv_out_data_81; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_82 = pipe6_io_pipe_phv_out_data_82; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_83 = pipe6_io_pipe_phv_out_data_83; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_84 = pipe6_io_pipe_phv_out_data_84; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_85 = pipe6_io_pipe_phv_out_data_85; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_86 = pipe6_io_pipe_phv_out_data_86; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_87 = pipe6_io_pipe_phv_out_data_87; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_88 = pipe6_io_pipe_phv_out_data_88; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_89 = pipe6_io_pipe_phv_out_data_89; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_90 = pipe6_io_pipe_phv_out_data_90; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_91 = pipe6_io_pipe_phv_out_data_91; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_92 = pipe6_io_pipe_phv_out_data_92; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_93 = pipe6_io_pipe_phv_out_data_93; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_94 = pipe6_io_pipe_phv_out_data_94; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_95 = pipe6_io_pipe_phv_out_data_95; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_96 = pipe6_io_pipe_phv_out_data_96; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_97 = pipe6_io_pipe_phv_out_data_97; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_98 = pipe6_io_pipe_phv_out_data_98; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_99 = pipe6_io_pipe_phv_out_data_99; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_100 = pipe6_io_pipe_phv_out_data_100; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_101 = pipe6_io_pipe_phv_out_data_101; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_102 = pipe6_io_pipe_phv_out_data_102; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_103 = pipe6_io_pipe_phv_out_data_103; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_104 = pipe6_io_pipe_phv_out_data_104; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_105 = pipe6_io_pipe_phv_out_data_105; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_106 = pipe6_io_pipe_phv_out_data_106; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_107 = pipe6_io_pipe_phv_out_data_107; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_108 = pipe6_io_pipe_phv_out_data_108; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_109 = pipe6_io_pipe_phv_out_data_109; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_110 = pipe6_io_pipe_phv_out_data_110; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_111 = pipe6_io_pipe_phv_out_data_111; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_112 = pipe6_io_pipe_phv_out_data_112; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_113 = pipe6_io_pipe_phv_out_data_113; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_114 = pipe6_io_pipe_phv_out_data_114; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_115 = pipe6_io_pipe_phv_out_data_115; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_116 = pipe6_io_pipe_phv_out_data_116; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_117 = pipe6_io_pipe_phv_out_data_117; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_118 = pipe6_io_pipe_phv_out_data_118; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_119 = pipe6_io_pipe_phv_out_data_119; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_120 = pipe6_io_pipe_phv_out_data_120; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_121 = pipe6_io_pipe_phv_out_data_121; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_122 = pipe6_io_pipe_phv_out_data_122; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_123 = pipe6_io_pipe_phv_out_data_123; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_124 = pipe6_io_pipe_phv_out_data_124; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_125 = pipe6_io_pipe_phv_out_data_125; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_126 = pipe6_io_pipe_phv_out_data_126; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_127 = pipe6_io_pipe_phv_out_data_127; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_128 = pipe6_io_pipe_phv_out_data_128; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_129 = pipe6_io_pipe_phv_out_data_129; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_130 = pipe6_io_pipe_phv_out_data_130; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_131 = pipe6_io_pipe_phv_out_data_131; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_132 = pipe6_io_pipe_phv_out_data_132; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_133 = pipe6_io_pipe_phv_out_data_133; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_134 = pipe6_io_pipe_phv_out_data_134; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_135 = pipe6_io_pipe_phv_out_data_135; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_136 = pipe6_io_pipe_phv_out_data_136; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_137 = pipe6_io_pipe_phv_out_data_137; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_138 = pipe6_io_pipe_phv_out_data_138; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_139 = pipe6_io_pipe_phv_out_data_139; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_140 = pipe6_io_pipe_phv_out_data_140; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_141 = pipe6_io_pipe_phv_out_data_141; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_142 = pipe6_io_pipe_phv_out_data_142; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_143 = pipe6_io_pipe_phv_out_data_143; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_144 = pipe6_io_pipe_phv_out_data_144; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_145 = pipe6_io_pipe_phv_out_data_145; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_146 = pipe6_io_pipe_phv_out_data_146; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_147 = pipe6_io_pipe_phv_out_data_147; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_148 = pipe6_io_pipe_phv_out_data_148; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_149 = pipe6_io_pipe_phv_out_data_149; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_150 = pipe6_io_pipe_phv_out_data_150; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_151 = pipe6_io_pipe_phv_out_data_151; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_152 = pipe6_io_pipe_phv_out_data_152; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_153 = pipe6_io_pipe_phv_out_data_153; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_154 = pipe6_io_pipe_phv_out_data_154; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_155 = pipe6_io_pipe_phv_out_data_155; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_156 = pipe6_io_pipe_phv_out_data_156; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_157 = pipe6_io_pipe_phv_out_data_157; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_158 = pipe6_io_pipe_phv_out_data_158; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_159 = pipe6_io_pipe_phv_out_data_159; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_160 = pipe6_io_pipe_phv_out_data_160; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_161 = pipe6_io_pipe_phv_out_data_161; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_162 = pipe6_io_pipe_phv_out_data_162; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_163 = pipe6_io_pipe_phv_out_data_163; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_164 = pipe6_io_pipe_phv_out_data_164; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_165 = pipe6_io_pipe_phv_out_data_165; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_166 = pipe6_io_pipe_phv_out_data_166; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_167 = pipe6_io_pipe_phv_out_data_167; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_168 = pipe6_io_pipe_phv_out_data_168; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_169 = pipe6_io_pipe_phv_out_data_169; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_170 = pipe6_io_pipe_phv_out_data_170; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_171 = pipe6_io_pipe_phv_out_data_171; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_172 = pipe6_io_pipe_phv_out_data_172; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_173 = pipe6_io_pipe_phv_out_data_173; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_174 = pipe6_io_pipe_phv_out_data_174; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_175 = pipe6_io_pipe_phv_out_data_175; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_176 = pipe6_io_pipe_phv_out_data_176; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_177 = pipe6_io_pipe_phv_out_data_177; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_178 = pipe6_io_pipe_phv_out_data_178; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_179 = pipe6_io_pipe_phv_out_data_179; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_180 = pipe6_io_pipe_phv_out_data_180; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_181 = pipe6_io_pipe_phv_out_data_181; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_182 = pipe6_io_pipe_phv_out_data_182; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_183 = pipe6_io_pipe_phv_out_data_183; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_184 = pipe6_io_pipe_phv_out_data_184; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_185 = pipe6_io_pipe_phv_out_data_185; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_186 = pipe6_io_pipe_phv_out_data_186; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_187 = pipe6_io_pipe_phv_out_data_187; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_188 = pipe6_io_pipe_phv_out_data_188; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_189 = pipe6_io_pipe_phv_out_data_189; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_190 = pipe6_io_pipe_phv_out_data_190; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_191 = pipe6_io_pipe_phv_out_data_191; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_192 = pipe6_io_pipe_phv_out_data_192; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_193 = pipe6_io_pipe_phv_out_data_193; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_194 = pipe6_io_pipe_phv_out_data_194; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_195 = pipe6_io_pipe_phv_out_data_195; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_196 = pipe6_io_pipe_phv_out_data_196; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_197 = pipe6_io_pipe_phv_out_data_197; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_198 = pipe6_io_pipe_phv_out_data_198; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_199 = pipe6_io_pipe_phv_out_data_199; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_200 = pipe6_io_pipe_phv_out_data_200; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_201 = pipe6_io_pipe_phv_out_data_201; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_202 = pipe6_io_pipe_phv_out_data_202; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_203 = pipe6_io_pipe_phv_out_data_203; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_204 = pipe6_io_pipe_phv_out_data_204; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_205 = pipe6_io_pipe_phv_out_data_205; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_206 = pipe6_io_pipe_phv_out_data_206; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_207 = pipe6_io_pipe_phv_out_data_207; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_208 = pipe6_io_pipe_phv_out_data_208; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_209 = pipe6_io_pipe_phv_out_data_209; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_210 = pipe6_io_pipe_phv_out_data_210; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_211 = pipe6_io_pipe_phv_out_data_211; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_212 = pipe6_io_pipe_phv_out_data_212; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_213 = pipe6_io_pipe_phv_out_data_213; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_214 = pipe6_io_pipe_phv_out_data_214; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_215 = pipe6_io_pipe_phv_out_data_215; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_216 = pipe6_io_pipe_phv_out_data_216; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_217 = pipe6_io_pipe_phv_out_data_217; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_218 = pipe6_io_pipe_phv_out_data_218; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_219 = pipe6_io_pipe_phv_out_data_219; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_220 = pipe6_io_pipe_phv_out_data_220; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_221 = pipe6_io_pipe_phv_out_data_221; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_222 = pipe6_io_pipe_phv_out_data_222; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_223 = pipe6_io_pipe_phv_out_data_223; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_224 = pipe6_io_pipe_phv_out_data_224; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_225 = pipe6_io_pipe_phv_out_data_225; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_226 = pipe6_io_pipe_phv_out_data_226; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_227 = pipe6_io_pipe_phv_out_data_227; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_228 = pipe6_io_pipe_phv_out_data_228; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_229 = pipe6_io_pipe_phv_out_data_229; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_230 = pipe6_io_pipe_phv_out_data_230; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_231 = pipe6_io_pipe_phv_out_data_231; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_232 = pipe6_io_pipe_phv_out_data_232; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_233 = pipe6_io_pipe_phv_out_data_233; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_234 = pipe6_io_pipe_phv_out_data_234; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_235 = pipe6_io_pipe_phv_out_data_235; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_236 = pipe6_io_pipe_phv_out_data_236; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_237 = pipe6_io_pipe_phv_out_data_237; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_238 = pipe6_io_pipe_phv_out_data_238; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_239 = pipe6_io_pipe_phv_out_data_239; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_240 = pipe6_io_pipe_phv_out_data_240; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_241 = pipe6_io_pipe_phv_out_data_241; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_242 = pipe6_io_pipe_phv_out_data_242; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_243 = pipe6_io_pipe_phv_out_data_243; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_244 = pipe6_io_pipe_phv_out_data_244; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_245 = pipe6_io_pipe_phv_out_data_245; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_246 = pipe6_io_pipe_phv_out_data_246; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_247 = pipe6_io_pipe_phv_out_data_247; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_248 = pipe6_io_pipe_phv_out_data_248; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_249 = pipe6_io_pipe_phv_out_data_249; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_250 = pipe6_io_pipe_phv_out_data_250; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_251 = pipe6_io_pipe_phv_out_data_251; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_252 = pipe6_io_pipe_phv_out_data_252; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_253 = pipe6_io_pipe_phv_out_data_253; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_254 = pipe6_io_pipe_phv_out_data_254; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_255 = pipe6_io_pipe_phv_out_data_255; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_256 = pipe6_io_pipe_phv_out_data_256; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_257 = pipe6_io_pipe_phv_out_data_257; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_258 = pipe6_io_pipe_phv_out_data_258; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_259 = pipe6_io_pipe_phv_out_data_259; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_260 = pipe6_io_pipe_phv_out_data_260; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_261 = pipe6_io_pipe_phv_out_data_261; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_262 = pipe6_io_pipe_phv_out_data_262; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_263 = pipe6_io_pipe_phv_out_data_263; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_264 = pipe6_io_pipe_phv_out_data_264; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_265 = pipe6_io_pipe_phv_out_data_265; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_266 = pipe6_io_pipe_phv_out_data_266; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_267 = pipe6_io_pipe_phv_out_data_267; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_268 = pipe6_io_pipe_phv_out_data_268; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_269 = pipe6_io_pipe_phv_out_data_269; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_270 = pipe6_io_pipe_phv_out_data_270; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_271 = pipe6_io_pipe_phv_out_data_271; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_272 = pipe6_io_pipe_phv_out_data_272; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_273 = pipe6_io_pipe_phv_out_data_273; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_274 = pipe6_io_pipe_phv_out_data_274; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_275 = pipe6_io_pipe_phv_out_data_275; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_276 = pipe6_io_pipe_phv_out_data_276; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_277 = pipe6_io_pipe_phv_out_data_277; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_278 = pipe6_io_pipe_phv_out_data_278; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_279 = pipe6_io_pipe_phv_out_data_279; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_280 = pipe6_io_pipe_phv_out_data_280; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_281 = pipe6_io_pipe_phv_out_data_281; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_282 = pipe6_io_pipe_phv_out_data_282; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_283 = pipe6_io_pipe_phv_out_data_283; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_284 = pipe6_io_pipe_phv_out_data_284; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_285 = pipe6_io_pipe_phv_out_data_285; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_286 = pipe6_io_pipe_phv_out_data_286; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_287 = pipe6_io_pipe_phv_out_data_287; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_288 = pipe6_io_pipe_phv_out_data_288; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_289 = pipe6_io_pipe_phv_out_data_289; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_290 = pipe6_io_pipe_phv_out_data_290; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_291 = pipe6_io_pipe_phv_out_data_291; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_292 = pipe6_io_pipe_phv_out_data_292; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_293 = pipe6_io_pipe_phv_out_data_293; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_294 = pipe6_io_pipe_phv_out_data_294; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_295 = pipe6_io_pipe_phv_out_data_295; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_296 = pipe6_io_pipe_phv_out_data_296; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_297 = pipe6_io_pipe_phv_out_data_297; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_298 = pipe6_io_pipe_phv_out_data_298; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_299 = pipe6_io_pipe_phv_out_data_299; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_300 = pipe6_io_pipe_phv_out_data_300; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_301 = pipe6_io_pipe_phv_out_data_301; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_302 = pipe6_io_pipe_phv_out_data_302; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_303 = pipe6_io_pipe_phv_out_data_303; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_304 = pipe6_io_pipe_phv_out_data_304; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_305 = pipe6_io_pipe_phv_out_data_305; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_306 = pipe6_io_pipe_phv_out_data_306; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_307 = pipe6_io_pipe_phv_out_data_307; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_308 = pipe6_io_pipe_phv_out_data_308; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_309 = pipe6_io_pipe_phv_out_data_309; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_310 = pipe6_io_pipe_phv_out_data_310; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_311 = pipe6_io_pipe_phv_out_data_311; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_312 = pipe6_io_pipe_phv_out_data_312; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_313 = pipe6_io_pipe_phv_out_data_313; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_314 = pipe6_io_pipe_phv_out_data_314; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_315 = pipe6_io_pipe_phv_out_data_315; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_316 = pipe6_io_pipe_phv_out_data_316; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_317 = pipe6_io_pipe_phv_out_data_317; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_318 = pipe6_io_pipe_phv_out_data_318; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_319 = pipe6_io_pipe_phv_out_data_319; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_320 = pipe6_io_pipe_phv_out_data_320; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_321 = pipe6_io_pipe_phv_out_data_321; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_322 = pipe6_io_pipe_phv_out_data_322; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_323 = pipe6_io_pipe_phv_out_data_323; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_324 = pipe6_io_pipe_phv_out_data_324; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_325 = pipe6_io_pipe_phv_out_data_325; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_326 = pipe6_io_pipe_phv_out_data_326; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_327 = pipe6_io_pipe_phv_out_data_327; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_328 = pipe6_io_pipe_phv_out_data_328; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_329 = pipe6_io_pipe_phv_out_data_329; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_330 = pipe6_io_pipe_phv_out_data_330; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_331 = pipe6_io_pipe_phv_out_data_331; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_332 = pipe6_io_pipe_phv_out_data_332; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_333 = pipe6_io_pipe_phv_out_data_333; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_334 = pipe6_io_pipe_phv_out_data_334; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_335 = pipe6_io_pipe_phv_out_data_335; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_336 = pipe6_io_pipe_phv_out_data_336; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_337 = pipe6_io_pipe_phv_out_data_337; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_338 = pipe6_io_pipe_phv_out_data_338; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_339 = pipe6_io_pipe_phv_out_data_339; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_340 = pipe6_io_pipe_phv_out_data_340; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_341 = pipe6_io_pipe_phv_out_data_341; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_342 = pipe6_io_pipe_phv_out_data_342; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_343 = pipe6_io_pipe_phv_out_data_343; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_344 = pipe6_io_pipe_phv_out_data_344; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_345 = pipe6_io_pipe_phv_out_data_345; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_346 = pipe6_io_pipe_phv_out_data_346; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_347 = pipe6_io_pipe_phv_out_data_347; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_348 = pipe6_io_pipe_phv_out_data_348; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_349 = pipe6_io_pipe_phv_out_data_349; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_350 = pipe6_io_pipe_phv_out_data_350; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_351 = pipe6_io_pipe_phv_out_data_351; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_352 = pipe6_io_pipe_phv_out_data_352; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_353 = pipe6_io_pipe_phv_out_data_353; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_354 = pipe6_io_pipe_phv_out_data_354; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_355 = pipe6_io_pipe_phv_out_data_355; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_356 = pipe6_io_pipe_phv_out_data_356; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_357 = pipe6_io_pipe_phv_out_data_357; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_358 = pipe6_io_pipe_phv_out_data_358; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_359 = pipe6_io_pipe_phv_out_data_359; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_360 = pipe6_io_pipe_phv_out_data_360; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_361 = pipe6_io_pipe_phv_out_data_361; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_362 = pipe6_io_pipe_phv_out_data_362; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_363 = pipe6_io_pipe_phv_out_data_363; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_364 = pipe6_io_pipe_phv_out_data_364; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_365 = pipe6_io_pipe_phv_out_data_365; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_366 = pipe6_io_pipe_phv_out_data_366; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_367 = pipe6_io_pipe_phv_out_data_367; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_368 = pipe6_io_pipe_phv_out_data_368; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_369 = pipe6_io_pipe_phv_out_data_369; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_370 = pipe6_io_pipe_phv_out_data_370; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_371 = pipe6_io_pipe_phv_out_data_371; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_372 = pipe6_io_pipe_phv_out_data_372; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_373 = pipe6_io_pipe_phv_out_data_373; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_374 = pipe6_io_pipe_phv_out_data_374; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_375 = pipe6_io_pipe_phv_out_data_375; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_376 = pipe6_io_pipe_phv_out_data_376; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_377 = pipe6_io_pipe_phv_out_data_377; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_378 = pipe6_io_pipe_phv_out_data_378; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_379 = pipe6_io_pipe_phv_out_data_379; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_380 = pipe6_io_pipe_phv_out_data_380; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_381 = pipe6_io_pipe_phv_out_data_381; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_382 = pipe6_io_pipe_phv_out_data_382; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_383 = pipe6_io_pipe_phv_out_data_383; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_384 = pipe6_io_pipe_phv_out_data_384; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_385 = pipe6_io_pipe_phv_out_data_385; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_386 = pipe6_io_pipe_phv_out_data_386; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_387 = pipe6_io_pipe_phv_out_data_387; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_388 = pipe6_io_pipe_phv_out_data_388; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_389 = pipe6_io_pipe_phv_out_data_389; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_390 = pipe6_io_pipe_phv_out_data_390; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_391 = pipe6_io_pipe_phv_out_data_391; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_392 = pipe6_io_pipe_phv_out_data_392; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_393 = pipe6_io_pipe_phv_out_data_393; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_394 = pipe6_io_pipe_phv_out_data_394; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_395 = pipe6_io_pipe_phv_out_data_395; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_396 = pipe6_io_pipe_phv_out_data_396; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_397 = pipe6_io_pipe_phv_out_data_397; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_398 = pipe6_io_pipe_phv_out_data_398; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_399 = pipe6_io_pipe_phv_out_data_399; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_400 = pipe6_io_pipe_phv_out_data_400; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_401 = pipe6_io_pipe_phv_out_data_401; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_402 = pipe6_io_pipe_phv_out_data_402; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_403 = pipe6_io_pipe_phv_out_data_403; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_404 = pipe6_io_pipe_phv_out_data_404; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_405 = pipe6_io_pipe_phv_out_data_405; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_406 = pipe6_io_pipe_phv_out_data_406; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_407 = pipe6_io_pipe_phv_out_data_407; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_408 = pipe6_io_pipe_phv_out_data_408; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_409 = pipe6_io_pipe_phv_out_data_409; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_410 = pipe6_io_pipe_phv_out_data_410; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_411 = pipe6_io_pipe_phv_out_data_411; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_412 = pipe6_io_pipe_phv_out_data_412; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_413 = pipe6_io_pipe_phv_out_data_413; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_414 = pipe6_io_pipe_phv_out_data_414; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_415 = pipe6_io_pipe_phv_out_data_415; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_416 = pipe6_io_pipe_phv_out_data_416; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_417 = pipe6_io_pipe_phv_out_data_417; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_418 = pipe6_io_pipe_phv_out_data_418; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_419 = pipe6_io_pipe_phv_out_data_419; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_420 = pipe6_io_pipe_phv_out_data_420; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_421 = pipe6_io_pipe_phv_out_data_421; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_422 = pipe6_io_pipe_phv_out_data_422; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_423 = pipe6_io_pipe_phv_out_data_423; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_424 = pipe6_io_pipe_phv_out_data_424; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_425 = pipe6_io_pipe_phv_out_data_425; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_426 = pipe6_io_pipe_phv_out_data_426; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_427 = pipe6_io_pipe_phv_out_data_427; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_428 = pipe6_io_pipe_phv_out_data_428; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_429 = pipe6_io_pipe_phv_out_data_429; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_430 = pipe6_io_pipe_phv_out_data_430; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_431 = pipe6_io_pipe_phv_out_data_431; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_432 = pipe6_io_pipe_phv_out_data_432; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_433 = pipe6_io_pipe_phv_out_data_433; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_434 = pipe6_io_pipe_phv_out_data_434; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_435 = pipe6_io_pipe_phv_out_data_435; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_436 = pipe6_io_pipe_phv_out_data_436; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_437 = pipe6_io_pipe_phv_out_data_437; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_438 = pipe6_io_pipe_phv_out_data_438; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_439 = pipe6_io_pipe_phv_out_data_439; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_440 = pipe6_io_pipe_phv_out_data_440; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_441 = pipe6_io_pipe_phv_out_data_441; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_442 = pipe6_io_pipe_phv_out_data_442; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_443 = pipe6_io_pipe_phv_out_data_443; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_444 = pipe6_io_pipe_phv_out_data_444; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_445 = pipe6_io_pipe_phv_out_data_445; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_446 = pipe6_io_pipe_phv_out_data_446; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_447 = pipe6_io_pipe_phv_out_data_447; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_448 = pipe6_io_pipe_phv_out_data_448; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_449 = pipe6_io_pipe_phv_out_data_449; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_450 = pipe6_io_pipe_phv_out_data_450; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_451 = pipe6_io_pipe_phv_out_data_451; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_452 = pipe6_io_pipe_phv_out_data_452; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_453 = pipe6_io_pipe_phv_out_data_453; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_454 = pipe6_io_pipe_phv_out_data_454; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_455 = pipe6_io_pipe_phv_out_data_455; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_456 = pipe6_io_pipe_phv_out_data_456; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_457 = pipe6_io_pipe_phv_out_data_457; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_458 = pipe6_io_pipe_phv_out_data_458; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_459 = pipe6_io_pipe_phv_out_data_459; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_460 = pipe6_io_pipe_phv_out_data_460; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_461 = pipe6_io_pipe_phv_out_data_461; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_462 = pipe6_io_pipe_phv_out_data_462; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_463 = pipe6_io_pipe_phv_out_data_463; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_464 = pipe6_io_pipe_phv_out_data_464; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_465 = pipe6_io_pipe_phv_out_data_465; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_466 = pipe6_io_pipe_phv_out_data_466; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_467 = pipe6_io_pipe_phv_out_data_467; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_468 = pipe6_io_pipe_phv_out_data_468; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_469 = pipe6_io_pipe_phv_out_data_469; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_470 = pipe6_io_pipe_phv_out_data_470; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_471 = pipe6_io_pipe_phv_out_data_471; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_472 = pipe6_io_pipe_phv_out_data_472; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_473 = pipe6_io_pipe_phv_out_data_473; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_474 = pipe6_io_pipe_phv_out_data_474; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_475 = pipe6_io_pipe_phv_out_data_475; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_476 = pipe6_io_pipe_phv_out_data_476; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_477 = pipe6_io_pipe_phv_out_data_477; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_478 = pipe6_io_pipe_phv_out_data_478; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_479 = pipe6_io_pipe_phv_out_data_479; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_480 = pipe6_io_pipe_phv_out_data_480; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_481 = pipe6_io_pipe_phv_out_data_481; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_482 = pipe6_io_pipe_phv_out_data_482; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_483 = pipe6_io_pipe_phv_out_data_483; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_484 = pipe6_io_pipe_phv_out_data_484; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_485 = pipe6_io_pipe_phv_out_data_485; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_486 = pipe6_io_pipe_phv_out_data_486; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_487 = pipe6_io_pipe_phv_out_data_487; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_488 = pipe6_io_pipe_phv_out_data_488; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_489 = pipe6_io_pipe_phv_out_data_489; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_490 = pipe6_io_pipe_phv_out_data_490; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_491 = pipe6_io_pipe_phv_out_data_491; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_492 = pipe6_io_pipe_phv_out_data_492; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_493 = pipe6_io_pipe_phv_out_data_493; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_494 = pipe6_io_pipe_phv_out_data_494; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_495 = pipe6_io_pipe_phv_out_data_495; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_496 = pipe6_io_pipe_phv_out_data_496; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_497 = pipe6_io_pipe_phv_out_data_497; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_498 = pipe6_io_pipe_phv_out_data_498; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_499 = pipe6_io_pipe_phv_out_data_499; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_500 = pipe6_io_pipe_phv_out_data_500; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_501 = pipe6_io_pipe_phv_out_data_501; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_502 = pipe6_io_pipe_phv_out_data_502; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_503 = pipe6_io_pipe_phv_out_data_503; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_504 = pipe6_io_pipe_phv_out_data_504; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_505 = pipe6_io_pipe_phv_out_data_505; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_506 = pipe6_io_pipe_phv_out_data_506; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_507 = pipe6_io_pipe_phv_out_data_507; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_508 = pipe6_io_pipe_phv_out_data_508; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_509 = pipe6_io_pipe_phv_out_data_509; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_510 = pipe6_io_pipe_phv_out_data_510; // @[executor.scala 530:27]
  assign io_pipe_phv_out_data_511 = pipe6_io_pipe_phv_out_data_511; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_0 = pipe6_io_pipe_phv_out_header_0; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_1 = pipe6_io_pipe_phv_out_header_1; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_2 = pipe6_io_pipe_phv_out_header_2; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_3 = pipe6_io_pipe_phv_out_header_3; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_4 = pipe6_io_pipe_phv_out_header_4; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_5 = pipe6_io_pipe_phv_out_header_5; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_6 = pipe6_io_pipe_phv_out_header_6; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_7 = pipe6_io_pipe_phv_out_header_7; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_8 = pipe6_io_pipe_phv_out_header_8; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_9 = pipe6_io_pipe_phv_out_header_9; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_10 = pipe6_io_pipe_phv_out_header_10; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_11 = pipe6_io_pipe_phv_out_header_11; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_12 = pipe6_io_pipe_phv_out_header_12; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_13 = pipe6_io_pipe_phv_out_header_13; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_14 = pipe6_io_pipe_phv_out_header_14; // @[executor.scala 530:27]
  assign io_pipe_phv_out_header_15 = pipe6_io_pipe_phv_out_header_15; // @[executor.scala 530:27]
  assign io_pipe_phv_out_parse_current_state = pipe6_io_pipe_phv_out_parse_current_state; // @[executor.scala 530:27]
  assign io_pipe_phv_out_parse_current_offset = pipe6_io_pipe_phv_out_parse_current_offset; // @[executor.scala 530:27]
  assign io_pipe_phv_out_parse_transition_field = pipe6_io_pipe_phv_out_parse_transition_field; // @[executor.scala 530:27]
  assign io_pipe_phv_out_next_processor_id = pipe6_io_pipe_phv_out_next_processor_id; // @[executor.scala 530:27]
  assign io_pipe_phv_out_next_config_id = pipe6_io_pipe_phv_out_next_config_id; // @[executor.scala 530:27]
  assign pipe1_clock = clock;
  assign pipe1_io_pipe_phv_in_data_0 = io_pipe_phv_in_data_0; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_1 = io_pipe_phv_in_data_1; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_2 = io_pipe_phv_in_data_2; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_3 = io_pipe_phv_in_data_3; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_4 = io_pipe_phv_in_data_4; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_5 = io_pipe_phv_in_data_5; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_6 = io_pipe_phv_in_data_6; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_7 = io_pipe_phv_in_data_7; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_8 = io_pipe_phv_in_data_8; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_9 = io_pipe_phv_in_data_9; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_10 = io_pipe_phv_in_data_10; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_11 = io_pipe_phv_in_data_11; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_12 = io_pipe_phv_in_data_12; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_13 = io_pipe_phv_in_data_13; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_14 = io_pipe_phv_in_data_14; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_15 = io_pipe_phv_in_data_15; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_16 = io_pipe_phv_in_data_16; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_17 = io_pipe_phv_in_data_17; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_18 = io_pipe_phv_in_data_18; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_19 = io_pipe_phv_in_data_19; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_20 = io_pipe_phv_in_data_20; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_21 = io_pipe_phv_in_data_21; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_22 = io_pipe_phv_in_data_22; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_23 = io_pipe_phv_in_data_23; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_24 = io_pipe_phv_in_data_24; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_25 = io_pipe_phv_in_data_25; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_26 = io_pipe_phv_in_data_26; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_27 = io_pipe_phv_in_data_27; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_28 = io_pipe_phv_in_data_28; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_29 = io_pipe_phv_in_data_29; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_30 = io_pipe_phv_in_data_30; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_31 = io_pipe_phv_in_data_31; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_32 = io_pipe_phv_in_data_32; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_33 = io_pipe_phv_in_data_33; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_34 = io_pipe_phv_in_data_34; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_35 = io_pipe_phv_in_data_35; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_36 = io_pipe_phv_in_data_36; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_37 = io_pipe_phv_in_data_37; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_38 = io_pipe_phv_in_data_38; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_39 = io_pipe_phv_in_data_39; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_40 = io_pipe_phv_in_data_40; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_41 = io_pipe_phv_in_data_41; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_42 = io_pipe_phv_in_data_42; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_43 = io_pipe_phv_in_data_43; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_44 = io_pipe_phv_in_data_44; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_45 = io_pipe_phv_in_data_45; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_46 = io_pipe_phv_in_data_46; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_47 = io_pipe_phv_in_data_47; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_48 = io_pipe_phv_in_data_48; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_49 = io_pipe_phv_in_data_49; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_50 = io_pipe_phv_in_data_50; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_51 = io_pipe_phv_in_data_51; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_52 = io_pipe_phv_in_data_52; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_53 = io_pipe_phv_in_data_53; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_54 = io_pipe_phv_in_data_54; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_55 = io_pipe_phv_in_data_55; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_56 = io_pipe_phv_in_data_56; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_57 = io_pipe_phv_in_data_57; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_58 = io_pipe_phv_in_data_58; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_59 = io_pipe_phv_in_data_59; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_60 = io_pipe_phv_in_data_60; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_61 = io_pipe_phv_in_data_61; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_62 = io_pipe_phv_in_data_62; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_63 = io_pipe_phv_in_data_63; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_64 = io_pipe_phv_in_data_64; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_65 = io_pipe_phv_in_data_65; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_66 = io_pipe_phv_in_data_66; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_67 = io_pipe_phv_in_data_67; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_68 = io_pipe_phv_in_data_68; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_69 = io_pipe_phv_in_data_69; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_70 = io_pipe_phv_in_data_70; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_71 = io_pipe_phv_in_data_71; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_72 = io_pipe_phv_in_data_72; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_73 = io_pipe_phv_in_data_73; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_74 = io_pipe_phv_in_data_74; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_75 = io_pipe_phv_in_data_75; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_76 = io_pipe_phv_in_data_76; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_77 = io_pipe_phv_in_data_77; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_78 = io_pipe_phv_in_data_78; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_79 = io_pipe_phv_in_data_79; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_80 = io_pipe_phv_in_data_80; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_81 = io_pipe_phv_in_data_81; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_82 = io_pipe_phv_in_data_82; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_83 = io_pipe_phv_in_data_83; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_84 = io_pipe_phv_in_data_84; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_85 = io_pipe_phv_in_data_85; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_86 = io_pipe_phv_in_data_86; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_87 = io_pipe_phv_in_data_87; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_88 = io_pipe_phv_in_data_88; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_89 = io_pipe_phv_in_data_89; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_90 = io_pipe_phv_in_data_90; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_91 = io_pipe_phv_in_data_91; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_92 = io_pipe_phv_in_data_92; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_93 = io_pipe_phv_in_data_93; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_94 = io_pipe_phv_in_data_94; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_95 = io_pipe_phv_in_data_95; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_96 = io_pipe_phv_in_data_96; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_97 = io_pipe_phv_in_data_97; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_98 = io_pipe_phv_in_data_98; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_99 = io_pipe_phv_in_data_99; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_100 = io_pipe_phv_in_data_100; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_101 = io_pipe_phv_in_data_101; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_102 = io_pipe_phv_in_data_102; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_103 = io_pipe_phv_in_data_103; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_104 = io_pipe_phv_in_data_104; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_105 = io_pipe_phv_in_data_105; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_106 = io_pipe_phv_in_data_106; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_107 = io_pipe_phv_in_data_107; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_108 = io_pipe_phv_in_data_108; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_109 = io_pipe_phv_in_data_109; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_110 = io_pipe_phv_in_data_110; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_111 = io_pipe_phv_in_data_111; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_112 = io_pipe_phv_in_data_112; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_113 = io_pipe_phv_in_data_113; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_114 = io_pipe_phv_in_data_114; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_115 = io_pipe_phv_in_data_115; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_116 = io_pipe_phv_in_data_116; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_117 = io_pipe_phv_in_data_117; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_118 = io_pipe_phv_in_data_118; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_119 = io_pipe_phv_in_data_119; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_120 = io_pipe_phv_in_data_120; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_121 = io_pipe_phv_in_data_121; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_122 = io_pipe_phv_in_data_122; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_123 = io_pipe_phv_in_data_123; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_124 = io_pipe_phv_in_data_124; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_125 = io_pipe_phv_in_data_125; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_126 = io_pipe_phv_in_data_126; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_127 = io_pipe_phv_in_data_127; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_128 = io_pipe_phv_in_data_128; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_129 = io_pipe_phv_in_data_129; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_130 = io_pipe_phv_in_data_130; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_131 = io_pipe_phv_in_data_131; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_132 = io_pipe_phv_in_data_132; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_133 = io_pipe_phv_in_data_133; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_134 = io_pipe_phv_in_data_134; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_135 = io_pipe_phv_in_data_135; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_136 = io_pipe_phv_in_data_136; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_137 = io_pipe_phv_in_data_137; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_138 = io_pipe_phv_in_data_138; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_139 = io_pipe_phv_in_data_139; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_140 = io_pipe_phv_in_data_140; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_141 = io_pipe_phv_in_data_141; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_142 = io_pipe_phv_in_data_142; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_143 = io_pipe_phv_in_data_143; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_144 = io_pipe_phv_in_data_144; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_145 = io_pipe_phv_in_data_145; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_146 = io_pipe_phv_in_data_146; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_147 = io_pipe_phv_in_data_147; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_148 = io_pipe_phv_in_data_148; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_149 = io_pipe_phv_in_data_149; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_150 = io_pipe_phv_in_data_150; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_151 = io_pipe_phv_in_data_151; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_152 = io_pipe_phv_in_data_152; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_153 = io_pipe_phv_in_data_153; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_154 = io_pipe_phv_in_data_154; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_155 = io_pipe_phv_in_data_155; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_156 = io_pipe_phv_in_data_156; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_157 = io_pipe_phv_in_data_157; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_158 = io_pipe_phv_in_data_158; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_159 = io_pipe_phv_in_data_159; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_160 = io_pipe_phv_in_data_160; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_161 = io_pipe_phv_in_data_161; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_162 = io_pipe_phv_in_data_162; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_163 = io_pipe_phv_in_data_163; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_164 = io_pipe_phv_in_data_164; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_165 = io_pipe_phv_in_data_165; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_166 = io_pipe_phv_in_data_166; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_167 = io_pipe_phv_in_data_167; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_168 = io_pipe_phv_in_data_168; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_169 = io_pipe_phv_in_data_169; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_170 = io_pipe_phv_in_data_170; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_171 = io_pipe_phv_in_data_171; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_172 = io_pipe_phv_in_data_172; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_173 = io_pipe_phv_in_data_173; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_174 = io_pipe_phv_in_data_174; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_175 = io_pipe_phv_in_data_175; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_176 = io_pipe_phv_in_data_176; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_177 = io_pipe_phv_in_data_177; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_178 = io_pipe_phv_in_data_178; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_179 = io_pipe_phv_in_data_179; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_180 = io_pipe_phv_in_data_180; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_181 = io_pipe_phv_in_data_181; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_182 = io_pipe_phv_in_data_182; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_183 = io_pipe_phv_in_data_183; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_184 = io_pipe_phv_in_data_184; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_185 = io_pipe_phv_in_data_185; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_186 = io_pipe_phv_in_data_186; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_187 = io_pipe_phv_in_data_187; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_188 = io_pipe_phv_in_data_188; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_189 = io_pipe_phv_in_data_189; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_190 = io_pipe_phv_in_data_190; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_191 = io_pipe_phv_in_data_191; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_192 = io_pipe_phv_in_data_192; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_193 = io_pipe_phv_in_data_193; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_194 = io_pipe_phv_in_data_194; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_195 = io_pipe_phv_in_data_195; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_196 = io_pipe_phv_in_data_196; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_197 = io_pipe_phv_in_data_197; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_198 = io_pipe_phv_in_data_198; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_199 = io_pipe_phv_in_data_199; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_200 = io_pipe_phv_in_data_200; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_201 = io_pipe_phv_in_data_201; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_202 = io_pipe_phv_in_data_202; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_203 = io_pipe_phv_in_data_203; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_204 = io_pipe_phv_in_data_204; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_205 = io_pipe_phv_in_data_205; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_206 = io_pipe_phv_in_data_206; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_207 = io_pipe_phv_in_data_207; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_208 = io_pipe_phv_in_data_208; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_209 = io_pipe_phv_in_data_209; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_210 = io_pipe_phv_in_data_210; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_211 = io_pipe_phv_in_data_211; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_212 = io_pipe_phv_in_data_212; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_213 = io_pipe_phv_in_data_213; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_214 = io_pipe_phv_in_data_214; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_215 = io_pipe_phv_in_data_215; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_216 = io_pipe_phv_in_data_216; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_217 = io_pipe_phv_in_data_217; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_218 = io_pipe_phv_in_data_218; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_219 = io_pipe_phv_in_data_219; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_220 = io_pipe_phv_in_data_220; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_221 = io_pipe_phv_in_data_221; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_222 = io_pipe_phv_in_data_222; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_223 = io_pipe_phv_in_data_223; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_224 = io_pipe_phv_in_data_224; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_225 = io_pipe_phv_in_data_225; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_226 = io_pipe_phv_in_data_226; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_227 = io_pipe_phv_in_data_227; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_228 = io_pipe_phv_in_data_228; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_229 = io_pipe_phv_in_data_229; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_230 = io_pipe_phv_in_data_230; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_231 = io_pipe_phv_in_data_231; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_232 = io_pipe_phv_in_data_232; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_233 = io_pipe_phv_in_data_233; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_234 = io_pipe_phv_in_data_234; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_235 = io_pipe_phv_in_data_235; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_236 = io_pipe_phv_in_data_236; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_237 = io_pipe_phv_in_data_237; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_238 = io_pipe_phv_in_data_238; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_239 = io_pipe_phv_in_data_239; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_240 = io_pipe_phv_in_data_240; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_241 = io_pipe_phv_in_data_241; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_242 = io_pipe_phv_in_data_242; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_243 = io_pipe_phv_in_data_243; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_244 = io_pipe_phv_in_data_244; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_245 = io_pipe_phv_in_data_245; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_246 = io_pipe_phv_in_data_246; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_247 = io_pipe_phv_in_data_247; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_248 = io_pipe_phv_in_data_248; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_249 = io_pipe_phv_in_data_249; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_250 = io_pipe_phv_in_data_250; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_251 = io_pipe_phv_in_data_251; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_252 = io_pipe_phv_in_data_252; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_253 = io_pipe_phv_in_data_253; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_254 = io_pipe_phv_in_data_254; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_255 = io_pipe_phv_in_data_255; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_256 = io_pipe_phv_in_data_256; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_257 = io_pipe_phv_in_data_257; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_258 = io_pipe_phv_in_data_258; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_259 = io_pipe_phv_in_data_259; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_260 = io_pipe_phv_in_data_260; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_261 = io_pipe_phv_in_data_261; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_262 = io_pipe_phv_in_data_262; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_263 = io_pipe_phv_in_data_263; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_264 = io_pipe_phv_in_data_264; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_265 = io_pipe_phv_in_data_265; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_266 = io_pipe_phv_in_data_266; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_267 = io_pipe_phv_in_data_267; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_268 = io_pipe_phv_in_data_268; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_269 = io_pipe_phv_in_data_269; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_270 = io_pipe_phv_in_data_270; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_271 = io_pipe_phv_in_data_271; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_272 = io_pipe_phv_in_data_272; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_273 = io_pipe_phv_in_data_273; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_274 = io_pipe_phv_in_data_274; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_275 = io_pipe_phv_in_data_275; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_276 = io_pipe_phv_in_data_276; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_277 = io_pipe_phv_in_data_277; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_278 = io_pipe_phv_in_data_278; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_279 = io_pipe_phv_in_data_279; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_280 = io_pipe_phv_in_data_280; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_281 = io_pipe_phv_in_data_281; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_282 = io_pipe_phv_in_data_282; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_283 = io_pipe_phv_in_data_283; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_284 = io_pipe_phv_in_data_284; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_285 = io_pipe_phv_in_data_285; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_286 = io_pipe_phv_in_data_286; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_287 = io_pipe_phv_in_data_287; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_288 = io_pipe_phv_in_data_288; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_289 = io_pipe_phv_in_data_289; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_290 = io_pipe_phv_in_data_290; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_291 = io_pipe_phv_in_data_291; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_292 = io_pipe_phv_in_data_292; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_293 = io_pipe_phv_in_data_293; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_294 = io_pipe_phv_in_data_294; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_295 = io_pipe_phv_in_data_295; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_296 = io_pipe_phv_in_data_296; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_297 = io_pipe_phv_in_data_297; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_298 = io_pipe_phv_in_data_298; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_299 = io_pipe_phv_in_data_299; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_300 = io_pipe_phv_in_data_300; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_301 = io_pipe_phv_in_data_301; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_302 = io_pipe_phv_in_data_302; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_303 = io_pipe_phv_in_data_303; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_304 = io_pipe_phv_in_data_304; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_305 = io_pipe_phv_in_data_305; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_306 = io_pipe_phv_in_data_306; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_307 = io_pipe_phv_in_data_307; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_308 = io_pipe_phv_in_data_308; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_309 = io_pipe_phv_in_data_309; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_310 = io_pipe_phv_in_data_310; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_311 = io_pipe_phv_in_data_311; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_312 = io_pipe_phv_in_data_312; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_313 = io_pipe_phv_in_data_313; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_314 = io_pipe_phv_in_data_314; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_315 = io_pipe_phv_in_data_315; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_316 = io_pipe_phv_in_data_316; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_317 = io_pipe_phv_in_data_317; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_318 = io_pipe_phv_in_data_318; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_319 = io_pipe_phv_in_data_319; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_320 = io_pipe_phv_in_data_320; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_321 = io_pipe_phv_in_data_321; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_322 = io_pipe_phv_in_data_322; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_323 = io_pipe_phv_in_data_323; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_324 = io_pipe_phv_in_data_324; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_325 = io_pipe_phv_in_data_325; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_326 = io_pipe_phv_in_data_326; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_327 = io_pipe_phv_in_data_327; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_328 = io_pipe_phv_in_data_328; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_329 = io_pipe_phv_in_data_329; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_330 = io_pipe_phv_in_data_330; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_331 = io_pipe_phv_in_data_331; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_332 = io_pipe_phv_in_data_332; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_333 = io_pipe_phv_in_data_333; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_334 = io_pipe_phv_in_data_334; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_335 = io_pipe_phv_in_data_335; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_336 = io_pipe_phv_in_data_336; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_337 = io_pipe_phv_in_data_337; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_338 = io_pipe_phv_in_data_338; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_339 = io_pipe_phv_in_data_339; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_340 = io_pipe_phv_in_data_340; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_341 = io_pipe_phv_in_data_341; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_342 = io_pipe_phv_in_data_342; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_343 = io_pipe_phv_in_data_343; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_344 = io_pipe_phv_in_data_344; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_345 = io_pipe_phv_in_data_345; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_346 = io_pipe_phv_in_data_346; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_347 = io_pipe_phv_in_data_347; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_348 = io_pipe_phv_in_data_348; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_349 = io_pipe_phv_in_data_349; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_350 = io_pipe_phv_in_data_350; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_351 = io_pipe_phv_in_data_351; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_352 = io_pipe_phv_in_data_352; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_353 = io_pipe_phv_in_data_353; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_354 = io_pipe_phv_in_data_354; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_355 = io_pipe_phv_in_data_355; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_356 = io_pipe_phv_in_data_356; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_357 = io_pipe_phv_in_data_357; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_358 = io_pipe_phv_in_data_358; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_359 = io_pipe_phv_in_data_359; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_360 = io_pipe_phv_in_data_360; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_361 = io_pipe_phv_in_data_361; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_362 = io_pipe_phv_in_data_362; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_363 = io_pipe_phv_in_data_363; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_364 = io_pipe_phv_in_data_364; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_365 = io_pipe_phv_in_data_365; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_366 = io_pipe_phv_in_data_366; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_367 = io_pipe_phv_in_data_367; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_368 = io_pipe_phv_in_data_368; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_369 = io_pipe_phv_in_data_369; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_370 = io_pipe_phv_in_data_370; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_371 = io_pipe_phv_in_data_371; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_372 = io_pipe_phv_in_data_372; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_373 = io_pipe_phv_in_data_373; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_374 = io_pipe_phv_in_data_374; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_375 = io_pipe_phv_in_data_375; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_376 = io_pipe_phv_in_data_376; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_377 = io_pipe_phv_in_data_377; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_378 = io_pipe_phv_in_data_378; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_379 = io_pipe_phv_in_data_379; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_380 = io_pipe_phv_in_data_380; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_381 = io_pipe_phv_in_data_381; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_382 = io_pipe_phv_in_data_382; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_383 = io_pipe_phv_in_data_383; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_384 = io_pipe_phv_in_data_384; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_385 = io_pipe_phv_in_data_385; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_386 = io_pipe_phv_in_data_386; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_387 = io_pipe_phv_in_data_387; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_388 = io_pipe_phv_in_data_388; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_389 = io_pipe_phv_in_data_389; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_390 = io_pipe_phv_in_data_390; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_391 = io_pipe_phv_in_data_391; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_392 = io_pipe_phv_in_data_392; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_393 = io_pipe_phv_in_data_393; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_394 = io_pipe_phv_in_data_394; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_395 = io_pipe_phv_in_data_395; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_396 = io_pipe_phv_in_data_396; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_397 = io_pipe_phv_in_data_397; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_398 = io_pipe_phv_in_data_398; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_399 = io_pipe_phv_in_data_399; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_400 = io_pipe_phv_in_data_400; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_401 = io_pipe_phv_in_data_401; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_402 = io_pipe_phv_in_data_402; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_403 = io_pipe_phv_in_data_403; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_404 = io_pipe_phv_in_data_404; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_405 = io_pipe_phv_in_data_405; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_406 = io_pipe_phv_in_data_406; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_407 = io_pipe_phv_in_data_407; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_408 = io_pipe_phv_in_data_408; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_409 = io_pipe_phv_in_data_409; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_410 = io_pipe_phv_in_data_410; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_411 = io_pipe_phv_in_data_411; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_412 = io_pipe_phv_in_data_412; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_413 = io_pipe_phv_in_data_413; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_414 = io_pipe_phv_in_data_414; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_415 = io_pipe_phv_in_data_415; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_416 = io_pipe_phv_in_data_416; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_417 = io_pipe_phv_in_data_417; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_418 = io_pipe_phv_in_data_418; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_419 = io_pipe_phv_in_data_419; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_420 = io_pipe_phv_in_data_420; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_421 = io_pipe_phv_in_data_421; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_422 = io_pipe_phv_in_data_422; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_423 = io_pipe_phv_in_data_423; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_424 = io_pipe_phv_in_data_424; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_425 = io_pipe_phv_in_data_425; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_426 = io_pipe_phv_in_data_426; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_427 = io_pipe_phv_in_data_427; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_428 = io_pipe_phv_in_data_428; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_429 = io_pipe_phv_in_data_429; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_430 = io_pipe_phv_in_data_430; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_431 = io_pipe_phv_in_data_431; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_432 = io_pipe_phv_in_data_432; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_433 = io_pipe_phv_in_data_433; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_434 = io_pipe_phv_in_data_434; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_435 = io_pipe_phv_in_data_435; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_436 = io_pipe_phv_in_data_436; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_437 = io_pipe_phv_in_data_437; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_438 = io_pipe_phv_in_data_438; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_439 = io_pipe_phv_in_data_439; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_440 = io_pipe_phv_in_data_440; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_441 = io_pipe_phv_in_data_441; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_442 = io_pipe_phv_in_data_442; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_443 = io_pipe_phv_in_data_443; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_444 = io_pipe_phv_in_data_444; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_445 = io_pipe_phv_in_data_445; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_446 = io_pipe_phv_in_data_446; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_447 = io_pipe_phv_in_data_447; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_448 = io_pipe_phv_in_data_448; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_449 = io_pipe_phv_in_data_449; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_450 = io_pipe_phv_in_data_450; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_451 = io_pipe_phv_in_data_451; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_452 = io_pipe_phv_in_data_452; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_453 = io_pipe_phv_in_data_453; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_454 = io_pipe_phv_in_data_454; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_455 = io_pipe_phv_in_data_455; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_456 = io_pipe_phv_in_data_456; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_457 = io_pipe_phv_in_data_457; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_458 = io_pipe_phv_in_data_458; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_459 = io_pipe_phv_in_data_459; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_460 = io_pipe_phv_in_data_460; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_461 = io_pipe_phv_in_data_461; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_462 = io_pipe_phv_in_data_462; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_463 = io_pipe_phv_in_data_463; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_464 = io_pipe_phv_in_data_464; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_465 = io_pipe_phv_in_data_465; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_466 = io_pipe_phv_in_data_466; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_467 = io_pipe_phv_in_data_467; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_468 = io_pipe_phv_in_data_468; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_469 = io_pipe_phv_in_data_469; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_470 = io_pipe_phv_in_data_470; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_471 = io_pipe_phv_in_data_471; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_472 = io_pipe_phv_in_data_472; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_473 = io_pipe_phv_in_data_473; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_474 = io_pipe_phv_in_data_474; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_475 = io_pipe_phv_in_data_475; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_476 = io_pipe_phv_in_data_476; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_477 = io_pipe_phv_in_data_477; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_478 = io_pipe_phv_in_data_478; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_479 = io_pipe_phv_in_data_479; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_480 = io_pipe_phv_in_data_480; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_481 = io_pipe_phv_in_data_481; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_482 = io_pipe_phv_in_data_482; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_483 = io_pipe_phv_in_data_483; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_484 = io_pipe_phv_in_data_484; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_485 = io_pipe_phv_in_data_485; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_486 = io_pipe_phv_in_data_486; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_487 = io_pipe_phv_in_data_487; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_488 = io_pipe_phv_in_data_488; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_489 = io_pipe_phv_in_data_489; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_490 = io_pipe_phv_in_data_490; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_491 = io_pipe_phv_in_data_491; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_492 = io_pipe_phv_in_data_492; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_493 = io_pipe_phv_in_data_493; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_494 = io_pipe_phv_in_data_494; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_495 = io_pipe_phv_in_data_495; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_496 = io_pipe_phv_in_data_496; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_497 = io_pipe_phv_in_data_497; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_498 = io_pipe_phv_in_data_498; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_499 = io_pipe_phv_in_data_499; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_500 = io_pipe_phv_in_data_500; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_501 = io_pipe_phv_in_data_501; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_502 = io_pipe_phv_in_data_502; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_503 = io_pipe_phv_in_data_503; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_504 = io_pipe_phv_in_data_504; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_505 = io_pipe_phv_in_data_505; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_506 = io_pipe_phv_in_data_506; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_507 = io_pipe_phv_in_data_507; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_508 = io_pipe_phv_in_data_508; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_509 = io_pipe_phv_in_data_509; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_510 = io_pipe_phv_in_data_510; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_data_511 = io_pipe_phv_in_data_511; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_0 = io_pipe_phv_in_header_0; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_1 = io_pipe_phv_in_header_1; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_2 = io_pipe_phv_in_header_2; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_3 = io_pipe_phv_in_header_3; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_4 = io_pipe_phv_in_header_4; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_5 = io_pipe_phv_in_header_5; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_6 = io_pipe_phv_in_header_6; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_7 = io_pipe_phv_in_header_7; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_8 = io_pipe_phv_in_header_8; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_9 = io_pipe_phv_in_header_9; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_10 = io_pipe_phv_in_header_10; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_11 = io_pipe_phv_in_header_11; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_12 = io_pipe_phv_in_header_12; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_13 = io_pipe_phv_in_header_13; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_14 = io_pipe_phv_in_header_14; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_header_15 = io_pipe_phv_in_header_15; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_parse_current_state = io_pipe_phv_in_parse_current_state; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_parse_current_offset = io_pipe_phv_in_parse_current_offset; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_parse_transition_field = io_pipe_phv_in_parse_transition_field; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_next_processor_id = io_pipe_phv_in_next_processor_id; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_next_config_id = io_pipe_phv_in_next_config_id; // @[executor.scala 496:26]
  assign pipe1_io_pipe_phv_in_is_valid_processor = io_pipe_phv_in_is_valid_processor; // @[executor.scala 496:26]
  assign pipe1_io_hit = io_hit; // @[executor.scala 497:26]
  assign pipe1_io_match_value = io_match_value; // @[executor.scala 498:26]
  assign pipe1_io_action_mod_en_0 = io_action_mod_en_0; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_en_1 = io_action_mod_en_1; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_addr = io_action_mod_addr; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_data_0 = io_action_mod_data_0; // @[executor.scala 499:26]
  assign pipe1_io_action_mod_data_1 = io_action_mod_data_1; // @[executor.scala 499:26]
  assign pipe2_clock = clock;
  assign pipe2_io_pipe_phv_in_data_0 = pipe1_io_pipe_phv_out_data_0; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_1 = pipe1_io_pipe_phv_out_data_1; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_2 = pipe1_io_pipe_phv_out_data_2; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_3 = pipe1_io_pipe_phv_out_data_3; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_4 = pipe1_io_pipe_phv_out_data_4; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_5 = pipe1_io_pipe_phv_out_data_5; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_6 = pipe1_io_pipe_phv_out_data_6; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_7 = pipe1_io_pipe_phv_out_data_7; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_8 = pipe1_io_pipe_phv_out_data_8; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_9 = pipe1_io_pipe_phv_out_data_9; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_10 = pipe1_io_pipe_phv_out_data_10; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_11 = pipe1_io_pipe_phv_out_data_11; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_12 = pipe1_io_pipe_phv_out_data_12; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_13 = pipe1_io_pipe_phv_out_data_13; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_14 = pipe1_io_pipe_phv_out_data_14; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_15 = pipe1_io_pipe_phv_out_data_15; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_16 = pipe1_io_pipe_phv_out_data_16; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_17 = pipe1_io_pipe_phv_out_data_17; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_18 = pipe1_io_pipe_phv_out_data_18; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_19 = pipe1_io_pipe_phv_out_data_19; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_20 = pipe1_io_pipe_phv_out_data_20; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_21 = pipe1_io_pipe_phv_out_data_21; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_22 = pipe1_io_pipe_phv_out_data_22; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_23 = pipe1_io_pipe_phv_out_data_23; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_24 = pipe1_io_pipe_phv_out_data_24; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_25 = pipe1_io_pipe_phv_out_data_25; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_26 = pipe1_io_pipe_phv_out_data_26; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_27 = pipe1_io_pipe_phv_out_data_27; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_28 = pipe1_io_pipe_phv_out_data_28; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_29 = pipe1_io_pipe_phv_out_data_29; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_30 = pipe1_io_pipe_phv_out_data_30; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_31 = pipe1_io_pipe_phv_out_data_31; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_32 = pipe1_io_pipe_phv_out_data_32; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_33 = pipe1_io_pipe_phv_out_data_33; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_34 = pipe1_io_pipe_phv_out_data_34; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_35 = pipe1_io_pipe_phv_out_data_35; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_36 = pipe1_io_pipe_phv_out_data_36; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_37 = pipe1_io_pipe_phv_out_data_37; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_38 = pipe1_io_pipe_phv_out_data_38; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_39 = pipe1_io_pipe_phv_out_data_39; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_40 = pipe1_io_pipe_phv_out_data_40; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_41 = pipe1_io_pipe_phv_out_data_41; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_42 = pipe1_io_pipe_phv_out_data_42; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_43 = pipe1_io_pipe_phv_out_data_43; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_44 = pipe1_io_pipe_phv_out_data_44; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_45 = pipe1_io_pipe_phv_out_data_45; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_46 = pipe1_io_pipe_phv_out_data_46; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_47 = pipe1_io_pipe_phv_out_data_47; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_48 = pipe1_io_pipe_phv_out_data_48; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_49 = pipe1_io_pipe_phv_out_data_49; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_50 = pipe1_io_pipe_phv_out_data_50; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_51 = pipe1_io_pipe_phv_out_data_51; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_52 = pipe1_io_pipe_phv_out_data_52; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_53 = pipe1_io_pipe_phv_out_data_53; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_54 = pipe1_io_pipe_phv_out_data_54; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_55 = pipe1_io_pipe_phv_out_data_55; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_56 = pipe1_io_pipe_phv_out_data_56; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_57 = pipe1_io_pipe_phv_out_data_57; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_58 = pipe1_io_pipe_phv_out_data_58; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_59 = pipe1_io_pipe_phv_out_data_59; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_60 = pipe1_io_pipe_phv_out_data_60; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_61 = pipe1_io_pipe_phv_out_data_61; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_62 = pipe1_io_pipe_phv_out_data_62; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_63 = pipe1_io_pipe_phv_out_data_63; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_64 = pipe1_io_pipe_phv_out_data_64; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_65 = pipe1_io_pipe_phv_out_data_65; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_66 = pipe1_io_pipe_phv_out_data_66; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_67 = pipe1_io_pipe_phv_out_data_67; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_68 = pipe1_io_pipe_phv_out_data_68; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_69 = pipe1_io_pipe_phv_out_data_69; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_70 = pipe1_io_pipe_phv_out_data_70; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_71 = pipe1_io_pipe_phv_out_data_71; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_72 = pipe1_io_pipe_phv_out_data_72; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_73 = pipe1_io_pipe_phv_out_data_73; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_74 = pipe1_io_pipe_phv_out_data_74; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_75 = pipe1_io_pipe_phv_out_data_75; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_76 = pipe1_io_pipe_phv_out_data_76; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_77 = pipe1_io_pipe_phv_out_data_77; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_78 = pipe1_io_pipe_phv_out_data_78; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_79 = pipe1_io_pipe_phv_out_data_79; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_80 = pipe1_io_pipe_phv_out_data_80; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_81 = pipe1_io_pipe_phv_out_data_81; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_82 = pipe1_io_pipe_phv_out_data_82; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_83 = pipe1_io_pipe_phv_out_data_83; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_84 = pipe1_io_pipe_phv_out_data_84; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_85 = pipe1_io_pipe_phv_out_data_85; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_86 = pipe1_io_pipe_phv_out_data_86; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_87 = pipe1_io_pipe_phv_out_data_87; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_88 = pipe1_io_pipe_phv_out_data_88; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_89 = pipe1_io_pipe_phv_out_data_89; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_90 = pipe1_io_pipe_phv_out_data_90; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_91 = pipe1_io_pipe_phv_out_data_91; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_92 = pipe1_io_pipe_phv_out_data_92; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_93 = pipe1_io_pipe_phv_out_data_93; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_94 = pipe1_io_pipe_phv_out_data_94; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_95 = pipe1_io_pipe_phv_out_data_95; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_96 = pipe1_io_pipe_phv_out_data_96; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_97 = pipe1_io_pipe_phv_out_data_97; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_98 = pipe1_io_pipe_phv_out_data_98; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_99 = pipe1_io_pipe_phv_out_data_99; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_100 = pipe1_io_pipe_phv_out_data_100; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_101 = pipe1_io_pipe_phv_out_data_101; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_102 = pipe1_io_pipe_phv_out_data_102; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_103 = pipe1_io_pipe_phv_out_data_103; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_104 = pipe1_io_pipe_phv_out_data_104; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_105 = pipe1_io_pipe_phv_out_data_105; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_106 = pipe1_io_pipe_phv_out_data_106; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_107 = pipe1_io_pipe_phv_out_data_107; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_108 = pipe1_io_pipe_phv_out_data_108; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_109 = pipe1_io_pipe_phv_out_data_109; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_110 = pipe1_io_pipe_phv_out_data_110; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_111 = pipe1_io_pipe_phv_out_data_111; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_112 = pipe1_io_pipe_phv_out_data_112; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_113 = pipe1_io_pipe_phv_out_data_113; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_114 = pipe1_io_pipe_phv_out_data_114; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_115 = pipe1_io_pipe_phv_out_data_115; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_116 = pipe1_io_pipe_phv_out_data_116; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_117 = pipe1_io_pipe_phv_out_data_117; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_118 = pipe1_io_pipe_phv_out_data_118; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_119 = pipe1_io_pipe_phv_out_data_119; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_120 = pipe1_io_pipe_phv_out_data_120; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_121 = pipe1_io_pipe_phv_out_data_121; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_122 = pipe1_io_pipe_phv_out_data_122; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_123 = pipe1_io_pipe_phv_out_data_123; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_124 = pipe1_io_pipe_phv_out_data_124; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_125 = pipe1_io_pipe_phv_out_data_125; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_126 = pipe1_io_pipe_phv_out_data_126; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_127 = pipe1_io_pipe_phv_out_data_127; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_128 = pipe1_io_pipe_phv_out_data_128; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_129 = pipe1_io_pipe_phv_out_data_129; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_130 = pipe1_io_pipe_phv_out_data_130; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_131 = pipe1_io_pipe_phv_out_data_131; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_132 = pipe1_io_pipe_phv_out_data_132; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_133 = pipe1_io_pipe_phv_out_data_133; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_134 = pipe1_io_pipe_phv_out_data_134; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_135 = pipe1_io_pipe_phv_out_data_135; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_136 = pipe1_io_pipe_phv_out_data_136; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_137 = pipe1_io_pipe_phv_out_data_137; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_138 = pipe1_io_pipe_phv_out_data_138; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_139 = pipe1_io_pipe_phv_out_data_139; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_140 = pipe1_io_pipe_phv_out_data_140; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_141 = pipe1_io_pipe_phv_out_data_141; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_142 = pipe1_io_pipe_phv_out_data_142; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_143 = pipe1_io_pipe_phv_out_data_143; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_144 = pipe1_io_pipe_phv_out_data_144; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_145 = pipe1_io_pipe_phv_out_data_145; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_146 = pipe1_io_pipe_phv_out_data_146; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_147 = pipe1_io_pipe_phv_out_data_147; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_148 = pipe1_io_pipe_phv_out_data_148; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_149 = pipe1_io_pipe_phv_out_data_149; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_150 = pipe1_io_pipe_phv_out_data_150; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_151 = pipe1_io_pipe_phv_out_data_151; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_152 = pipe1_io_pipe_phv_out_data_152; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_153 = pipe1_io_pipe_phv_out_data_153; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_154 = pipe1_io_pipe_phv_out_data_154; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_155 = pipe1_io_pipe_phv_out_data_155; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_156 = pipe1_io_pipe_phv_out_data_156; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_157 = pipe1_io_pipe_phv_out_data_157; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_158 = pipe1_io_pipe_phv_out_data_158; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_159 = pipe1_io_pipe_phv_out_data_159; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_160 = pipe1_io_pipe_phv_out_data_160; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_161 = pipe1_io_pipe_phv_out_data_161; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_162 = pipe1_io_pipe_phv_out_data_162; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_163 = pipe1_io_pipe_phv_out_data_163; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_164 = pipe1_io_pipe_phv_out_data_164; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_165 = pipe1_io_pipe_phv_out_data_165; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_166 = pipe1_io_pipe_phv_out_data_166; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_167 = pipe1_io_pipe_phv_out_data_167; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_168 = pipe1_io_pipe_phv_out_data_168; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_169 = pipe1_io_pipe_phv_out_data_169; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_170 = pipe1_io_pipe_phv_out_data_170; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_171 = pipe1_io_pipe_phv_out_data_171; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_172 = pipe1_io_pipe_phv_out_data_172; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_173 = pipe1_io_pipe_phv_out_data_173; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_174 = pipe1_io_pipe_phv_out_data_174; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_175 = pipe1_io_pipe_phv_out_data_175; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_176 = pipe1_io_pipe_phv_out_data_176; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_177 = pipe1_io_pipe_phv_out_data_177; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_178 = pipe1_io_pipe_phv_out_data_178; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_179 = pipe1_io_pipe_phv_out_data_179; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_180 = pipe1_io_pipe_phv_out_data_180; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_181 = pipe1_io_pipe_phv_out_data_181; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_182 = pipe1_io_pipe_phv_out_data_182; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_183 = pipe1_io_pipe_phv_out_data_183; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_184 = pipe1_io_pipe_phv_out_data_184; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_185 = pipe1_io_pipe_phv_out_data_185; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_186 = pipe1_io_pipe_phv_out_data_186; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_187 = pipe1_io_pipe_phv_out_data_187; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_188 = pipe1_io_pipe_phv_out_data_188; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_189 = pipe1_io_pipe_phv_out_data_189; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_190 = pipe1_io_pipe_phv_out_data_190; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_191 = pipe1_io_pipe_phv_out_data_191; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_192 = pipe1_io_pipe_phv_out_data_192; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_193 = pipe1_io_pipe_phv_out_data_193; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_194 = pipe1_io_pipe_phv_out_data_194; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_195 = pipe1_io_pipe_phv_out_data_195; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_196 = pipe1_io_pipe_phv_out_data_196; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_197 = pipe1_io_pipe_phv_out_data_197; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_198 = pipe1_io_pipe_phv_out_data_198; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_199 = pipe1_io_pipe_phv_out_data_199; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_200 = pipe1_io_pipe_phv_out_data_200; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_201 = pipe1_io_pipe_phv_out_data_201; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_202 = pipe1_io_pipe_phv_out_data_202; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_203 = pipe1_io_pipe_phv_out_data_203; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_204 = pipe1_io_pipe_phv_out_data_204; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_205 = pipe1_io_pipe_phv_out_data_205; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_206 = pipe1_io_pipe_phv_out_data_206; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_207 = pipe1_io_pipe_phv_out_data_207; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_208 = pipe1_io_pipe_phv_out_data_208; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_209 = pipe1_io_pipe_phv_out_data_209; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_210 = pipe1_io_pipe_phv_out_data_210; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_211 = pipe1_io_pipe_phv_out_data_211; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_212 = pipe1_io_pipe_phv_out_data_212; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_213 = pipe1_io_pipe_phv_out_data_213; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_214 = pipe1_io_pipe_phv_out_data_214; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_215 = pipe1_io_pipe_phv_out_data_215; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_216 = pipe1_io_pipe_phv_out_data_216; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_217 = pipe1_io_pipe_phv_out_data_217; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_218 = pipe1_io_pipe_phv_out_data_218; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_219 = pipe1_io_pipe_phv_out_data_219; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_220 = pipe1_io_pipe_phv_out_data_220; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_221 = pipe1_io_pipe_phv_out_data_221; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_222 = pipe1_io_pipe_phv_out_data_222; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_223 = pipe1_io_pipe_phv_out_data_223; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_224 = pipe1_io_pipe_phv_out_data_224; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_225 = pipe1_io_pipe_phv_out_data_225; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_226 = pipe1_io_pipe_phv_out_data_226; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_227 = pipe1_io_pipe_phv_out_data_227; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_228 = pipe1_io_pipe_phv_out_data_228; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_229 = pipe1_io_pipe_phv_out_data_229; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_230 = pipe1_io_pipe_phv_out_data_230; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_231 = pipe1_io_pipe_phv_out_data_231; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_232 = pipe1_io_pipe_phv_out_data_232; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_233 = pipe1_io_pipe_phv_out_data_233; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_234 = pipe1_io_pipe_phv_out_data_234; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_235 = pipe1_io_pipe_phv_out_data_235; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_236 = pipe1_io_pipe_phv_out_data_236; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_237 = pipe1_io_pipe_phv_out_data_237; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_238 = pipe1_io_pipe_phv_out_data_238; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_239 = pipe1_io_pipe_phv_out_data_239; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_240 = pipe1_io_pipe_phv_out_data_240; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_241 = pipe1_io_pipe_phv_out_data_241; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_242 = pipe1_io_pipe_phv_out_data_242; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_243 = pipe1_io_pipe_phv_out_data_243; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_244 = pipe1_io_pipe_phv_out_data_244; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_245 = pipe1_io_pipe_phv_out_data_245; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_246 = pipe1_io_pipe_phv_out_data_246; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_247 = pipe1_io_pipe_phv_out_data_247; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_248 = pipe1_io_pipe_phv_out_data_248; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_249 = pipe1_io_pipe_phv_out_data_249; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_250 = pipe1_io_pipe_phv_out_data_250; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_251 = pipe1_io_pipe_phv_out_data_251; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_252 = pipe1_io_pipe_phv_out_data_252; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_253 = pipe1_io_pipe_phv_out_data_253; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_254 = pipe1_io_pipe_phv_out_data_254; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_255 = pipe1_io_pipe_phv_out_data_255; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_256 = pipe1_io_pipe_phv_out_data_256; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_257 = pipe1_io_pipe_phv_out_data_257; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_258 = pipe1_io_pipe_phv_out_data_258; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_259 = pipe1_io_pipe_phv_out_data_259; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_260 = pipe1_io_pipe_phv_out_data_260; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_261 = pipe1_io_pipe_phv_out_data_261; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_262 = pipe1_io_pipe_phv_out_data_262; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_263 = pipe1_io_pipe_phv_out_data_263; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_264 = pipe1_io_pipe_phv_out_data_264; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_265 = pipe1_io_pipe_phv_out_data_265; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_266 = pipe1_io_pipe_phv_out_data_266; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_267 = pipe1_io_pipe_phv_out_data_267; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_268 = pipe1_io_pipe_phv_out_data_268; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_269 = pipe1_io_pipe_phv_out_data_269; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_270 = pipe1_io_pipe_phv_out_data_270; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_271 = pipe1_io_pipe_phv_out_data_271; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_272 = pipe1_io_pipe_phv_out_data_272; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_273 = pipe1_io_pipe_phv_out_data_273; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_274 = pipe1_io_pipe_phv_out_data_274; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_275 = pipe1_io_pipe_phv_out_data_275; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_276 = pipe1_io_pipe_phv_out_data_276; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_277 = pipe1_io_pipe_phv_out_data_277; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_278 = pipe1_io_pipe_phv_out_data_278; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_279 = pipe1_io_pipe_phv_out_data_279; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_280 = pipe1_io_pipe_phv_out_data_280; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_281 = pipe1_io_pipe_phv_out_data_281; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_282 = pipe1_io_pipe_phv_out_data_282; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_283 = pipe1_io_pipe_phv_out_data_283; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_284 = pipe1_io_pipe_phv_out_data_284; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_285 = pipe1_io_pipe_phv_out_data_285; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_286 = pipe1_io_pipe_phv_out_data_286; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_287 = pipe1_io_pipe_phv_out_data_287; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_288 = pipe1_io_pipe_phv_out_data_288; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_289 = pipe1_io_pipe_phv_out_data_289; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_290 = pipe1_io_pipe_phv_out_data_290; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_291 = pipe1_io_pipe_phv_out_data_291; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_292 = pipe1_io_pipe_phv_out_data_292; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_293 = pipe1_io_pipe_phv_out_data_293; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_294 = pipe1_io_pipe_phv_out_data_294; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_295 = pipe1_io_pipe_phv_out_data_295; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_296 = pipe1_io_pipe_phv_out_data_296; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_297 = pipe1_io_pipe_phv_out_data_297; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_298 = pipe1_io_pipe_phv_out_data_298; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_299 = pipe1_io_pipe_phv_out_data_299; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_300 = pipe1_io_pipe_phv_out_data_300; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_301 = pipe1_io_pipe_phv_out_data_301; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_302 = pipe1_io_pipe_phv_out_data_302; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_303 = pipe1_io_pipe_phv_out_data_303; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_304 = pipe1_io_pipe_phv_out_data_304; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_305 = pipe1_io_pipe_phv_out_data_305; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_306 = pipe1_io_pipe_phv_out_data_306; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_307 = pipe1_io_pipe_phv_out_data_307; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_308 = pipe1_io_pipe_phv_out_data_308; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_309 = pipe1_io_pipe_phv_out_data_309; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_310 = pipe1_io_pipe_phv_out_data_310; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_311 = pipe1_io_pipe_phv_out_data_311; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_312 = pipe1_io_pipe_phv_out_data_312; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_313 = pipe1_io_pipe_phv_out_data_313; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_314 = pipe1_io_pipe_phv_out_data_314; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_315 = pipe1_io_pipe_phv_out_data_315; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_316 = pipe1_io_pipe_phv_out_data_316; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_317 = pipe1_io_pipe_phv_out_data_317; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_318 = pipe1_io_pipe_phv_out_data_318; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_319 = pipe1_io_pipe_phv_out_data_319; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_320 = pipe1_io_pipe_phv_out_data_320; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_321 = pipe1_io_pipe_phv_out_data_321; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_322 = pipe1_io_pipe_phv_out_data_322; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_323 = pipe1_io_pipe_phv_out_data_323; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_324 = pipe1_io_pipe_phv_out_data_324; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_325 = pipe1_io_pipe_phv_out_data_325; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_326 = pipe1_io_pipe_phv_out_data_326; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_327 = pipe1_io_pipe_phv_out_data_327; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_328 = pipe1_io_pipe_phv_out_data_328; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_329 = pipe1_io_pipe_phv_out_data_329; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_330 = pipe1_io_pipe_phv_out_data_330; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_331 = pipe1_io_pipe_phv_out_data_331; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_332 = pipe1_io_pipe_phv_out_data_332; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_333 = pipe1_io_pipe_phv_out_data_333; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_334 = pipe1_io_pipe_phv_out_data_334; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_335 = pipe1_io_pipe_phv_out_data_335; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_336 = pipe1_io_pipe_phv_out_data_336; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_337 = pipe1_io_pipe_phv_out_data_337; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_338 = pipe1_io_pipe_phv_out_data_338; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_339 = pipe1_io_pipe_phv_out_data_339; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_340 = pipe1_io_pipe_phv_out_data_340; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_341 = pipe1_io_pipe_phv_out_data_341; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_342 = pipe1_io_pipe_phv_out_data_342; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_343 = pipe1_io_pipe_phv_out_data_343; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_344 = pipe1_io_pipe_phv_out_data_344; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_345 = pipe1_io_pipe_phv_out_data_345; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_346 = pipe1_io_pipe_phv_out_data_346; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_347 = pipe1_io_pipe_phv_out_data_347; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_348 = pipe1_io_pipe_phv_out_data_348; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_349 = pipe1_io_pipe_phv_out_data_349; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_350 = pipe1_io_pipe_phv_out_data_350; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_351 = pipe1_io_pipe_phv_out_data_351; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_352 = pipe1_io_pipe_phv_out_data_352; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_353 = pipe1_io_pipe_phv_out_data_353; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_354 = pipe1_io_pipe_phv_out_data_354; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_355 = pipe1_io_pipe_phv_out_data_355; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_356 = pipe1_io_pipe_phv_out_data_356; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_357 = pipe1_io_pipe_phv_out_data_357; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_358 = pipe1_io_pipe_phv_out_data_358; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_359 = pipe1_io_pipe_phv_out_data_359; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_360 = pipe1_io_pipe_phv_out_data_360; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_361 = pipe1_io_pipe_phv_out_data_361; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_362 = pipe1_io_pipe_phv_out_data_362; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_363 = pipe1_io_pipe_phv_out_data_363; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_364 = pipe1_io_pipe_phv_out_data_364; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_365 = pipe1_io_pipe_phv_out_data_365; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_366 = pipe1_io_pipe_phv_out_data_366; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_367 = pipe1_io_pipe_phv_out_data_367; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_368 = pipe1_io_pipe_phv_out_data_368; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_369 = pipe1_io_pipe_phv_out_data_369; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_370 = pipe1_io_pipe_phv_out_data_370; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_371 = pipe1_io_pipe_phv_out_data_371; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_372 = pipe1_io_pipe_phv_out_data_372; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_373 = pipe1_io_pipe_phv_out_data_373; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_374 = pipe1_io_pipe_phv_out_data_374; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_375 = pipe1_io_pipe_phv_out_data_375; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_376 = pipe1_io_pipe_phv_out_data_376; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_377 = pipe1_io_pipe_phv_out_data_377; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_378 = pipe1_io_pipe_phv_out_data_378; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_379 = pipe1_io_pipe_phv_out_data_379; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_380 = pipe1_io_pipe_phv_out_data_380; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_381 = pipe1_io_pipe_phv_out_data_381; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_382 = pipe1_io_pipe_phv_out_data_382; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_383 = pipe1_io_pipe_phv_out_data_383; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_384 = pipe1_io_pipe_phv_out_data_384; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_385 = pipe1_io_pipe_phv_out_data_385; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_386 = pipe1_io_pipe_phv_out_data_386; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_387 = pipe1_io_pipe_phv_out_data_387; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_388 = pipe1_io_pipe_phv_out_data_388; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_389 = pipe1_io_pipe_phv_out_data_389; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_390 = pipe1_io_pipe_phv_out_data_390; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_391 = pipe1_io_pipe_phv_out_data_391; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_392 = pipe1_io_pipe_phv_out_data_392; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_393 = pipe1_io_pipe_phv_out_data_393; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_394 = pipe1_io_pipe_phv_out_data_394; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_395 = pipe1_io_pipe_phv_out_data_395; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_396 = pipe1_io_pipe_phv_out_data_396; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_397 = pipe1_io_pipe_phv_out_data_397; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_398 = pipe1_io_pipe_phv_out_data_398; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_399 = pipe1_io_pipe_phv_out_data_399; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_400 = pipe1_io_pipe_phv_out_data_400; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_401 = pipe1_io_pipe_phv_out_data_401; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_402 = pipe1_io_pipe_phv_out_data_402; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_403 = pipe1_io_pipe_phv_out_data_403; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_404 = pipe1_io_pipe_phv_out_data_404; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_405 = pipe1_io_pipe_phv_out_data_405; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_406 = pipe1_io_pipe_phv_out_data_406; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_407 = pipe1_io_pipe_phv_out_data_407; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_408 = pipe1_io_pipe_phv_out_data_408; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_409 = pipe1_io_pipe_phv_out_data_409; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_410 = pipe1_io_pipe_phv_out_data_410; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_411 = pipe1_io_pipe_phv_out_data_411; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_412 = pipe1_io_pipe_phv_out_data_412; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_413 = pipe1_io_pipe_phv_out_data_413; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_414 = pipe1_io_pipe_phv_out_data_414; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_415 = pipe1_io_pipe_phv_out_data_415; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_416 = pipe1_io_pipe_phv_out_data_416; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_417 = pipe1_io_pipe_phv_out_data_417; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_418 = pipe1_io_pipe_phv_out_data_418; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_419 = pipe1_io_pipe_phv_out_data_419; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_420 = pipe1_io_pipe_phv_out_data_420; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_421 = pipe1_io_pipe_phv_out_data_421; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_422 = pipe1_io_pipe_phv_out_data_422; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_423 = pipe1_io_pipe_phv_out_data_423; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_424 = pipe1_io_pipe_phv_out_data_424; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_425 = pipe1_io_pipe_phv_out_data_425; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_426 = pipe1_io_pipe_phv_out_data_426; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_427 = pipe1_io_pipe_phv_out_data_427; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_428 = pipe1_io_pipe_phv_out_data_428; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_429 = pipe1_io_pipe_phv_out_data_429; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_430 = pipe1_io_pipe_phv_out_data_430; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_431 = pipe1_io_pipe_phv_out_data_431; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_432 = pipe1_io_pipe_phv_out_data_432; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_433 = pipe1_io_pipe_phv_out_data_433; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_434 = pipe1_io_pipe_phv_out_data_434; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_435 = pipe1_io_pipe_phv_out_data_435; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_436 = pipe1_io_pipe_phv_out_data_436; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_437 = pipe1_io_pipe_phv_out_data_437; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_438 = pipe1_io_pipe_phv_out_data_438; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_439 = pipe1_io_pipe_phv_out_data_439; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_440 = pipe1_io_pipe_phv_out_data_440; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_441 = pipe1_io_pipe_phv_out_data_441; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_442 = pipe1_io_pipe_phv_out_data_442; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_443 = pipe1_io_pipe_phv_out_data_443; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_444 = pipe1_io_pipe_phv_out_data_444; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_445 = pipe1_io_pipe_phv_out_data_445; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_446 = pipe1_io_pipe_phv_out_data_446; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_447 = pipe1_io_pipe_phv_out_data_447; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_448 = pipe1_io_pipe_phv_out_data_448; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_449 = pipe1_io_pipe_phv_out_data_449; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_450 = pipe1_io_pipe_phv_out_data_450; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_451 = pipe1_io_pipe_phv_out_data_451; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_452 = pipe1_io_pipe_phv_out_data_452; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_453 = pipe1_io_pipe_phv_out_data_453; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_454 = pipe1_io_pipe_phv_out_data_454; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_455 = pipe1_io_pipe_phv_out_data_455; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_456 = pipe1_io_pipe_phv_out_data_456; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_457 = pipe1_io_pipe_phv_out_data_457; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_458 = pipe1_io_pipe_phv_out_data_458; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_459 = pipe1_io_pipe_phv_out_data_459; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_460 = pipe1_io_pipe_phv_out_data_460; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_461 = pipe1_io_pipe_phv_out_data_461; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_462 = pipe1_io_pipe_phv_out_data_462; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_463 = pipe1_io_pipe_phv_out_data_463; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_464 = pipe1_io_pipe_phv_out_data_464; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_465 = pipe1_io_pipe_phv_out_data_465; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_466 = pipe1_io_pipe_phv_out_data_466; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_467 = pipe1_io_pipe_phv_out_data_467; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_468 = pipe1_io_pipe_phv_out_data_468; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_469 = pipe1_io_pipe_phv_out_data_469; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_470 = pipe1_io_pipe_phv_out_data_470; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_471 = pipe1_io_pipe_phv_out_data_471; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_472 = pipe1_io_pipe_phv_out_data_472; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_473 = pipe1_io_pipe_phv_out_data_473; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_474 = pipe1_io_pipe_phv_out_data_474; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_475 = pipe1_io_pipe_phv_out_data_475; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_476 = pipe1_io_pipe_phv_out_data_476; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_477 = pipe1_io_pipe_phv_out_data_477; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_478 = pipe1_io_pipe_phv_out_data_478; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_479 = pipe1_io_pipe_phv_out_data_479; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_480 = pipe1_io_pipe_phv_out_data_480; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_481 = pipe1_io_pipe_phv_out_data_481; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_482 = pipe1_io_pipe_phv_out_data_482; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_483 = pipe1_io_pipe_phv_out_data_483; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_484 = pipe1_io_pipe_phv_out_data_484; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_485 = pipe1_io_pipe_phv_out_data_485; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_486 = pipe1_io_pipe_phv_out_data_486; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_487 = pipe1_io_pipe_phv_out_data_487; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_488 = pipe1_io_pipe_phv_out_data_488; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_489 = pipe1_io_pipe_phv_out_data_489; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_490 = pipe1_io_pipe_phv_out_data_490; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_491 = pipe1_io_pipe_phv_out_data_491; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_492 = pipe1_io_pipe_phv_out_data_492; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_493 = pipe1_io_pipe_phv_out_data_493; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_494 = pipe1_io_pipe_phv_out_data_494; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_495 = pipe1_io_pipe_phv_out_data_495; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_496 = pipe1_io_pipe_phv_out_data_496; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_497 = pipe1_io_pipe_phv_out_data_497; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_498 = pipe1_io_pipe_phv_out_data_498; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_499 = pipe1_io_pipe_phv_out_data_499; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_500 = pipe1_io_pipe_phv_out_data_500; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_501 = pipe1_io_pipe_phv_out_data_501; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_502 = pipe1_io_pipe_phv_out_data_502; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_503 = pipe1_io_pipe_phv_out_data_503; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_504 = pipe1_io_pipe_phv_out_data_504; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_505 = pipe1_io_pipe_phv_out_data_505; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_506 = pipe1_io_pipe_phv_out_data_506; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_507 = pipe1_io_pipe_phv_out_data_507; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_508 = pipe1_io_pipe_phv_out_data_508; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_509 = pipe1_io_pipe_phv_out_data_509; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_510 = pipe1_io_pipe_phv_out_data_510; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_data_511 = pipe1_io_pipe_phv_out_data_511; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_0 = pipe1_io_pipe_phv_out_header_0; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_1 = pipe1_io_pipe_phv_out_header_1; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_2 = pipe1_io_pipe_phv_out_header_2; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_3 = pipe1_io_pipe_phv_out_header_3; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_4 = pipe1_io_pipe_phv_out_header_4; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_5 = pipe1_io_pipe_phv_out_header_5; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_6 = pipe1_io_pipe_phv_out_header_6; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_7 = pipe1_io_pipe_phv_out_header_7; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_8 = pipe1_io_pipe_phv_out_header_8; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_9 = pipe1_io_pipe_phv_out_header_9; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_10 = pipe1_io_pipe_phv_out_header_10; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_11 = pipe1_io_pipe_phv_out_header_11; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_12 = pipe1_io_pipe_phv_out_header_12; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_13 = pipe1_io_pipe_phv_out_header_13; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_14 = pipe1_io_pipe_phv_out_header_14; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_header_15 = pipe1_io_pipe_phv_out_header_15; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_parse_current_state = pipe1_io_pipe_phv_out_parse_current_state; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_parse_current_offset = pipe1_io_pipe_phv_out_parse_current_offset; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_parse_transition_field = pipe1_io_pipe_phv_out_parse_transition_field; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_next_processor_id = pipe1_io_pipe_phv_out_next_processor_id; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_next_config_id = pipe1_io_pipe_phv_out_next_config_id; // @[executor.scala 501:26]
  assign pipe2_io_pipe_phv_in_is_valid_processor = pipe1_io_pipe_phv_out_is_valid_processor; // @[executor.scala 501:26]
  assign pipe2_io_args_in_0 = pipe1_io_args_out_0; // @[executor.scala 502:26]
  assign pipe2_io_args_in_1 = pipe1_io_args_out_1; // @[executor.scala 502:26]
  assign pipe2_io_args_in_2 = pipe1_io_args_out_2; // @[executor.scala 502:26]
  assign pipe2_io_args_in_3 = pipe1_io_args_out_3; // @[executor.scala 502:26]
  assign pipe2_io_args_in_4 = pipe1_io_args_out_4; // @[executor.scala 502:26]
  assign pipe2_io_args_in_5 = pipe1_io_args_out_5; // @[executor.scala 502:26]
  assign pipe2_io_args_in_6 = pipe1_io_args_out_6; // @[executor.scala 502:26]
  assign pipe2_io_vliw_in_0 = pipe1_io_vliw_out_0; // @[executor.scala 503:26]
  assign pipe2_io_vliw_in_1 = pipe1_io_vliw_out_1; // @[executor.scala 503:26]
  assign pipe2_io_vliw_in_2 = pipe1_io_vliw_out_2; // @[executor.scala 503:26]
  assign pipe2_io_vliw_in_3 = pipe1_io_vliw_out_3; // @[executor.scala 503:26]
  assign pipe3_clock = clock;
  assign pipe3_io_pipe_phv_in_data_0 = pipe2_io_pipe_phv_out_data_0; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_1 = pipe2_io_pipe_phv_out_data_1; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_2 = pipe2_io_pipe_phv_out_data_2; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_3 = pipe2_io_pipe_phv_out_data_3; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_4 = pipe2_io_pipe_phv_out_data_4; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_5 = pipe2_io_pipe_phv_out_data_5; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_6 = pipe2_io_pipe_phv_out_data_6; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_7 = pipe2_io_pipe_phv_out_data_7; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_8 = pipe2_io_pipe_phv_out_data_8; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_9 = pipe2_io_pipe_phv_out_data_9; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_10 = pipe2_io_pipe_phv_out_data_10; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_11 = pipe2_io_pipe_phv_out_data_11; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_12 = pipe2_io_pipe_phv_out_data_12; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_13 = pipe2_io_pipe_phv_out_data_13; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_14 = pipe2_io_pipe_phv_out_data_14; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_15 = pipe2_io_pipe_phv_out_data_15; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_16 = pipe2_io_pipe_phv_out_data_16; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_17 = pipe2_io_pipe_phv_out_data_17; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_18 = pipe2_io_pipe_phv_out_data_18; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_19 = pipe2_io_pipe_phv_out_data_19; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_20 = pipe2_io_pipe_phv_out_data_20; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_21 = pipe2_io_pipe_phv_out_data_21; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_22 = pipe2_io_pipe_phv_out_data_22; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_23 = pipe2_io_pipe_phv_out_data_23; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_24 = pipe2_io_pipe_phv_out_data_24; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_25 = pipe2_io_pipe_phv_out_data_25; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_26 = pipe2_io_pipe_phv_out_data_26; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_27 = pipe2_io_pipe_phv_out_data_27; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_28 = pipe2_io_pipe_phv_out_data_28; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_29 = pipe2_io_pipe_phv_out_data_29; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_30 = pipe2_io_pipe_phv_out_data_30; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_31 = pipe2_io_pipe_phv_out_data_31; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_32 = pipe2_io_pipe_phv_out_data_32; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_33 = pipe2_io_pipe_phv_out_data_33; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_34 = pipe2_io_pipe_phv_out_data_34; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_35 = pipe2_io_pipe_phv_out_data_35; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_36 = pipe2_io_pipe_phv_out_data_36; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_37 = pipe2_io_pipe_phv_out_data_37; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_38 = pipe2_io_pipe_phv_out_data_38; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_39 = pipe2_io_pipe_phv_out_data_39; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_40 = pipe2_io_pipe_phv_out_data_40; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_41 = pipe2_io_pipe_phv_out_data_41; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_42 = pipe2_io_pipe_phv_out_data_42; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_43 = pipe2_io_pipe_phv_out_data_43; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_44 = pipe2_io_pipe_phv_out_data_44; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_45 = pipe2_io_pipe_phv_out_data_45; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_46 = pipe2_io_pipe_phv_out_data_46; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_47 = pipe2_io_pipe_phv_out_data_47; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_48 = pipe2_io_pipe_phv_out_data_48; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_49 = pipe2_io_pipe_phv_out_data_49; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_50 = pipe2_io_pipe_phv_out_data_50; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_51 = pipe2_io_pipe_phv_out_data_51; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_52 = pipe2_io_pipe_phv_out_data_52; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_53 = pipe2_io_pipe_phv_out_data_53; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_54 = pipe2_io_pipe_phv_out_data_54; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_55 = pipe2_io_pipe_phv_out_data_55; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_56 = pipe2_io_pipe_phv_out_data_56; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_57 = pipe2_io_pipe_phv_out_data_57; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_58 = pipe2_io_pipe_phv_out_data_58; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_59 = pipe2_io_pipe_phv_out_data_59; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_60 = pipe2_io_pipe_phv_out_data_60; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_61 = pipe2_io_pipe_phv_out_data_61; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_62 = pipe2_io_pipe_phv_out_data_62; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_63 = pipe2_io_pipe_phv_out_data_63; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_64 = pipe2_io_pipe_phv_out_data_64; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_65 = pipe2_io_pipe_phv_out_data_65; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_66 = pipe2_io_pipe_phv_out_data_66; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_67 = pipe2_io_pipe_phv_out_data_67; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_68 = pipe2_io_pipe_phv_out_data_68; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_69 = pipe2_io_pipe_phv_out_data_69; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_70 = pipe2_io_pipe_phv_out_data_70; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_71 = pipe2_io_pipe_phv_out_data_71; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_72 = pipe2_io_pipe_phv_out_data_72; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_73 = pipe2_io_pipe_phv_out_data_73; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_74 = pipe2_io_pipe_phv_out_data_74; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_75 = pipe2_io_pipe_phv_out_data_75; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_76 = pipe2_io_pipe_phv_out_data_76; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_77 = pipe2_io_pipe_phv_out_data_77; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_78 = pipe2_io_pipe_phv_out_data_78; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_79 = pipe2_io_pipe_phv_out_data_79; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_80 = pipe2_io_pipe_phv_out_data_80; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_81 = pipe2_io_pipe_phv_out_data_81; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_82 = pipe2_io_pipe_phv_out_data_82; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_83 = pipe2_io_pipe_phv_out_data_83; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_84 = pipe2_io_pipe_phv_out_data_84; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_85 = pipe2_io_pipe_phv_out_data_85; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_86 = pipe2_io_pipe_phv_out_data_86; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_87 = pipe2_io_pipe_phv_out_data_87; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_88 = pipe2_io_pipe_phv_out_data_88; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_89 = pipe2_io_pipe_phv_out_data_89; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_90 = pipe2_io_pipe_phv_out_data_90; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_91 = pipe2_io_pipe_phv_out_data_91; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_92 = pipe2_io_pipe_phv_out_data_92; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_93 = pipe2_io_pipe_phv_out_data_93; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_94 = pipe2_io_pipe_phv_out_data_94; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_95 = pipe2_io_pipe_phv_out_data_95; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_96 = pipe2_io_pipe_phv_out_data_96; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_97 = pipe2_io_pipe_phv_out_data_97; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_98 = pipe2_io_pipe_phv_out_data_98; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_99 = pipe2_io_pipe_phv_out_data_99; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_100 = pipe2_io_pipe_phv_out_data_100; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_101 = pipe2_io_pipe_phv_out_data_101; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_102 = pipe2_io_pipe_phv_out_data_102; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_103 = pipe2_io_pipe_phv_out_data_103; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_104 = pipe2_io_pipe_phv_out_data_104; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_105 = pipe2_io_pipe_phv_out_data_105; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_106 = pipe2_io_pipe_phv_out_data_106; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_107 = pipe2_io_pipe_phv_out_data_107; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_108 = pipe2_io_pipe_phv_out_data_108; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_109 = pipe2_io_pipe_phv_out_data_109; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_110 = pipe2_io_pipe_phv_out_data_110; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_111 = pipe2_io_pipe_phv_out_data_111; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_112 = pipe2_io_pipe_phv_out_data_112; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_113 = pipe2_io_pipe_phv_out_data_113; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_114 = pipe2_io_pipe_phv_out_data_114; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_115 = pipe2_io_pipe_phv_out_data_115; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_116 = pipe2_io_pipe_phv_out_data_116; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_117 = pipe2_io_pipe_phv_out_data_117; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_118 = pipe2_io_pipe_phv_out_data_118; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_119 = pipe2_io_pipe_phv_out_data_119; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_120 = pipe2_io_pipe_phv_out_data_120; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_121 = pipe2_io_pipe_phv_out_data_121; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_122 = pipe2_io_pipe_phv_out_data_122; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_123 = pipe2_io_pipe_phv_out_data_123; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_124 = pipe2_io_pipe_phv_out_data_124; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_125 = pipe2_io_pipe_phv_out_data_125; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_126 = pipe2_io_pipe_phv_out_data_126; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_127 = pipe2_io_pipe_phv_out_data_127; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_128 = pipe2_io_pipe_phv_out_data_128; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_129 = pipe2_io_pipe_phv_out_data_129; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_130 = pipe2_io_pipe_phv_out_data_130; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_131 = pipe2_io_pipe_phv_out_data_131; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_132 = pipe2_io_pipe_phv_out_data_132; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_133 = pipe2_io_pipe_phv_out_data_133; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_134 = pipe2_io_pipe_phv_out_data_134; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_135 = pipe2_io_pipe_phv_out_data_135; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_136 = pipe2_io_pipe_phv_out_data_136; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_137 = pipe2_io_pipe_phv_out_data_137; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_138 = pipe2_io_pipe_phv_out_data_138; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_139 = pipe2_io_pipe_phv_out_data_139; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_140 = pipe2_io_pipe_phv_out_data_140; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_141 = pipe2_io_pipe_phv_out_data_141; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_142 = pipe2_io_pipe_phv_out_data_142; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_143 = pipe2_io_pipe_phv_out_data_143; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_144 = pipe2_io_pipe_phv_out_data_144; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_145 = pipe2_io_pipe_phv_out_data_145; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_146 = pipe2_io_pipe_phv_out_data_146; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_147 = pipe2_io_pipe_phv_out_data_147; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_148 = pipe2_io_pipe_phv_out_data_148; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_149 = pipe2_io_pipe_phv_out_data_149; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_150 = pipe2_io_pipe_phv_out_data_150; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_151 = pipe2_io_pipe_phv_out_data_151; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_152 = pipe2_io_pipe_phv_out_data_152; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_153 = pipe2_io_pipe_phv_out_data_153; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_154 = pipe2_io_pipe_phv_out_data_154; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_155 = pipe2_io_pipe_phv_out_data_155; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_156 = pipe2_io_pipe_phv_out_data_156; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_157 = pipe2_io_pipe_phv_out_data_157; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_158 = pipe2_io_pipe_phv_out_data_158; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_159 = pipe2_io_pipe_phv_out_data_159; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_160 = pipe2_io_pipe_phv_out_data_160; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_161 = pipe2_io_pipe_phv_out_data_161; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_162 = pipe2_io_pipe_phv_out_data_162; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_163 = pipe2_io_pipe_phv_out_data_163; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_164 = pipe2_io_pipe_phv_out_data_164; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_165 = pipe2_io_pipe_phv_out_data_165; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_166 = pipe2_io_pipe_phv_out_data_166; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_167 = pipe2_io_pipe_phv_out_data_167; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_168 = pipe2_io_pipe_phv_out_data_168; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_169 = pipe2_io_pipe_phv_out_data_169; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_170 = pipe2_io_pipe_phv_out_data_170; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_171 = pipe2_io_pipe_phv_out_data_171; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_172 = pipe2_io_pipe_phv_out_data_172; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_173 = pipe2_io_pipe_phv_out_data_173; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_174 = pipe2_io_pipe_phv_out_data_174; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_175 = pipe2_io_pipe_phv_out_data_175; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_176 = pipe2_io_pipe_phv_out_data_176; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_177 = pipe2_io_pipe_phv_out_data_177; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_178 = pipe2_io_pipe_phv_out_data_178; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_179 = pipe2_io_pipe_phv_out_data_179; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_180 = pipe2_io_pipe_phv_out_data_180; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_181 = pipe2_io_pipe_phv_out_data_181; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_182 = pipe2_io_pipe_phv_out_data_182; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_183 = pipe2_io_pipe_phv_out_data_183; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_184 = pipe2_io_pipe_phv_out_data_184; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_185 = pipe2_io_pipe_phv_out_data_185; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_186 = pipe2_io_pipe_phv_out_data_186; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_187 = pipe2_io_pipe_phv_out_data_187; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_188 = pipe2_io_pipe_phv_out_data_188; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_189 = pipe2_io_pipe_phv_out_data_189; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_190 = pipe2_io_pipe_phv_out_data_190; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_191 = pipe2_io_pipe_phv_out_data_191; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_192 = pipe2_io_pipe_phv_out_data_192; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_193 = pipe2_io_pipe_phv_out_data_193; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_194 = pipe2_io_pipe_phv_out_data_194; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_195 = pipe2_io_pipe_phv_out_data_195; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_196 = pipe2_io_pipe_phv_out_data_196; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_197 = pipe2_io_pipe_phv_out_data_197; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_198 = pipe2_io_pipe_phv_out_data_198; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_199 = pipe2_io_pipe_phv_out_data_199; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_200 = pipe2_io_pipe_phv_out_data_200; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_201 = pipe2_io_pipe_phv_out_data_201; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_202 = pipe2_io_pipe_phv_out_data_202; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_203 = pipe2_io_pipe_phv_out_data_203; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_204 = pipe2_io_pipe_phv_out_data_204; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_205 = pipe2_io_pipe_phv_out_data_205; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_206 = pipe2_io_pipe_phv_out_data_206; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_207 = pipe2_io_pipe_phv_out_data_207; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_208 = pipe2_io_pipe_phv_out_data_208; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_209 = pipe2_io_pipe_phv_out_data_209; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_210 = pipe2_io_pipe_phv_out_data_210; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_211 = pipe2_io_pipe_phv_out_data_211; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_212 = pipe2_io_pipe_phv_out_data_212; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_213 = pipe2_io_pipe_phv_out_data_213; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_214 = pipe2_io_pipe_phv_out_data_214; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_215 = pipe2_io_pipe_phv_out_data_215; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_216 = pipe2_io_pipe_phv_out_data_216; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_217 = pipe2_io_pipe_phv_out_data_217; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_218 = pipe2_io_pipe_phv_out_data_218; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_219 = pipe2_io_pipe_phv_out_data_219; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_220 = pipe2_io_pipe_phv_out_data_220; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_221 = pipe2_io_pipe_phv_out_data_221; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_222 = pipe2_io_pipe_phv_out_data_222; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_223 = pipe2_io_pipe_phv_out_data_223; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_224 = pipe2_io_pipe_phv_out_data_224; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_225 = pipe2_io_pipe_phv_out_data_225; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_226 = pipe2_io_pipe_phv_out_data_226; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_227 = pipe2_io_pipe_phv_out_data_227; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_228 = pipe2_io_pipe_phv_out_data_228; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_229 = pipe2_io_pipe_phv_out_data_229; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_230 = pipe2_io_pipe_phv_out_data_230; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_231 = pipe2_io_pipe_phv_out_data_231; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_232 = pipe2_io_pipe_phv_out_data_232; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_233 = pipe2_io_pipe_phv_out_data_233; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_234 = pipe2_io_pipe_phv_out_data_234; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_235 = pipe2_io_pipe_phv_out_data_235; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_236 = pipe2_io_pipe_phv_out_data_236; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_237 = pipe2_io_pipe_phv_out_data_237; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_238 = pipe2_io_pipe_phv_out_data_238; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_239 = pipe2_io_pipe_phv_out_data_239; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_240 = pipe2_io_pipe_phv_out_data_240; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_241 = pipe2_io_pipe_phv_out_data_241; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_242 = pipe2_io_pipe_phv_out_data_242; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_243 = pipe2_io_pipe_phv_out_data_243; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_244 = pipe2_io_pipe_phv_out_data_244; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_245 = pipe2_io_pipe_phv_out_data_245; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_246 = pipe2_io_pipe_phv_out_data_246; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_247 = pipe2_io_pipe_phv_out_data_247; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_248 = pipe2_io_pipe_phv_out_data_248; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_249 = pipe2_io_pipe_phv_out_data_249; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_250 = pipe2_io_pipe_phv_out_data_250; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_251 = pipe2_io_pipe_phv_out_data_251; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_252 = pipe2_io_pipe_phv_out_data_252; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_253 = pipe2_io_pipe_phv_out_data_253; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_254 = pipe2_io_pipe_phv_out_data_254; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_255 = pipe2_io_pipe_phv_out_data_255; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_256 = pipe2_io_pipe_phv_out_data_256; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_257 = pipe2_io_pipe_phv_out_data_257; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_258 = pipe2_io_pipe_phv_out_data_258; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_259 = pipe2_io_pipe_phv_out_data_259; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_260 = pipe2_io_pipe_phv_out_data_260; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_261 = pipe2_io_pipe_phv_out_data_261; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_262 = pipe2_io_pipe_phv_out_data_262; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_263 = pipe2_io_pipe_phv_out_data_263; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_264 = pipe2_io_pipe_phv_out_data_264; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_265 = pipe2_io_pipe_phv_out_data_265; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_266 = pipe2_io_pipe_phv_out_data_266; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_267 = pipe2_io_pipe_phv_out_data_267; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_268 = pipe2_io_pipe_phv_out_data_268; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_269 = pipe2_io_pipe_phv_out_data_269; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_270 = pipe2_io_pipe_phv_out_data_270; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_271 = pipe2_io_pipe_phv_out_data_271; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_272 = pipe2_io_pipe_phv_out_data_272; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_273 = pipe2_io_pipe_phv_out_data_273; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_274 = pipe2_io_pipe_phv_out_data_274; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_275 = pipe2_io_pipe_phv_out_data_275; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_276 = pipe2_io_pipe_phv_out_data_276; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_277 = pipe2_io_pipe_phv_out_data_277; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_278 = pipe2_io_pipe_phv_out_data_278; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_279 = pipe2_io_pipe_phv_out_data_279; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_280 = pipe2_io_pipe_phv_out_data_280; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_281 = pipe2_io_pipe_phv_out_data_281; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_282 = pipe2_io_pipe_phv_out_data_282; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_283 = pipe2_io_pipe_phv_out_data_283; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_284 = pipe2_io_pipe_phv_out_data_284; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_285 = pipe2_io_pipe_phv_out_data_285; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_286 = pipe2_io_pipe_phv_out_data_286; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_287 = pipe2_io_pipe_phv_out_data_287; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_288 = pipe2_io_pipe_phv_out_data_288; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_289 = pipe2_io_pipe_phv_out_data_289; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_290 = pipe2_io_pipe_phv_out_data_290; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_291 = pipe2_io_pipe_phv_out_data_291; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_292 = pipe2_io_pipe_phv_out_data_292; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_293 = pipe2_io_pipe_phv_out_data_293; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_294 = pipe2_io_pipe_phv_out_data_294; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_295 = pipe2_io_pipe_phv_out_data_295; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_296 = pipe2_io_pipe_phv_out_data_296; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_297 = pipe2_io_pipe_phv_out_data_297; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_298 = pipe2_io_pipe_phv_out_data_298; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_299 = pipe2_io_pipe_phv_out_data_299; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_300 = pipe2_io_pipe_phv_out_data_300; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_301 = pipe2_io_pipe_phv_out_data_301; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_302 = pipe2_io_pipe_phv_out_data_302; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_303 = pipe2_io_pipe_phv_out_data_303; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_304 = pipe2_io_pipe_phv_out_data_304; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_305 = pipe2_io_pipe_phv_out_data_305; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_306 = pipe2_io_pipe_phv_out_data_306; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_307 = pipe2_io_pipe_phv_out_data_307; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_308 = pipe2_io_pipe_phv_out_data_308; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_309 = pipe2_io_pipe_phv_out_data_309; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_310 = pipe2_io_pipe_phv_out_data_310; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_311 = pipe2_io_pipe_phv_out_data_311; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_312 = pipe2_io_pipe_phv_out_data_312; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_313 = pipe2_io_pipe_phv_out_data_313; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_314 = pipe2_io_pipe_phv_out_data_314; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_315 = pipe2_io_pipe_phv_out_data_315; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_316 = pipe2_io_pipe_phv_out_data_316; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_317 = pipe2_io_pipe_phv_out_data_317; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_318 = pipe2_io_pipe_phv_out_data_318; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_319 = pipe2_io_pipe_phv_out_data_319; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_320 = pipe2_io_pipe_phv_out_data_320; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_321 = pipe2_io_pipe_phv_out_data_321; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_322 = pipe2_io_pipe_phv_out_data_322; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_323 = pipe2_io_pipe_phv_out_data_323; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_324 = pipe2_io_pipe_phv_out_data_324; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_325 = pipe2_io_pipe_phv_out_data_325; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_326 = pipe2_io_pipe_phv_out_data_326; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_327 = pipe2_io_pipe_phv_out_data_327; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_328 = pipe2_io_pipe_phv_out_data_328; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_329 = pipe2_io_pipe_phv_out_data_329; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_330 = pipe2_io_pipe_phv_out_data_330; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_331 = pipe2_io_pipe_phv_out_data_331; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_332 = pipe2_io_pipe_phv_out_data_332; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_333 = pipe2_io_pipe_phv_out_data_333; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_334 = pipe2_io_pipe_phv_out_data_334; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_335 = pipe2_io_pipe_phv_out_data_335; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_336 = pipe2_io_pipe_phv_out_data_336; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_337 = pipe2_io_pipe_phv_out_data_337; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_338 = pipe2_io_pipe_phv_out_data_338; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_339 = pipe2_io_pipe_phv_out_data_339; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_340 = pipe2_io_pipe_phv_out_data_340; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_341 = pipe2_io_pipe_phv_out_data_341; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_342 = pipe2_io_pipe_phv_out_data_342; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_343 = pipe2_io_pipe_phv_out_data_343; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_344 = pipe2_io_pipe_phv_out_data_344; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_345 = pipe2_io_pipe_phv_out_data_345; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_346 = pipe2_io_pipe_phv_out_data_346; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_347 = pipe2_io_pipe_phv_out_data_347; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_348 = pipe2_io_pipe_phv_out_data_348; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_349 = pipe2_io_pipe_phv_out_data_349; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_350 = pipe2_io_pipe_phv_out_data_350; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_351 = pipe2_io_pipe_phv_out_data_351; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_352 = pipe2_io_pipe_phv_out_data_352; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_353 = pipe2_io_pipe_phv_out_data_353; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_354 = pipe2_io_pipe_phv_out_data_354; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_355 = pipe2_io_pipe_phv_out_data_355; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_356 = pipe2_io_pipe_phv_out_data_356; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_357 = pipe2_io_pipe_phv_out_data_357; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_358 = pipe2_io_pipe_phv_out_data_358; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_359 = pipe2_io_pipe_phv_out_data_359; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_360 = pipe2_io_pipe_phv_out_data_360; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_361 = pipe2_io_pipe_phv_out_data_361; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_362 = pipe2_io_pipe_phv_out_data_362; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_363 = pipe2_io_pipe_phv_out_data_363; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_364 = pipe2_io_pipe_phv_out_data_364; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_365 = pipe2_io_pipe_phv_out_data_365; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_366 = pipe2_io_pipe_phv_out_data_366; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_367 = pipe2_io_pipe_phv_out_data_367; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_368 = pipe2_io_pipe_phv_out_data_368; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_369 = pipe2_io_pipe_phv_out_data_369; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_370 = pipe2_io_pipe_phv_out_data_370; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_371 = pipe2_io_pipe_phv_out_data_371; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_372 = pipe2_io_pipe_phv_out_data_372; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_373 = pipe2_io_pipe_phv_out_data_373; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_374 = pipe2_io_pipe_phv_out_data_374; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_375 = pipe2_io_pipe_phv_out_data_375; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_376 = pipe2_io_pipe_phv_out_data_376; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_377 = pipe2_io_pipe_phv_out_data_377; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_378 = pipe2_io_pipe_phv_out_data_378; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_379 = pipe2_io_pipe_phv_out_data_379; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_380 = pipe2_io_pipe_phv_out_data_380; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_381 = pipe2_io_pipe_phv_out_data_381; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_382 = pipe2_io_pipe_phv_out_data_382; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_383 = pipe2_io_pipe_phv_out_data_383; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_384 = pipe2_io_pipe_phv_out_data_384; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_385 = pipe2_io_pipe_phv_out_data_385; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_386 = pipe2_io_pipe_phv_out_data_386; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_387 = pipe2_io_pipe_phv_out_data_387; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_388 = pipe2_io_pipe_phv_out_data_388; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_389 = pipe2_io_pipe_phv_out_data_389; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_390 = pipe2_io_pipe_phv_out_data_390; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_391 = pipe2_io_pipe_phv_out_data_391; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_392 = pipe2_io_pipe_phv_out_data_392; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_393 = pipe2_io_pipe_phv_out_data_393; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_394 = pipe2_io_pipe_phv_out_data_394; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_395 = pipe2_io_pipe_phv_out_data_395; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_396 = pipe2_io_pipe_phv_out_data_396; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_397 = pipe2_io_pipe_phv_out_data_397; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_398 = pipe2_io_pipe_phv_out_data_398; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_399 = pipe2_io_pipe_phv_out_data_399; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_400 = pipe2_io_pipe_phv_out_data_400; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_401 = pipe2_io_pipe_phv_out_data_401; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_402 = pipe2_io_pipe_phv_out_data_402; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_403 = pipe2_io_pipe_phv_out_data_403; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_404 = pipe2_io_pipe_phv_out_data_404; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_405 = pipe2_io_pipe_phv_out_data_405; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_406 = pipe2_io_pipe_phv_out_data_406; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_407 = pipe2_io_pipe_phv_out_data_407; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_408 = pipe2_io_pipe_phv_out_data_408; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_409 = pipe2_io_pipe_phv_out_data_409; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_410 = pipe2_io_pipe_phv_out_data_410; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_411 = pipe2_io_pipe_phv_out_data_411; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_412 = pipe2_io_pipe_phv_out_data_412; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_413 = pipe2_io_pipe_phv_out_data_413; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_414 = pipe2_io_pipe_phv_out_data_414; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_415 = pipe2_io_pipe_phv_out_data_415; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_416 = pipe2_io_pipe_phv_out_data_416; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_417 = pipe2_io_pipe_phv_out_data_417; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_418 = pipe2_io_pipe_phv_out_data_418; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_419 = pipe2_io_pipe_phv_out_data_419; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_420 = pipe2_io_pipe_phv_out_data_420; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_421 = pipe2_io_pipe_phv_out_data_421; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_422 = pipe2_io_pipe_phv_out_data_422; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_423 = pipe2_io_pipe_phv_out_data_423; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_424 = pipe2_io_pipe_phv_out_data_424; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_425 = pipe2_io_pipe_phv_out_data_425; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_426 = pipe2_io_pipe_phv_out_data_426; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_427 = pipe2_io_pipe_phv_out_data_427; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_428 = pipe2_io_pipe_phv_out_data_428; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_429 = pipe2_io_pipe_phv_out_data_429; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_430 = pipe2_io_pipe_phv_out_data_430; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_431 = pipe2_io_pipe_phv_out_data_431; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_432 = pipe2_io_pipe_phv_out_data_432; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_433 = pipe2_io_pipe_phv_out_data_433; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_434 = pipe2_io_pipe_phv_out_data_434; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_435 = pipe2_io_pipe_phv_out_data_435; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_436 = pipe2_io_pipe_phv_out_data_436; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_437 = pipe2_io_pipe_phv_out_data_437; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_438 = pipe2_io_pipe_phv_out_data_438; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_439 = pipe2_io_pipe_phv_out_data_439; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_440 = pipe2_io_pipe_phv_out_data_440; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_441 = pipe2_io_pipe_phv_out_data_441; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_442 = pipe2_io_pipe_phv_out_data_442; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_443 = pipe2_io_pipe_phv_out_data_443; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_444 = pipe2_io_pipe_phv_out_data_444; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_445 = pipe2_io_pipe_phv_out_data_445; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_446 = pipe2_io_pipe_phv_out_data_446; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_447 = pipe2_io_pipe_phv_out_data_447; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_448 = pipe2_io_pipe_phv_out_data_448; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_449 = pipe2_io_pipe_phv_out_data_449; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_450 = pipe2_io_pipe_phv_out_data_450; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_451 = pipe2_io_pipe_phv_out_data_451; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_452 = pipe2_io_pipe_phv_out_data_452; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_453 = pipe2_io_pipe_phv_out_data_453; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_454 = pipe2_io_pipe_phv_out_data_454; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_455 = pipe2_io_pipe_phv_out_data_455; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_456 = pipe2_io_pipe_phv_out_data_456; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_457 = pipe2_io_pipe_phv_out_data_457; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_458 = pipe2_io_pipe_phv_out_data_458; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_459 = pipe2_io_pipe_phv_out_data_459; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_460 = pipe2_io_pipe_phv_out_data_460; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_461 = pipe2_io_pipe_phv_out_data_461; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_462 = pipe2_io_pipe_phv_out_data_462; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_463 = pipe2_io_pipe_phv_out_data_463; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_464 = pipe2_io_pipe_phv_out_data_464; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_465 = pipe2_io_pipe_phv_out_data_465; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_466 = pipe2_io_pipe_phv_out_data_466; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_467 = pipe2_io_pipe_phv_out_data_467; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_468 = pipe2_io_pipe_phv_out_data_468; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_469 = pipe2_io_pipe_phv_out_data_469; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_470 = pipe2_io_pipe_phv_out_data_470; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_471 = pipe2_io_pipe_phv_out_data_471; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_472 = pipe2_io_pipe_phv_out_data_472; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_473 = pipe2_io_pipe_phv_out_data_473; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_474 = pipe2_io_pipe_phv_out_data_474; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_475 = pipe2_io_pipe_phv_out_data_475; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_476 = pipe2_io_pipe_phv_out_data_476; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_477 = pipe2_io_pipe_phv_out_data_477; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_478 = pipe2_io_pipe_phv_out_data_478; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_479 = pipe2_io_pipe_phv_out_data_479; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_480 = pipe2_io_pipe_phv_out_data_480; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_481 = pipe2_io_pipe_phv_out_data_481; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_482 = pipe2_io_pipe_phv_out_data_482; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_483 = pipe2_io_pipe_phv_out_data_483; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_484 = pipe2_io_pipe_phv_out_data_484; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_485 = pipe2_io_pipe_phv_out_data_485; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_486 = pipe2_io_pipe_phv_out_data_486; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_487 = pipe2_io_pipe_phv_out_data_487; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_488 = pipe2_io_pipe_phv_out_data_488; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_489 = pipe2_io_pipe_phv_out_data_489; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_490 = pipe2_io_pipe_phv_out_data_490; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_491 = pipe2_io_pipe_phv_out_data_491; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_492 = pipe2_io_pipe_phv_out_data_492; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_493 = pipe2_io_pipe_phv_out_data_493; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_494 = pipe2_io_pipe_phv_out_data_494; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_495 = pipe2_io_pipe_phv_out_data_495; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_496 = pipe2_io_pipe_phv_out_data_496; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_497 = pipe2_io_pipe_phv_out_data_497; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_498 = pipe2_io_pipe_phv_out_data_498; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_499 = pipe2_io_pipe_phv_out_data_499; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_500 = pipe2_io_pipe_phv_out_data_500; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_501 = pipe2_io_pipe_phv_out_data_501; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_502 = pipe2_io_pipe_phv_out_data_502; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_503 = pipe2_io_pipe_phv_out_data_503; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_504 = pipe2_io_pipe_phv_out_data_504; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_505 = pipe2_io_pipe_phv_out_data_505; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_506 = pipe2_io_pipe_phv_out_data_506; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_507 = pipe2_io_pipe_phv_out_data_507; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_508 = pipe2_io_pipe_phv_out_data_508; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_509 = pipe2_io_pipe_phv_out_data_509; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_510 = pipe2_io_pipe_phv_out_data_510; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_data_511 = pipe2_io_pipe_phv_out_data_511; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_0 = pipe2_io_pipe_phv_out_header_0; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_1 = pipe2_io_pipe_phv_out_header_1; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_2 = pipe2_io_pipe_phv_out_header_2; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_3 = pipe2_io_pipe_phv_out_header_3; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_4 = pipe2_io_pipe_phv_out_header_4; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_5 = pipe2_io_pipe_phv_out_header_5; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_6 = pipe2_io_pipe_phv_out_header_6; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_7 = pipe2_io_pipe_phv_out_header_7; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_8 = pipe2_io_pipe_phv_out_header_8; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_9 = pipe2_io_pipe_phv_out_header_9; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_10 = pipe2_io_pipe_phv_out_header_10; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_11 = pipe2_io_pipe_phv_out_header_11; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_12 = pipe2_io_pipe_phv_out_header_12; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_13 = pipe2_io_pipe_phv_out_header_13; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_14 = pipe2_io_pipe_phv_out_header_14; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_header_15 = pipe2_io_pipe_phv_out_header_15; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_parse_current_state = pipe2_io_pipe_phv_out_parse_current_state; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_parse_current_offset = pipe2_io_pipe_phv_out_parse_current_offset; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_parse_transition_field = pipe2_io_pipe_phv_out_parse_transition_field; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_next_processor_id = pipe2_io_pipe_phv_out_next_processor_id; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_next_config_id = pipe2_io_pipe_phv_out_next_config_id; // @[executor.scala 505:26]
  assign pipe3_io_pipe_phv_in_is_valid_processor = pipe2_io_pipe_phv_out_is_valid_processor; // @[executor.scala 505:26]
  assign pipe3_io_args_in_0 = pipe2_io_args_out_0; // @[executor.scala 506:26]
  assign pipe3_io_args_in_1 = pipe2_io_args_out_1; // @[executor.scala 506:26]
  assign pipe3_io_args_in_2 = pipe2_io_args_out_2; // @[executor.scala 506:26]
  assign pipe3_io_args_in_3 = pipe2_io_args_out_3; // @[executor.scala 506:26]
  assign pipe3_io_args_in_4 = pipe2_io_args_out_4; // @[executor.scala 506:26]
  assign pipe3_io_args_in_5 = pipe2_io_args_out_5; // @[executor.scala 506:26]
  assign pipe3_io_args_in_6 = pipe2_io_args_out_6; // @[executor.scala 506:26]
  assign pipe3_io_vliw_in_0 = pipe2_io_vliw_out_0; // @[executor.scala 507:26]
  assign pipe3_io_vliw_in_1 = pipe2_io_vliw_out_1; // @[executor.scala 507:26]
  assign pipe3_io_vliw_in_2 = pipe2_io_vliw_out_2; // @[executor.scala 507:26]
  assign pipe3_io_vliw_in_3 = pipe2_io_vliw_out_3; // @[executor.scala 507:26]
  assign pipe3_io_offset_in_0 = pipe2_io_offset_out_0; // @[executor.scala 508:26]
  assign pipe3_io_offset_in_1 = pipe2_io_offset_out_1; // @[executor.scala 508:26]
  assign pipe3_io_offset_in_2 = pipe2_io_offset_out_2; // @[executor.scala 508:26]
  assign pipe3_io_offset_in_3 = pipe2_io_offset_out_3; // @[executor.scala 508:26]
  assign pipe3_io_length_in_0 = pipe2_io_length_out_0; // @[executor.scala 509:26]
  assign pipe3_io_length_in_1 = pipe2_io_length_out_1; // @[executor.scala 509:26]
  assign pipe3_io_length_in_2 = pipe2_io_length_out_2; // @[executor.scala 509:26]
  assign pipe3_io_length_in_3 = pipe2_io_length_out_3; // @[executor.scala 509:26]
  assign pipe4_clock = clock;
  assign pipe4_io_pipe_phv_in_data_0 = pipe3_io_pipe_phv_out_data_0; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_1 = pipe3_io_pipe_phv_out_data_1; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_2 = pipe3_io_pipe_phv_out_data_2; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_3 = pipe3_io_pipe_phv_out_data_3; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_4 = pipe3_io_pipe_phv_out_data_4; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_5 = pipe3_io_pipe_phv_out_data_5; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_6 = pipe3_io_pipe_phv_out_data_6; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_7 = pipe3_io_pipe_phv_out_data_7; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_8 = pipe3_io_pipe_phv_out_data_8; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_9 = pipe3_io_pipe_phv_out_data_9; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_10 = pipe3_io_pipe_phv_out_data_10; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_11 = pipe3_io_pipe_phv_out_data_11; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_12 = pipe3_io_pipe_phv_out_data_12; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_13 = pipe3_io_pipe_phv_out_data_13; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_14 = pipe3_io_pipe_phv_out_data_14; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_15 = pipe3_io_pipe_phv_out_data_15; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_16 = pipe3_io_pipe_phv_out_data_16; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_17 = pipe3_io_pipe_phv_out_data_17; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_18 = pipe3_io_pipe_phv_out_data_18; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_19 = pipe3_io_pipe_phv_out_data_19; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_20 = pipe3_io_pipe_phv_out_data_20; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_21 = pipe3_io_pipe_phv_out_data_21; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_22 = pipe3_io_pipe_phv_out_data_22; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_23 = pipe3_io_pipe_phv_out_data_23; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_24 = pipe3_io_pipe_phv_out_data_24; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_25 = pipe3_io_pipe_phv_out_data_25; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_26 = pipe3_io_pipe_phv_out_data_26; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_27 = pipe3_io_pipe_phv_out_data_27; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_28 = pipe3_io_pipe_phv_out_data_28; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_29 = pipe3_io_pipe_phv_out_data_29; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_30 = pipe3_io_pipe_phv_out_data_30; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_31 = pipe3_io_pipe_phv_out_data_31; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_32 = pipe3_io_pipe_phv_out_data_32; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_33 = pipe3_io_pipe_phv_out_data_33; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_34 = pipe3_io_pipe_phv_out_data_34; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_35 = pipe3_io_pipe_phv_out_data_35; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_36 = pipe3_io_pipe_phv_out_data_36; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_37 = pipe3_io_pipe_phv_out_data_37; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_38 = pipe3_io_pipe_phv_out_data_38; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_39 = pipe3_io_pipe_phv_out_data_39; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_40 = pipe3_io_pipe_phv_out_data_40; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_41 = pipe3_io_pipe_phv_out_data_41; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_42 = pipe3_io_pipe_phv_out_data_42; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_43 = pipe3_io_pipe_phv_out_data_43; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_44 = pipe3_io_pipe_phv_out_data_44; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_45 = pipe3_io_pipe_phv_out_data_45; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_46 = pipe3_io_pipe_phv_out_data_46; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_47 = pipe3_io_pipe_phv_out_data_47; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_48 = pipe3_io_pipe_phv_out_data_48; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_49 = pipe3_io_pipe_phv_out_data_49; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_50 = pipe3_io_pipe_phv_out_data_50; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_51 = pipe3_io_pipe_phv_out_data_51; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_52 = pipe3_io_pipe_phv_out_data_52; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_53 = pipe3_io_pipe_phv_out_data_53; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_54 = pipe3_io_pipe_phv_out_data_54; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_55 = pipe3_io_pipe_phv_out_data_55; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_56 = pipe3_io_pipe_phv_out_data_56; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_57 = pipe3_io_pipe_phv_out_data_57; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_58 = pipe3_io_pipe_phv_out_data_58; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_59 = pipe3_io_pipe_phv_out_data_59; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_60 = pipe3_io_pipe_phv_out_data_60; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_61 = pipe3_io_pipe_phv_out_data_61; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_62 = pipe3_io_pipe_phv_out_data_62; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_63 = pipe3_io_pipe_phv_out_data_63; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_64 = pipe3_io_pipe_phv_out_data_64; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_65 = pipe3_io_pipe_phv_out_data_65; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_66 = pipe3_io_pipe_phv_out_data_66; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_67 = pipe3_io_pipe_phv_out_data_67; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_68 = pipe3_io_pipe_phv_out_data_68; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_69 = pipe3_io_pipe_phv_out_data_69; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_70 = pipe3_io_pipe_phv_out_data_70; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_71 = pipe3_io_pipe_phv_out_data_71; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_72 = pipe3_io_pipe_phv_out_data_72; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_73 = pipe3_io_pipe_phv_out_data_73; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_74 = pipe3_io_pipe_phv_out_data_74; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_75 = pipe3_io_pipe_phv_out_data_75; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_76 = pipe3_io_pipe_phv_out_data_76; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_77 = pipe3_io_pipe_phv_out_data_77; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_78 = pipe3_io_pipe_phv_out_data_78; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_79 = pipe3_io_pipe_phv_out_data_79; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_80 = pipe3_io_pipe_phv_out_data_80; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_81 = pipe3_io_pipe_phv_out_data_81; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_82 = pipe3_io_pipe_phv_out_data_82; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_83 = pipe3_io_pipe_phv_out_data_83; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_84 = pipe3_io_pipe_phv_out_data_84; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_85 = pipe3_io_pipe_phv_out_data_85; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_86 = pipe3_io_pipe_phv_out_data_86; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_87 = pipe3_io_pipe_phv_out_data_87; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_88 = pipe3_io_pipe_phv_out_data_88; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_89 = pipe3_io_pipe_phv_out_data_89; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_90 = pipe3_io_pipe_phv_out_data_90; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_91 = pipe3_io_pipe_phv_out_data_91; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_92 = pipe3_io_pipe_phv_out_data_92; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_93 = pipe3_io_pipe_phv_out_data_93; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_94 = pipe3_io_pipe_phv_out_data_94; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_95 = pipe3_io_pipe_phv_out_data_95; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_96 = pipe3_io_pipe_phv_out_data_96; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_97 = pipe3_io_pipe_phv_out_data_97; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_98 = pipe3_io_pipe_phv_out_data_98; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_99 = pipe3_io_pipe_phv_out_data_99; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_100 = pipe3_io_pipe_phv_out_data_100; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_101 = pipe3_io_pipe_phv_out_data_101; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_102 = pipe3_io_pipe_phv_out_data_102; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_103 = pipe3_io_pipe_phv_out_data_103; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_104 = pipe3_io_pipe_phv_out_data_104; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_105 = pipe3_io_pipe_phv_out_data_105; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_106 = pipe3_io_pipe_phv_out_data_106; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_107 = pipe3_io_pipe_phv_out_data_107; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_108 = pipe3_io_pipe_phv_out_data_108; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_109 = pipe3_io_pipe_phv_out_data_109; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_110 = pipe3_io_pipe_phv_out_data_110; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_111 = pipe3_io_pipe_phv_out_data_111; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_112 = pipe3_io_pipe_phv_out_data_112; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_113 = pipe3_io_pipe_phv_out_data_113; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_114 = pipe3_io_pipe_phv_out_data_114; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_115 = pipe3_io_pipe_phv_out_data_115; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_116 = pipe3_io_pipe_phv_out_data_116; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_117 = pipe3_io_pipe_phv_out_data_117; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_118 = pipe3_io_pipe_phv_out_data_118; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_119 = pipe3_io_pipe_phv_out_data_119; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_120 = pipe3_io_pipe_phv_out_data_120; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_121 = pipe3_io_pipe_phv_out_data_121; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_122 = pipe3_io_pipe_phv_out_data_122; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_123 = pipe3_io_pipe_phv_out_data_123; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_124 = pipe3_io_pipe_phv_out_data_124; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_125 = pipe3_io_pipe_phv_out_data_125; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_126 = pipe3_io_pipe_phv_out_data_126; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_127 = pipe3_io_pipe_phv_out_data_127; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_128 = pipe3_io_pipe_phv_out_data_128; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_129 = pipe3_io_pipe_phv_out_data_129; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_130 = pipe3_io_pipe_phv_out_data_130; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_131 = pipe3_io_pipe_phv_out_data_131; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_132 = pipe3_io_pipe_phv_out_data_132; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_133 = pipe3_io_pipe_phv_out_data_133; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_134 = pipe3_io_pipe_phv_out_data_134; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_135 = pipe3_io_pipe_phv_out_data_135; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_136 = pipe3_io_pipe_phv_out_data_136; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_137 = pipe3_io_pipe_phv_out_data_137; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_138 = pipe3_io_pipe_phv_out_data_138; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_139 = pipe3_io_pipe_phv_out_data_139; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_140 = pipe3_io_pipe_phv_out_data_140; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_141 = pipe3_io_pipe_phv_out_data_141; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_142 = pipe3_io_pipe_phv_out_data_142; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_143 = pipe3_io_pipe_phv_out_data_143; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_144 = pipe3_io_pipe_phv_out_data_144; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_145 = pipe3_io_pipe_phv_out_data_145; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_146 = pipe3_io_pipe_phv_out_data_146; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_147 = pipe3_io_pipe_phv_out_data_147; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_148 = pipe3_io_pipe_phv_out_data_148; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_149 = pipe3_io_pipe_phv_out_data_149; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_150 = pipe3_io_pipe_phv_out_data_150; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_151 = pipe3_io_pipe_phv_out_data_151; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_152 = pipe3_io_pipe_phv_out_data_152; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_153 = pipe3_io_pipe_phv_out_data_153; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_154 = pipe3_io_pipe_phv_out_data_154; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_155 = pipe3_io_pipe_phv_out_data_155; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_156 = pipe3_io_pipe_phv_out_data_156; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_157 = pipe3_io_pipe_phv_out_data_157; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_158 = pipe3_io_pipe_phv_out_data_158; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_159 = pipe3_io_pipe_phv_out_data_159; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_160 = pipe3_io_pipe_phv_out_data_160; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_161 = pipe3_io_pipe_phv_out_data_161; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_162 = pipe3_io_pipe_phv_out_data_162; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_163 = pipe3_io_pipe_phv_out_data_163; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_164 = pipe3_io_pipe_phv_out_data_164; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_165 = pipe3_io_pipe_phv_out_data_165; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_166 = pipe3_io_pipe_phv_out_data_166; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_167 = pipe3_io_pipe_phv_out_data_167; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_168 = pipe3_io_pipe_phv_out_data_168; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_169 = pipe3_io_pipe_phv_out_data_169; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_170 = pipe3_io_pipe_phv_out_data_170; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_171 = pipe3_io_pipe_phv_out_data_171; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_172 = pipe3_io_pipe_phv_out_data_172; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_173 = pipe3_io_pipe_phv_out_data_173; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_174 = pipe3_io_pipe_phv_out_data_174; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_175 = pipe3_io_pipe_phv_out_data_175; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_176 = pipe3_io_pipe_phv_out_data_176; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_177 = pipe3_io_pipe_phv_out_data_177; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_178 = pipe3_io_pipe_phv_out_data_178; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_179 = pipe3_io_pipe_phv_out_data_179; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_180 = pipe3_io_pipe_phv_out_data_180; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_181 = pipe3_io_pipe_phv_out_data_181; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_182 = pipe3_io_pipe_phv_out_data_182; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_183 = pipe3_io_pipe_phv_out_data_183; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_184 = pipe3_io_pipe_phv_out_data_184; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_185 = pipe3_io_pipe_phv_out_data_185; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_186 = pipe3_io_pipe_phv_out_data_186; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_187 = pipe3_io_pipe_phv_out_data_187; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_188 = pipe3_io_pipe_phv_out_data_188; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_189 = pipe3_io_pipe_phv_out_data_189; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_190 = pipe3_io_pipe_phv_out_data_190; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_191 = pipe3_io_pipe_phv_out_data_191; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_192 = pipe3_io_pipe_phv_out_data_192; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_193 = pipe3_io_pipe_phv_out_data_193; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_194 = pipe3_io_pipe_phv_out_data_194; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_195 = pipe3_io_pipe_phv_out_data_195; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_196 = pipe3_io_pipe_phv_out_data_196; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_197 = pipe3_io_pipe_phv_out_data_197; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_198 = pipe3_io_pipe_phv_out_data_198; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_199 = pipe3_io_pipe_phv_out_data_199; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_200 = pipe3_io_pipe_phv_out_data_200; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_201 = pipe3_io_pipe_phv_out_data_201; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_202 = pipe3_io_pipe_phv_out_data_202; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_203 = pipe3_io_pipe_phv_out_data_203; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_204 = pipe3_io_pipe_phv_out_data_204; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_205 = pipe3_io_pipe_phv_out_data_205; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_206 = pipe3_io_pipe_phv_out_data_206; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_207 = pipe3_io_pipe_phv_out_data_207; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_208 = pipe3_io_pipe_phv_out_data_208; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_209 = pipe3_io_pipe_phv_out_data_209; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_210 = pipe3_io_pipe_phv_out_data_210; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_211 = pipe3_io_pipe_phv_out_data_211; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_212 = pipe3_io_pipe_phv_out_data_212; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_213 = pipe3_io_pipe_phv_out_data_213; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_214 = pipe3_io_pipe_phv_out_data_214; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_215 = pipe3_io_pipe_phv_out_data_215; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_216 = pipe3_io_pipe_phv_out_data_216; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_217 = pipe3_io_pipe_phv_out_data_217; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_218 = pipe3_io_pipe_phv_out_data_218; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_219 = pipe3_io_pipe_phv_out_data_219; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_220 = pipe3_io_pipe_phv_out_data_220; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_221 = pipe3_io_pipe_phv_out_data_221; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_222 = pipe3_io_pipe_phv_out_data_222; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_223 = pipe3_io_pipe_phv_out_data_223; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_224 = pipe3_io_pipe_phv_out_data_224; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_225 = pipe3_io_pipe_phv_out_data_225; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_226 = pipe3_io_pipe_phv_out_data_226; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_227 = pipe3_io_pipe_phv_out_data_227; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_228 = pipe3_io_pipe_phv_out_data_228; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_229 = pipe3_io_pipe_phv_out_data_229; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_230 = pipe3_io_pipe_phv_out_data_230; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_231 = pipe3_io_pipe_phv_out_data_231; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_232 = pipe3_io_pipe_phv_out_data_232; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_233 = pipe3_io_pipe_phv_out_data_233; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_234 = pipe3_io_pipe_phv_out_data_234; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_235 = pipe3_io_pipe_phv_out_data_235; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_236 = pipe3_io_pipe_phv_out_data_236; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_237 = pipe3_io_pipe_phv_out_data_237; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_238 = pipe3_io_pipe_phv_out_data_238; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_239 = pipe3_io_pipe_phv_out_data_239; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_240 = pipe3_io_pipe_phv_out_data_240; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_241 = pipe3_io_pipe_phv_out_data_241; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_242 = pipe3_io_pipe_phv_out_data_242; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_243 = pipe3_io_pipe_phv_out_data_243; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_244 = pipe3_io_pipe_phv_out_data_244; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_245 = pipe3_io_pipe_phv_out_data_245; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_246 = pipe3_io_pipe_phv_out_data_246; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_247 = pipe3_io_pipe_phv_out_data_247; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_248 = pipe3_io_pipe_phv_out_data_248; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_249 = pipe3_io_pipe_phv_out_data_249; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_250 = pipe3_io_pipe_phv_out_data_250; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_251 = pipe3_io_pipe_phv_out_data_251; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_252 = pipe3_io_pipe_phv_out_data_252; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_253 = pipe3_io_pipe_phv_out_data_253; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_254 = pipe3_io_pipe_phv_out_data_254; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_255 = pipe3_io_pipe_phv_out_data_255; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_256 = pipe3_io_pipe_phv_out_data_256; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_257 = pipe3_io_pipe_phv_out_data_257; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_258 = pipe3_io_pipe_phv_out_data_258; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_259 = pipe3_io_pipe_phv_out_data_259; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_260 = pipe3_io_pipe_phv_out_data_260; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_261 = pipe3_io_pipe_phv_out_data_261; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_262 = pipe3_io_pipe_phv_out_data_262; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_263 = pipe3_io_pipe_phv_out_data_263; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_264 = pipe3_io_pipe_phv_out_data_264; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_265 = pipe3_io_pipe_phv_out_data_265; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_266 = pipe3_io_pipe_phv_out_data_266; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_267 = pipe3_io_pipe_phv_out_data_267; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_268 = pipe3_io_pipe_phv_out_data_268; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_269 = pipe3_io_pipe_phv_out_data_269; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_270 = pipe3_io_pipe_phv_out_data_270; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_271 = pipe3_io_pipe_phv_out_data_271; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_272 = pipe3_io_pipe_phv_out_data_272; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_273 = pipe3_io_pipe_phv_out_data_273; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_274 = pipe3_io_pipe_phv_out_data_274; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_275 = pipe3_io_pipe_phv_out_data_275; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_276 = pipe3_io_pipe_phv_out_data_276; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_277 = pipe3_io_pipe_phv_out_data_277; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_278 = pipe3_io_pipe_phv_out_data_278; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_279 = pipe3_io_pipe_phv_out_data_279; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_280 = pipe3_io_pipe_phv_out_data_280; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_281 = pipe3_io_pipe_phv_out_data_281; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_282 = pipe3_io_pipe_phv_out_data_282; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_283 = pipe3_io_pipe_phv_out_data_283; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_284 = pipe3_io_pipe_phv_out_data_284; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_285 = pipe3_io_pipe_phv_out_data_285; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_286 = pipe3_io_pipe_phv_out_data_286; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_287 = pipe3_io_pipe_phv_out_data_287; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_288 = pipe3_io_pipe_phv_out_data_288; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_289 = pipe3_io_pipe_phv_out_data_289; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_290 = pipe3_io_pipe_phv_out_data_290; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_291 = pipe3_io_pipe_phv_out_data_291; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_292 = pipe3_io_pipe_phv_out_data_292; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_293 = pipe3_io_pipe_phv_out_data_293; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_294 = pipe3_io_pipe_phv_out_data_294; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_295 = pipe3_io_pipe_phv_out_data_295; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_296 = pipe3_io_pipe_phv_out_data_296; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_297 = pipe3_io_pipe_phv_out_data_297; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_298 = pipe3_io_pipe_phv_out_data_298; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_299 = pipe3_io_pipe_phv_out_data_299; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_300 = pipe3_io_pipe_phv_out_data_300; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_301 = pipe3_io_pipe_phv_out_data_301; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_302 = pipe3_io_pipe_phv_out_data_302; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_303 = pipe3_io_pipe_phv_out_data_303; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_304 = pipe3_io_pipe_phv_out_data_304; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_305 = pipe3_io_pipe_phv_out_data_305; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_306 = pipe3_io_pipe_phv_out_data_306; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_307 = pipe3_io_pipe_phv_out_data_307; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_308 = pipe3_io_pipe_phv_out_data_308; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_309 = pipe3_io_pipe_phv_out_data_309; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_310 = pipe3_io_pipe_phv_out_data_310; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_311 = pipe3_io_pipe_phv_out_data_311; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_312 = pipe3_io_pipe_phv_out_data_312; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_313 = pipe3_io_pipe_phv_out_data_313; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_314 = pipe3_io_pipe_phv_out_data_314; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_315 = pipe3_io_pipe_phv_out_data_315; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_316 = pipe3_io_pipe_phv_out_data_316; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_317 = pipe3_io_pipe_phv_out_data_317; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_318 = pipe3_io_pipe_phv_out_data_318; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_319 = pipe3_io_pipe_phv_out_data_319; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_320 = pipe3_io_pipe_phv_out_data_320; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_321 = pipe3_io_pipe_phv_out_data_321; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_322 = pipe3_io_pipe_phv_out_data_322; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_323 = pipe3_io_pipe_phv_out_data_323; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_324 = pipe3_io_pipe_phv_out_data_324; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_325 = pipe3_io_pipe_phv_out_data_325; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_326 = pipe3_io_pipe_phv_out_data_326; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_327 = pipe3_io_pipe_phv_out_data_327; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_328 = pipe3_io_pipe_phv_out_data_328; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_329 = pipe3_io_pipe_phv_out_data_329; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_330 = pipe3_io_pipe_phv_out_data_330; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_331 = pipe3_io_pipe_phv_out_data_331; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_332 = pipe3_io_pipe_phv_out_data_332; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_333 = pipe3_io_pipe_phv_out_data_333; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_334 = pipe3_io_pipe_phv_out_data_334; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_335 = pipe3_io_pipe_phv_out_data_335; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_336 = pipe3_io_pipe_phv_out_data_336; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_337 = pipe3_io_pipe_phv_out_data_337; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_338 = pipe3_io_pipe_phv_out_data_338; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_339 = pipe3_io_pipe_phv_out_data_339; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_340 = pipe3_io_pipe_phv_out_data_340; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_341 = pipe3_io_pipe_phv_out_data_341; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_342 = pipe3_io_pipe_phv_out_data_342; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_343 = pipe3_io_pipe_phv_out_data_343; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_344 = pipe3_io_pipe_phv_out_data_344; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_345 = pipe3_io_pipe_phv_out_data_345; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_346 = pipe3_io_pipe_phv_out_data_346; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_347 = pipe3_io_pipe_phv_out_data_347; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_348 = pipe3_io_pipe_phv_out_data_348; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_349 = pipe3_io_pipe_phv_out_data_349; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_350 = pipe3_io_pipe_phv_out_data_350; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_351 = pipe3_io_pipe_phv_out_data_351; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_352 = pipe3_io_pipe_phv_out_data_352; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_353 = pipe3_io_pipe_phv_out_data_353; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_354 = pipe3_io_pipe_phv_out_data_354; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_355 = pipe3_io_pipe_phv_out_data_355; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_356 = pipe3_io_pipe_phv_out_data_356; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_357 = pipe3_io_pipe_phv_out_data_357; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_358 = pipe3_io_pipe_phv_out_data_358; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_359 = pipe3_io_pipe_phv_out_data_359; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_360 = pipe3_io_pipe_phv_out_data_360; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_361 = pipe3_io_pipe_phv_out_data_361; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_362 = pipe3_io_pipe_phv_out_data_362; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_363 = pipe3_io_pipe_phv_out_data_363; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_364 = pipe3_io_pipe_phv_out_data_364; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_365 = pipe3_io_pipe_phv_out_data_365; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_366 = pipe3_io_pipe_phv_out_data_366; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_367 = pipe3_io_pipe_phv_out_data_367; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_368 = pipe3_io_pipe_phv_out_data_368; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_369 = pipe3_io_pipe_phv_out_data_369; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_370 = pipe3_io_pipe_phv_out_data_370; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_371 = pipe3_io_pipe_phv_out_data_371; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_372 = pipe3_io_pipe_phv_out_data_372; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_373 = pipe3_io_pipe_phv_out_data_373; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_374 = pipe3_io_pipe_phv_out_data_374; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_375 = pipe3_io_pipe_phv_out_data_375; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_376 = pipe3_io_pipe_phv_out_data_376; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_377 = pipe3_io_pipe_phv_out_data_377; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_378 = pipe3_io_pipe_phv_out_data_378; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_379 = pipe3_io_pipe_phv_out_data_379; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_380 = pipe3_io_pipe_phv_out_data_380; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_381 = pipe3_io_pipe_phv_out_data_381; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_382 = pipe3_io_pipe_phv_out_data_382; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_383 = pipe3_io_pipe_phv_out_data_383; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_384 = pipe3_io_pipe_phv_out_data_384; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_385 = pipe3_io_pipe_phv_out_data_385; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_386 = pipe3_io_pipe_phv_out_data_386; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_387 = pipe3_io_pipe_phv_out_data_387; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_388 = pipe3_io_pipe_phv_out_data_388; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_389 = pipe3_io_pipe_phv_out_data_389; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_390 = pipe3_io_pipe_phv_out_data_390; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_391 = pipe3_io_pipe_phv_out_data_391; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_392 = pipe3_io_pipe_phv_out_data_392; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_393 = pipe3_io_pipe_phv_out_data_393; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_394 = pipe3_io_pipe_phv_out_data_394; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_395 = pipe3_io_pipe_phv_out_data_395; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_396 = pipe3_io_pipe_phv_out_data_396; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_397 = pipe3_io_pipe_phv_out_data_397; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_398 = pipe3_io_pipe_phv_out_data_398; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_399 = pipe3_io_pipe_phv_out_data_399; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_400 = pipe3_io_pipe_phv_out_data_400; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_401 = pipe3_io_pipe_phv_out_data_401; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_402 = pipe3_io_pipe_phv_out_data_402; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_403 = pipe3_io_pipe_phv_out_data_403; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_404 = pipe3_io_pipe_phv_out_data_404; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_405 = pipe3_io_pipe_phv_out_data_405; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_406 = pipe3_io_pipe_phv_out_data_406; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_407 = pipe3_io_pipe_phv_out_data_407; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_408 = pipe3_io_pipe_phv_out_data_408; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_409 = pipe3_io_pipe_phv_out_data_409; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_410 = pipe3_io_pipe_phv_out_data_410; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_411 = pipe3_io_pipe_phv_out_data_411; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_412 = pipe3_io_pipe_phv_out_data_412; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_413 = pipe3_io_pipe_phv_out_data_413; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_414 = pipe3_io_pipe_phv_out_data_414; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_415 = pipe3_io_pipe_phv_out_data_415; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_416 = pipe3_io_pipe_phv_out_data_416; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_417 = pipe3_io_pipe_phv_out_data_417; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_418 = pipe3_io_pipe_phv_out_data_418; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_419 = pipe3_io_pipe_phv_out_data_419; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_420 = pipe3_io_pipe_phv_out_data_420; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_421 = pipe3_io_pipe_phv_out_data_421; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_422 = pipe3_io_pipe_phv_out_data_422; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_423 = pipe3_io_pipe_phv_out_data_423; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_424 = pipe3_io_pipe_phv_out_data_424; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_425 = pipe3_io_pipe_phv_out_data_425; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_426 = pipe3_io_pipe_phv_out_data_426; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_427 = pipe3_io_pipe_phv_out_data_427; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_428 = pipe3_io_pipe_phv_out_data_428; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_429 = pipe3_io_pipe_phv_out_data_429; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_430 = pipe3_io_pipe_phv_out_data_430; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_431 = pipe3_io_pipe_phv_out_data_431; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_432 = pipe3_io_pipe_phv_out_data_432; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_433 = pipe3_io_pipe_phv_out_data_433; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_434 = pipe3_io_pipe_phv_out_data_434; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_435 = pipe3_io_pipe_phv_out_data_435; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_436 = pipe3_io_pipe_phv_out_data_436; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_437 = pipe3_io_pipe_phv_out_data_437; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_438 = pipe3_io_pipe_phv_out_data_438; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_439 = pipe3_io_pipe_phv_out_data_439; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_440 = pipe3_io_pipe_phv_out_data_440; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_441 = pipe3_io_pipe_phv_out_data_441; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_442 = pipe3_io_pipe_phv_out_data_442; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_443 = pipe3_io_pipe_phv_out_data_443; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_444 = pipe3_io_pipe_phv_out_data_444; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_445 = pipe3_io_pipe_phv_out_data_445; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_446 = pipe3_io_pipe_phv_out_data_446; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_447 = pipe3_io_pipe_phv_out_data_447; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_448 = pipe3_io_pipe_phv_out_data_448; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_449 = pipe3_io_pipe_phv_out_data_449; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_450 = pipe3_io_pipe_phv_out_data_450; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_451 = pipe3_io_pipe_phv_out_data_451; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_452 = pipe3_io_pipe_phv_out_data_452; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_453 = pipe3_io_pipe_phv_out_data_453; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_454 = pipe3_io_pipe_phv_out_data_454; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_455 = pipe3_io_pipe_phv_out_data_455; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_456 = pipe3_io_pipe_phv_out_data_456; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_457 = pipe3_io_pipe_phv_out_data_457; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_458 = pipe3_io_pipe_phv_out_data_458; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_459 = pipe3_io_pipe_phv_out_data_459; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_460 = pipe3_io_pipe_phv_out_data_460; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_461 = pipe3_io_pipe_phv_out_data_461; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_462 = pipe3_io_pipe_phv_out_data_462; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_463 = pipe3_io_pipe_phv_out_data_463; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_464 = pipe3_io_pipe_phv_out_data_464; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_465 = pipe3_io_pipe_phv_out_data_465; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_466 = pipe3_io_pipe_phv_out_data_466; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_467 = pipe3_io_pipe_phv_out_data_467; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_468 = pipe3_io_pipe_phv_out_data_468; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_469 = pipe3_io_pipe_phv_out_data_469; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_470 = pipe3_io_pipe_phv_out_data_470; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_471 = pipe3_io_pipe_phv_out_data_471; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_472 = pipe3_io_pipe_phv_out_data_472; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_473 = pipe3_io_pipe_phv_out_data_473; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_474 = pipe3_io_pipe_phv_out_data_474; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_475 = pipe3_io_pipe_phv_out_data_475; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_476 = pipe3_io_pipe_phv_out_data_476; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_477 = pipe3_io_pipe_phv_out_data_477; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_478 = pipe3_io_pipe_phv_out_data_478; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_479 = pipe3_io_pipe_phv_out_data_479; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_480 = pipe3_io_pipe_phv_out_data_480; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_481 = pipe3_io_pipe_phv_out_data_481; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_482 = pipe3_io_pipe_phv_out_data_482; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_483 = pipe3_io_pipe_phv_out_data_483; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_484 = pipe3_io_pipe_phv_out_data_484; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_485 = pipe3_io_pipe_phv_out_data_485; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_486 = pipe3_io_pipe_phv_out_data_486; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_487 = pipe3_io_pipe_phv_out_data_487; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_488 = pipe3_io_pipe_phv_out_data_488; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_489 = pipe3_io_pipe_phv_out_data_489; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_490 = pipe3_io_pipe_phv_out_data_490; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_491 = pipe3_io_pipe_phv_out_data_491; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_492 = pipe3_io_pipe_phv_out_data_492; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_493 = pipe3_io_pipe_phv_out_data_493; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_494 = pipe3_io_pipe_phv_out_data_494; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_495 = pipe3_io_pipe_phv_out_data_495; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_496 = pipe3_io_pipe_phv_out_data_496; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_497 = pipe3_io_pipe_phv_out_data_497; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_498 = pipe3_io_pipe_phv_out_data_498; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_499 = pipe3_io_pipe_phv_out_data_499; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_500 = pipe3_io_pipe_phv_out_data_500; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_501 = pipe3_io_pipe_phv_out_data_501; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_502 = pipe3_io_pipe_phv_out_data_502; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_503 = pipe3_io_pipe_phv_out_data_503; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_504 = pipe3_io_pipe_phv_out_data_504; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_505 = pipe3_io_pipe_phv_out_data_505; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_506 = pipe3_io_pipe_phv_out_data_506; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_507 = pipe3_io_pipe_phv_out_data_507; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_508 = pipe3_io_pipe_phv_out_data_508; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_509 = pipe3_io_pipe_phv_out_data_509; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_510 = pipe3_io_pipe_phv_out_data_510; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_data_511 = pipe3_io_pipe_phv_out_data_511; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_0 = pipe3_io_pipe_phv_out_header_0; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_1 = pipe3_io_pipe_phv_out_header_1; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_2 = pipe3_io_pipe_phv_out_header_2; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_3 = pipe3_io_pipe_phv_out_header_3; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_4 = pipe3_io_pipe_phv_out_header_4; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_5 = pipe3_io_pipe_phv_out_header_5; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_6 = pipe3_io_pipe_phv_out_header_6; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_7 = pipe3_io_pipe_phv_out_header_7; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_8 = pipe3_io_pipe_phv_out_header_8; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_9 = pipe3_io_pipe_phv_out_header_9; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_10 = pipe3_io_pipe_phv_out_header_10; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_11 = pipe3_io_pipe_phv_out_header_11; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_12 = pipe3_io_pipe_phv_out_header_12; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_13 = pipe3_io_pipe_phv_out_header_13; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_14 = pipe3_io_pipe_phv_out_header_14; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_header_15 = pipe3_io_pipe_phv_out_header_15; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_parse_current_state = pipe3_io_pipe_phv_out_parse_current_state; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_parse_current_offset = pipe3_io_pipe_phv_out_parse_current_offset; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_parse_transition_field = pipe3_io_pipe_phv_out_parse_transition_field; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_next_processor_id = pipe3_io_pipe_phv_out_next_processor_id; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_next_config_id = pipe3_io_pipe_phv_out_next_config_id; // @[executor.scala 511:27]
  assign pipe4_io_pipe_phv_in_is_valid_processor = pipe3_io_pipe_phv_out_is_valid_processor; // @[executor.scala 511:27]
  assign pipe4_io_vliw_in_0 = pipe3_io_vliw_out_0; // @[executor.scala 512:27]
  assign pipe4_io_vliw_in_1 = pipe3_io_vliw_out_1; // @[executor.scala 512:27]
  assign pipe4_io_vliw_in_2 = pipe3_io_vliw_out_2; // @[executor.scala 512:27]
  assign pipe4_io_vliw_in_3 = pipe3_io_vliw_out_3; // @[executor.scala 512:27]
  assign pipe4_io_field_in_0 = pipe3_io_field_out_0; // @[executor.scala 513:27]
  assign pipe4_io_field_in_1 = pipe3_io_field_out_1; // @[executor.scala 513:27]
  assign pipe4_io_field_in_2 = pipe3_io_field_out_2; // @[executor.scala 513:27]
  assign pipe4_io_field_in_3 = pipe3_io_field_out_3; // @[executor.scala 513:27]
  assign pipe4_io_mask_in_0 = pipe3_io_mask_out_0; // @[executor.scala 514:27]
  assign pipe4_io_mask_in_1 = pipe3_io_mask_out_1; // @[executor.scala 514:27]
  assign pipe4_io_mask_in_2 = pipe3_io_mask_out_2; // @[executor.scala 514:27]
  assign pipe4_io_mask_in_3 = pipe3_io_mask_out_3; // @[executor.scala 514:27]
  assign pipe4_io_bias_in_0 = pipe3_io_bias_out_0; // @[executor.scala 515:27]
  assign pipe4_io_bias_in_1 = pipe3_io_bias_out_1; // @[executor.scala 515:27]
  assign pipe4_io_bias_in_2 = pipe3_io_bias_out_2; // @[executor.scala 515:27]
  assign pipe4_io_bias_in_3 = pipe3_io_bias_out_3; // @[executor.scala 515:27]
  assign pipe5_clock = clock;
  assign pipe5_io_pipe_phv_in_data_0 = pipe4_io_pipe_phv_out_data_0; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_1 = pipe4_io_pipe_phv_out_data_1; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_2 = pipe4_io_pipe_phv_out_data_2; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_3 = pipe4_io_pipe_phv_out_data_3; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_4 = pipe4_io_pipe_phv_out_data_4; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_5 = pipe4_io_pipe_phv_out_data_5; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_6 = pipe4_io_pipe_phv_out_data_6; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_7 = pipe4_io_pipe_phv_out_data_7; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_8 = pipe4_io_pipe_phv_out_data_8; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_9 = pipe4_io_pipe_phv_out_data_9; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_10 = pipe4_io_pipe_phv_out_data_10; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_11 = pipe4_io_pipe_phv_out_data_11; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_12 = pipe4_io_pipe_phv_out_data_12; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_13 = pipe4_io_pipe_phv_out_data_13; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_14 = pipe4_io_pipe_phv_out_data_14; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_15 = pipe4_io_pipe_phv_out_data_15; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_16 = pipe4_io_pipe_phv_out_data_16; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_17 = pipe4_io_pipe_phv_out_data_17; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_18 = pipe4_io_pipe_phv_out_data_18; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_19 = pipe4_io_pipe_phv_out_data_19; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_20 = pipe4_io_pipe_phv_out_data_20; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_21 = pipe4_io_pipe_phv_out_data_21; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_22 = pipe4_io_pipe_phv_out_data_22; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_23 = pipe4_io_pipe_phv_out_data_23; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_24 = pipe4_io_pipe_phv_out_data_24; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_25 = pipe4_io_pipe_phv_out_data_25; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_26 = pipe4_io_pipe_phv_out_data_26; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_27 = pipe4_io_pipe_phv_out_data_27; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_28 = pipe4_io_pipe_phv_out_data_28; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_29 = pipe4_io_pipe_phv_out_data_29; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_30 = pipe4_io_pipe_phv_out_data_30; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_31 = pipe4_io_pipe_phv_out_data_31; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_32 = pipe4_io_pipe_phv_out_data_32; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_33 = pipe4_io_pipe_phv_out_data_33; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_34 = pipe4_io_pipe_phv_out_data_34; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_35 = pipe4_io_pipe_phv_out_data_35; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_36 = pipe4_io_pipe_phv_out_data_36; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_37 = pipe4_io_pipe_phv_out_data_37; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_38 = pipe4_io_pipe_phv_out_data_38; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_39 = pipe4_io_pipe_phv_out_data_39; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_40 = pipe4_io_pipe_phv_out_data_40; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_41 = pipe4_io_pipe_phv_out_data_41; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_42 = pipe4_io_pipe_phv_out_data_42; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_43 = pipe4_io_pipe_phv_out_data_43; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_44 = pipe4_io_pipe_phv_out_data_44; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_45 = pipe4_io_pipe_phv_out_data_45; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_46 = pipe4_io_pipe_phv_out_data_46; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_47 = pipe4_io_pipe_phv_out_data_47; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_48 = pipe4_io_pipe_phv_out_data_48; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_49 = pipe4_io_pipe_phv_out_data_49; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_50 = pipe4_io_pipe_phv_out_data_50; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_51 = pipe4_io_pipe_phv_out_data_51; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_52 = pipe4_io_pipe_phv_out_data_52; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_53 = pipe4_io_pipe_phv_out_data_53; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_54 = pipe4_io_pipe_phv_out_data_54; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_55 = pipe4_io_pipe_phv_out_data_55; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_56 = pipe4_io_pipe_phv_out_data_56; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_57 = pipe4_io_pipe_phv_out_data_57; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_58 = pipe4_io_pipe_phv_out_data_58; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_59 = pipe4_io_pipe_phv_out_data_59; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_60 = pipe4_io_pipe_phv_out_data_60; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_61 = pipe4_io_pipe_phv_out_data_61; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_62 = pipe4_io_pipe_phv_out_data_62; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_63 = pipe4_io_pipe_phv_out_data_63; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_64 = pipe4_io_pipe_phv_out_data_64; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_65 = pipe4_io_pipe_phv_out_data_65; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_66 = pipe4_io_pipe_phv_out_data_66; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_67 = pipe4_io_pipe_phv_out_data_67; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_68 = pipe4_io_pipe_phv_out_data_68; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_69 = pipe4_io_pipe_phv_out_data_69; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_70 = pipe4_io_pipe_phv_out_data_70; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_71 = pipe4_io_pipe_phv_out_data_71; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_72 = pipe4_io_pipe_phv_out_data_72; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_73 = pipe4_io_pipe_phv_out_data_73; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_74 = pipe4_io_pipe_phv_out_data_74; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_75 = pipe4_io_pipe_phv_out_data_75; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_76 = pipe4_io_pipe_phv_out_data_76; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_77 = pipe4_io_pipe_phv_out_data_77; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_78 = pipe4_io_pipe_phv_out_data_78; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_79 = pipe4_io_pipe_phv_out_data_79; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_80 = pipe4_io_pipe_phv_out_data_80; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_81 = pipe4_io_pipe_phv_out_data_81; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_82 = pipe4_io_pipe_phv_out_data_82; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_83 = pipe4_io_pipe_phv_out_data_83; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_84 = pipe4_io_pipe_phv_out_data_84; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_85 = pipe4_io_pipe_phv_out_data_85; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_86 = pipe4_io_pipe_phv_out_data_86; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_87 = pipe4_io_pipe_phv_out_data_87; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_88 = pipe4_io_pipe_phv_out_data_88; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_89 = pipe4_io_pipe_phv_out_data_89; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_90 = pipe4_io_pipe_phv_out_data_90; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_91 = pipe4_io_pipe_phv_out_data_91; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_92 = pipe4_io_pipe_phv_out_data_92; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_93 = pipe4_io_pipe_phv_out_data_93; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_94 = pipe4_io_pipe_phv_out_data_94; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_95 = pipe4_io_pipe_phv_out_data_95; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_96 = pipe4_io_pipe_phv_out_data_96; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_97 = pipe4_io_pipe_phv_out_data_97; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_98 = pipe4_io_pipe_phv_out_data_98; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_99 = pipe4_io_pipe_phv_out_data_99; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_100 = pipe4_io_pipe_phv_out_data_100; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_101 = pipe4_io_pipe_phv_out_data_101; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_102 = pipe4_io_pipe_phv_out_data_102; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_103 = pipe4_io_pipe_phv_out_data_103; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_104 = pipe4_io_pipe_phv_out_data_104; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_105 = pipe4_io_pipe_phv_out_data_105; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_106 = pipe4_io_pipe_phv_out_data_106; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_107 = pipe4_io_pipe_phv_out_data_107; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_108 = pipe4_io_pipe_phv_out_data_108; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_109 = pipe4_io_pipe_phv_out_data_109; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_110 = pipe4_io_pipe_phv_out_data_110; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_111 = pipe4_io_pipe_phv_out_data_111; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_112 = pipe4_io_pipe_phv_out_data_112; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_113 = pipe4_io_pipe_phv_out_data_113; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_114 = pipe4_io_pipe_phv_out_data_114; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_115 = pipe4_io_pipe_phv_out_data_115; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_116 = pipe4_io_pipe_phv_out_data_116; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_117 = pipe4_io_pipe_phv_out_data_117; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_118 = pipe4_io_pipe_phv_out_data_118; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_119 = pipe4_io_pipe_phv_out_data_119; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_120 = pipe4_io_pipe_phv_out_data_120; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_121 = pipe4_io_pipe_phv_out_data_121; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_122 = pipe4_io_pipe_phv_out_data_122; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_123 = pipe4_io_pipe_phv_out_data_123; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_124 = pipe4_io_pipe_phv_out_data_124; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_125 = pipe4_io_pipe_phv_out_data_125; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_126 = pipe4_io_pipe_phv_out_data_126; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_127 = pipe4_io_pipe_phv_out_data_127; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_128 = pipe4_io_pipe_phv_out_data_128; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_129 = pipe4_io_pipe_phv_out_data_129; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_130 = pipe4_io_pipe_phv_out_data_130; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_131 = pipe4_io_pipe_phv_out_data_131; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_132 = pipe4_io_pipe_phv_out_data_132; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_133 = pipe4_io_pipe_phv_out_data_133; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_134 = pipe4_io_pipe_phv_out_data_134; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_135 = pipe4_io_pipe_phv_out_data_135; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_136 = pipe4_io_pipe_phv_out_data_136; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_137 = pipe4_io_pipe_phv_out_data_137; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_138 = pipe4_io_pipe_phv_out_data_138; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_139 = pipe4_io_pipe_phv_out_data_139; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_140 = pipe4_io_pipe_phv_out_data_140; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_141 = pipe4_io_pipe_phv_out_data_141; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_142 = pipe4_io_pipe_phv_out_data_142; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_143 = pipe4_io_pipe_phv_out_data_143; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_144 = pipe4_io_pipe_phv_out_data_144; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_145 = pipe4_io_pipe_phv_out_data_145; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_146 = pipe4_io_pipe_phv_out_data_146; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_147 = pipe4_io_pipe_phv_out_data_147; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_148 = pipe4_io_pipe_phv_out_data_148; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_149 = pipe4_io_pipe_phv_out_data_149; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_150 = pipe4_io_pipe_phv_out_data_150; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_151 = pipe4_io_pipe_phv_out_data_151; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_152 = pipe4_io_pipe_phv_out_data_152; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_153 = pipe4_io_pipe_phv_out_data_153; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_154 = pipe4_io_pipe_phv_out_data_154; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_155 = pipe4_io_pipe_phv_out_data_155; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_156 = pipe4_io_pipe_phv_out_data_156; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_157 = pipe4_io_pipe_phv_out_data_157; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_158 = pipe4_io_pipe_phv_out_data_158; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_159 = pipe4_io_pipe_phv_out_data_159; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_160 = pipe4_io_pipe_phv_out_data_160; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_161 = pipe4_io_pipe_phv_out_data_161; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_162 = pipe4_io_pipe_phv_out_data_162; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_163 = pipe4_io_pipe_phv_out_data_163; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_164 = pipe4_io_pipe_phv_out_data_164; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_165 = pipe4_io_pipe_phv_out_data_165; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_166 = pipe4_io_pipe_phv_out_data_166; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_167 = pipe4_io_pipe_phv_out_data_167; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_168 = pipe4_io_pipe_phv_out_data_168; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_169 = pipe4_io_pipe_phv_out_data_169; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_170 = pipe4_io_pipe_phv_out_data_170; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_171 = pipe4_io_pipe_phv_out_data_171; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_172 = pipe4_io_pipe_phv_out_data_172; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_173 = pipe4_io_pipe_phv_out_data_173; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_174 = pipe4_io_pipe_phv_out_data_174; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_175 = pipe4_io_pipe_phv_out_data_175; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_176 = pipe4_io_pipe_phv_out_data_176; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_177 = pipe4_io_pipe_phv_out_data_177; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_178 = pipe4_io_pipe_phv_out_data_178; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_179 = pipe4_io_pipe_phv_out_data_179; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_180 = pipe4_io_pipe_phv_out_data_180; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_181 = pipe4_io_pipe_phv_out_data_181; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_182 = pipe4_io_pipe_phv_out_data_182; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_183 = pipe4_io_pipe_phv_out_data_183; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_184 = pipe4_io_pipe_phv_out_data_184; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_185 = pipe4_io_pipe_phv_out_data_185; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_186 = pipe4_io_pipe_phv_out_data_186; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_187 = pipe4_io_pipe_phv_out_data_187; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_188 = pipe4_io_pipe_phv_out_data_188; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_189 = pipe4_io_pipe_phv_out_data_189; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_190 = pipe4_io_pipe_phv_out_data_190; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_191 = pipe4_io_pipe_phv_out_data_191; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_192 = pipe4_io_pipe_phv_out_data_192; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_193 = pipe4_io_pipe_phv_out_data_193; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_194 = pipe4_io_pipe_phv_out_data_194; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_195 = pipe4_io_pipe_phv_out_data_195; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_196 = pipe4_io_pipe_phv_out_data_196; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_197 = pipe4_io_pipe_phv_out_data_197; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_198 = pipe4_io_pipe_phv_out_data_198; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_199 = pipe4_io_pipe_phv_out_data_199; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_200 = pipe4_io_pipe_phv_out_data_200; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_201 = pipe4_io_pipe_phv_out_data_201; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_202 = pipe4_io_pipe_phv_out_data_202; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_203 = pipe4_io_pipe_phv_out_data_203; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_204 = pipe4_io_pipe_phv_out_data_204; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_205 = pipe4_io_pipe_phv_out_data_205; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_206 = pipe4_io_pipe_phv_out_data_206; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_207 = pipe4_io_pipe_phv_out_data_207; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_208 = pipe4_io_pipe_phv_out_data_208; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_209 = pipe4_io_pipe_phv_out_data_209; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_210 = pipe4_io_pipe_phv_out_data_210; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_211 = pipe4_io_pipe_phv_out_data_211; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_212 = pipe4_io_pipe_phv_out_data_212; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_213 = pipe4_io_pipe_phv_out_data_213; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_214 = pipe4_io_pipe_phv_out_data_214; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_215 = pipe4_io_pipe_phv_out_data_215; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_216 = pipe4_io_pipe_phv_out_data_216; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_217 = pipe4_io_pipe_phv_out_data_217; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_218 = pipe4_io_pipe_phv_out_data_218; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_219 = pipe4_io_pipe_phv_out_data_219; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_220 = pipe4_io_pipe_phv_out_data_220; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_221 = pipe4_io_pipe_phv_out_data_221; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_222 = pipe4_io_pipe_phv_out_data_222; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_223 = pipe4_io_pipe_phv_out_data_223; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_224 = pipe4_io_pipe_phv_out_data_224; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_225 = pipe4_io_pipe_phv_out_data_225; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_226 = pipe4_io_pipe_phv_out_data_226; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_227 = pipe4_io_pipe_phv_out_data_227; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_228 = pipe4_io_pipe_phv_out_data_228; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_229 = pipe4_io_pipe_phv_out_data_229; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_230 = pipe4_io_pipe_phv_out_data_230; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_231 = pipe4_io_pipe_phv_out_data_231; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_232 = pipe4_io_pipe_phv_out_data_232; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_233 = pipe4_io_pipe_phv_out_data_233; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_234 = pipe4_io_pipe_phv_out_data_234; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_235 = pipe4_io_pipe_phv_out_data_235; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_236 = pipe4_io_pipe_phv_out_data_236; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_237 = pipe4_io_pipe_phv_out_data_237; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_238 = pipe4_io_pipe_phv_out_data_238; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_239 = pipe4_io_pipe_phv_out_data_239; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_240 = pipe4_io_pipe_phv_out_data_240; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_241 = pipe4_io_pipe_phv_out_data_241; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_242 = pipe4_io_pipe_phv_out_data_242; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_243 = pipe4_io_pipe_phv_out_data_243; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_244 = pipe4_io_pipe_phv_out_data_244; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_245 = pipe4_io_pipe_phv_out_data_245; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_246 = pipe4_io_pipe_phv_out_data_246; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_247 = pipe4_io_pipe_phv_out_data_247; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_248 = pipe4_io_pipe_phv_out_data_248; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_249 = pipe4_io_pipe_phv_out_data_249; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_250 = pipe4_io_pipe_phv_out_data_250; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_251 = pipe4_io_pipe_phv_out_data_251; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_252 = pipe4_io_pipe_phv_out_data_252; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_253 = pipe4_io_pipe_phv_out_data_253; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_254 = pipe4_io_pipe_phv_out_data_254; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_255 = pipe4_io_pipe_phv_out_data_255; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_256 = pipe4_io_pipe_phv_out_data_256; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_257 = pipe4_io_pipe_phv_out_data_257; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_258 = pipe4_io_pipe_phv_out_data_258; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_259 = pipe4_io_pipe_phv_out_data_259; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_260 = pipe4_io_pipe_phv_out_data_260; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_261 = pipe4_io_pipe_phv_out_data_261; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_262 = pipe4_io_pipe_phv_out_data_262; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_263 = pipe4_io_pipe_phv_out_data_263; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_264 = pipe4_io_pipe_phv_out_data_264; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_265 = pipe4_io_pipe_phv_out_data_265; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_266 = pipe4_io_pipe_phv_out_data_266; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_267 = pipe4_io_pipe_phv_out_data_267; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_268 = pipe4_io_pipe_phv_out_data_268; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_269 = pipe4_io_pipe_phv_out_data_269; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_270 = pipe4_io_pipe_phv_out_data_270; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_271 = pipe4_io_pipe_phv_out_data_271; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_272 = pipe4_io_pipe_phv_out_data_272; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_273 = pipe4_io_pipe_phv_out_data_273; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_274 = pipe4_io_pipe_phv_out_data_274; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_275 = pipe4_io_pipe_phv_out_data_275; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_276 = pipe4_io_pipe_phv_out_data_276; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_277 = pipe4_io_pipe_phv_out_data_277; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_278 = pipe4_io_pipe_phv_out_data_278; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_279 = pipe4_io_pipe_phv_out_data_279; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_280 = pipe4_io_pipe_phv_out_data_280; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_281 = pipe4_io_pipe_phv_out_data_281; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_282 = pipe4_io_pipe_phv_out_data_282; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_283 = pipe4_io_pipe_phv_out_data_283; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_284 = pipe4_io_pipe_phv_out_data_284; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_285 = pipe4_io_pipe_phv_out_data_285; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_286 = pipe4_io_pipe_phv_out_data_286; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_287 = pipe4_io_pipe_phv_out_data_287; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_288 = pipe4_io_pipe_phv_out_data_288; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_289 = pipe4_io_pipe_phv_out_data_289; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_290 = pipe4_io_pipe_phv_out_data_290; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_291 = pipe4_io_pipe_phv_out_data_291; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_292 = pipe4_io_pipe_phv_out_data_292; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_293 = pipe4_io_pipe_phv_out_data_293; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_294 = pipe4_io_pipe_phv_out_data_294; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_295 = pipe4_io_pipe_phv_out_data_295; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_296 = pipe4_io_pipe_phv_out_data_296; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_297 = pipe4_io_pipe_phv_out_data_297; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_298 = pipe4_io_pipe_phv_out_data_298; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_299 = pipe4_io_pipe_phv_out_data_299; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_300 = pipe4_io_pipe_phv_out_data_300; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_301 = pipe4_io_pipe_phv_out_data_301; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_302 = pipe4_io_pipe_phv_out_data_302; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_303 = pipe4_io_pipe_phv_out_data_303; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_304 = pipe4_io_pipe_phv_out_data_304; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_305 = pipe4_io_pipe_phv_out_data_305; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_306 = pipe4_io_pipe_phv_out_data_306; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_307 = pipe4_io_pipe_phv_out_data_307; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_308 = pipe4_io_pipe_phv_out_data_308; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_309 = pipe4_io_pipe_phv_out_data_309; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_310 = pipe4_io_pipe_phv_out_data_310; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_311 = pipe4_io_pipe_phv_out_data_311; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_312 = pipe4_io_pipe_phv_out_data_312; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_313 = pipe4_io_pipe_phv_out_data_313; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_314 = pipe4_io_pipe_phv_out_data_314; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_315 = pipe4_io_pipe_phv_out_data_315; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_316 = pipe4_io_pipe_phv_out_data_316; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_317 = pipe4_io_pipe_phv_out_data_317; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_318 = pipe4_io_pipe_phv_out_data_318; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_319 = pipe4_io_pipe_phv_out_data_319; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_320 = pipe4_io_pipe_phv_out_data_320; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_321 = pipe4_io_pipe_phv_out_data_321; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_322 = pipe4_io_pipe_phv_out_data_322; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_323 = pipe4_io_pipe_phv_out_data_323; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_324 = pipe4_io_pipe_phv_out_data_324; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_325 = pipe4_io_pipe_phv_out_data_325; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_326 = pipe4_io_pipe_phv_out_data_326; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_327 = pipe4_io_pipe_phv_out_data_327; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_328 = pipe4_io_pipe_phv_out_data_328; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_329 = pipe4_io_pipe_phv_out_data_329; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_330 = pipe4_io_pipe_phv_out_data_330; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_331 = pipe4_io_pipe_phv_out_data_331; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_332 = pipe4_io_pipe_phv_out_data_332; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_333 = pipe4_io_pipe_phv_out_data_333; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_334 = pipe4_io_pipe_phv_out_data_334; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_335 = pipe4_io_pipe_phv_out_data_335; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_336 = pipe4_io_pipe_phv_out_data_336; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_337 = pipe4_io_pipe_phv_out_data_337; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_338 = pipe4_io_pipe_phv_out_data_338; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_339 = pipe4_io_pipe_phv_out_data_339; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_340 = pipe4_io_pipe_phv_out_data_340; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_341 = pipe4_io_pipe_phv_out_data_341; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_342 = pipe4_io_pipe_phv_out_data_342; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_343 = pipe4_io_pipe_phv_out_data_343; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_344 = pipe4_io_pipe_phv_out_data_344; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_345 = pipe4_io_pipe_phv_out_data_345; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_346 = pipe4_io_pipe_phv_out_data_346; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_347 = pipe4_io_pipe_phv_out_data_347; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_348 = pipe4_io_pipe_phv_out_data_348; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_349 = pipe4_io_pipe_phv_out_data_349; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_350 = pipe4_io_pipe_phv_out_data_350; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_351 = pipe4_io_pipe_phv_out_data_351; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_352 = pipe4_io_pipe_phv_out_data_352; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_353 = pipe4_io_pipe_phv_out_data_353; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_354 = pipe4_io_pipe_phv_out_data_354; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_355 = pipe4_io_pipe_phv_out_data_355; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_356 = pipe4_io_pipe_phv_out_data_356; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_357 = pipe4_io_pipe_phv_out_data_357; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_358 = pipe4_io_pipe_phv_out_data_358; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_359 = pipe4_io_pipe_phv_out_data_359; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_360 = pipe4_io_pipe_phv_out_data_360; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_361 = pipe4_io_pipe_phv_out_data_361; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_362 = pipe4_io_pipe_phv_out_data_362; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_363 = pipe4_io_pipe_phv_out_data_363; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_364 = pipe4_io_pipe_phv_out_data_364; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_365 = pipe4_io_pipe_phv_out_data_365; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_366 = pipe4_io_pipe_phv_out_data_366; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_367 = pipe4_io_pipe_phv_out_data_367; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_368 = pipe4_io_pipe_phv_out_data_368; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_369 = pipe4_io_pipe_phv_out_data_369; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_370 = pipe4_io_pipe_phv_out_data_370; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_371 = pipe4_io_pipe_phv_out_data_371; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_372 = pipe4_io_pipe_phv_out_data_372; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_373 = pipe4_io_pipe_phv_out_data_373; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_374 = pipe4_io_pipe_phv_out_data_374; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_375 = pipe4_io_pipe_phv_out_data_375; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_376 = pipe4_io_pipe_phv_out_data_376; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_377 = pipe4_io_pipe_phv_out_data_377; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_378 = pipe4_io_pipe_phv_out_data_378; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_379 = pipe4_io_pipe_phv_out_data_379; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_380 = pipe4_io_pipe_phv_out_data_380; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_381 = pipe4_io_pipe_phv_out_data_381; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_382 = pipe4_io_pipe_phv_out_data_382; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_383 = pipe4_io_pipe_phv_out_data_383; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_384 = pipe4_io_pipe_phv_out_data_384; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_385 = pipe4_io_pipe_phv_out_data_385; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_386 = pipe4_io_pipe_phv_out_data_386; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_387 = pipe4_io_pipe_phv_out_data_387; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_388 = pipe4_io_pipe_phv_out_data_388; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_389 = pipe4_io_pipe_phv_out_data_389; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_390 = pipe4_io_pipe_phv_out_data_390; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_391 = pipe4_io_pipe_phv_out_data_391; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_392 = pipe4_io_pipe_phv_out_data_392; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_393 = pipe4_io_pipe_phv_out_data_393; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_394 = pipe4_io_pipe_phv_out_data_394; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_395 = pipe4_io_pipe_phv_out_data_395; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_396 = pipe4_io_pipe_phv_out_data_396; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_397 = pipe4_io_pipe_phv_out_data_397; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_398 = pipe4_io_pipe_phv_out_data_398; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_399 = pipe4_io_pipe_phv_out_data_399; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_400 = pipe4_io_pipe_phv_out_data_400; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_401 = pipe4_io_pipe_phv_out_data_401; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_402 = pipe4_io_pipe_phv_out_data_402; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_403 = pipe4_io_pipe_phv_out_data_403; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_404 = pipe4_io_pipe_phv_out_data_404; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_405 = pipe4_io_pipe_phv_out_data_405; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_406 = pipe4_io_pipe_phv_out_data_406; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_407 = pipe4_io_pipe_phv_out_data_407; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_408 = pipe4_io_pipe_phv_out_data_408; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_409 = pipe4_io_pipe_phv_out_data_409; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_410 = pipe4_io_pipe_phv_out_data_410; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_411 = pipe4_io_pipe_phv_out_data_411; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_412 = pipe4_io_pipe_phv_out_data_412; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_413 = pipe4_io_pipe_phv_out_data_413; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_414 = pipe4_io_pipe_phv_out_data_414; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_415 = pipe4_io_pipe_phv_out_data_415; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_416 = pipe4_io_pipe_phv_out_data_416; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_417 = pipe4_io_pipe_phv_out_data_417; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_418 = pipe4_io_pipe_phv_out_data_418; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_419 = pipe4_io_pipe_phv_out_data_419; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_420 = pipe4_io_pipe_phv_out_data_420; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_421 = pipe4_io_pipe_phv_out_data_421; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_422 = pipe4_io_pipe_phv_out_data_422; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_423 = pipe4_io_pipe_phv_out_data_423; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_424 = pipe4_io_pipe_phv_out_data_424; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_425 = pipe4_io_pipe_phv_out_data_425; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_426 = pipe4_io_pipe_phv_out_data_426; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_427 = pipe4_io_pipe_phv_out_data_427; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_428 = pipe4_io_pipe_phv_out_data_428; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_429 = pipe4_io_pipe_phv_out_data_429; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_430 = pipe4_io_pipe_phv_out_data_430; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_431 = pipe4_io_pipe_phv_out_data_431; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_432 = pipe4_io_pipe_phv_out_data_432; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_433 = pipe4_io_pipe_phv_out_data_433; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_434 = pipe4_io_pipe_phv_out_data_434; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_435 = pipe4_io_pipe_phv_out_data_435; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_436 = pipe4_io_pipe_phv_out_data_436; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_437 = pipe4_io_pipe_phv_out_data_437; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_438 = pipe4_io_pipe_phv_out_data_438; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_439 = pipe4_io_pipe_phv_out_data_439; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_440 = pipe4_io_pipe_phv_out_data_440; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_441 = pipe4_io_pipe_phv_out_data_441; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_442 = pipe4_io_pipe_phv_out_data_442; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_443 = pipe4_io_pipe_phv_out_data_443; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_444 = pipe4_io_pipe_phv_out_data_444; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_445 = pipe4_io_pipe_phv_out_data_445; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_446 = pipe4_io_pipe_phv_out_data_446; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_447 = pipe4_io_pipe_phv_out_data_447; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_448 = pipe4_io_pipe_phv_out_data_448; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_449 = pipe4_io_pipe_phv_out_data_449; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_450 = pipe4_io_pipe_phv_out_data_450; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_451 = pipe4_io_pipe_phv_out_data_451; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_452 = pipe4_io_pipe_phv_out_data_452; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_453 = pipe4_io_pipe_phv_out_data_453; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_454 = pipe4_io_pipe_phv_out_data_454; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_455 = pipe4_io_pipe_phv_out_data_455; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_456 = pipe4_io_pipe_phv_out_data_456; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_457 = pipe4_io_pipe_phv_out_data_457; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_458 = pipe4_io_pipe_phv_out_data_458; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_459 = pipe4_io_pipe_phv_out_data_459; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_460 = pipe4_io_pipe_phv_out_data_460; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_461 = pipe4_io_pipe_phv_out_data_461; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_462 = pipe4_io_pipe_phv_out_data_462; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_463 = pipe4_io_pipe_phv_out_data_463; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_464 = pipe4_io_pipe_phv_out_data_464; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_465 = pipe4_io_pipe_phv_out_data_465; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_466 = pipe4_io_pipe_phv_out_data_466; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_467 = pipe4_io_pipe_phv_out_data_467; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_468 = pipe4_io_pipe_phv_out_data_468; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_469 = pipe4_io_pipe_phv_out_data_469; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_470 = pipe4_io_pipe_phv_out_data_470; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_471 = pipe4_io_pipe_phv_out_data_471; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_472 = pipe4_io_pipe_phv_out_data_472; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_473 = pipe4_io_pipe_phv_out_data_473; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_474 = pipe4_io_pipe_phv_out_data_474; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_475 = pipe4_io_pipe_phv_out_data_475; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_476 = pipe4_io_pipe_phv_out_data_476; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_477 = pipe4_io_pipe_phv_out_data_477; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_478 = pipe4_io_pipe_phv_out_data_478; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_479 = pipe4_io_pipe_phv_out_data_479; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_480 = pipe4_io_pipe_phv_out_data_480; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_481 = pipe4_io_pipe_phv_out_data_481; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_482 = pipe4_io_pipe_phv_out_data_482; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_483 = pipe4_io_pipe_phv_out_data_483; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_484 = pipe4_io_pipe_phv_out_data_484; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_485 = pipe4_io_pipe_phv_out_data_485; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_486 = pipe4_io_pipe_phv_out_data_486; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_487 = pipe4_io_pipe_phv_out_data_487; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_488 = pipe4_io_pipe_phv_out_data_488; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_489 = pipe4_io_pipe_phv_out_data_489; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_490 = pipe4_io_pipe_phv_out_data_490; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_491 = pipe4_io_pipe_phv_out_data_491; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_492 = pipe4_io_pipe_phv_out_data_492; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_493 = pipe4_io_pipe_phv_out_data_493; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_494 = pipe4_io_pipe_phv_out_data_494; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_495 = pipe4_io_pipe_phv_out_data_495; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_496 = pipe4_io_pipe_phv_out_data_496; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_497 = pipe4_io_pipe_phv_out_data_497; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_498 = pipe4_io_pipe_phv_out_data_498; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_499 = pipe4_io_pipe_phv_out_data_499; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_500 = pipe4_io_pipe_phv_out_data_500; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_501 = pipe4_io_pipe_phv_out_data_501; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_502 = pipe4_io_pipe_phv_out_data_502; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_503 = pipe4_io_pipe_phv_out_data_503; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_504 = pipe4_io_pipe_phv_out_data_504; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_505 = pipe4_io_pipe_phv_out_data_505; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_506 = pipe4_io_pipe_phv_out_data_506; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_507 = pipe4_io_pipe_phv_out_data_507; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_508 = pipe4_io_pipe_phv_out_data_508; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_509 = pipe4_io_pipe_phv_out_data_509; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_510 = pipe4_io_pipe_phv_out_data_510; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_data_511 = pipe4_io_pipe_phv_out_data_511; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_0 = pipe4_io_pipe_phv_out_header_0; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_1 = pipe4_io_pipe_phv_out_header_1; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_2 = pipe4_io_pipe_phv_out_header_2; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_3 = pipe4_io_pipe_phv_out_header_3; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_4 = pipe4_io_pipe_phv_out_header_4; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_5 = pipe4_io_pipe_phv_out_header_5; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_6 = pipe4_io_pipe_phv_out_header_6; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_7 = pipe4_io_pipe_phv_out_header_7; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_8 = pipe4_io_pipe_phv_out_header_8; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_9 = pipe4_io_pipe_phv_out_header_9; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_10 = pipe4_io_pipe_phv_out_header_10; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_11 = pipe4_io_pipe_phv_out_header_11; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_12 = pipe4_io_pipe_phv_out_header_12; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_13 = pipe4_io_pipe_phv_out_header_13; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_14 = pipe4_io_pipe_phv_out_header_14; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_header_15 = pipe4_io_pipe_phv_out_header_15; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_parse_current_state = pipe4_io_pipe_phv_out_parse_current_state; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_parse_current_offset = pipe4_io_pipe_phv_out_parse_current_offset; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_parse_transition_field = pipe4_io_pipe_phv_out_parse_transition_field; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_next_processor_id = pipe4_io_pipe_phv_out_next_processor_id; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_next_config_id = pipe4_io_pipe_phv_out_next_config_id; // @[executor.scala 517:26]
  assign pipe5_io_pipe_phv_in_is_valid_processor = pipe4_io_pipe_phv_out_is_valid_processor; // @[executor.scala 517:26]
  assign pipe5_io_vliw_in_0 = pipe4_io_vliw_out_0; // @[executor.scala 518:26]
  assign pipe5_io_vliw_in_1 = pipe4_io_vliw_out_1; // @[executor.scala 518:26]
  assign pipe5_io_vliw_in_2 = pipe4_io_vliw_out_2; // @[executor.scala 518:26]
  assign pipe5_io_vliw_in_3 = pipe4_io_vliw_out_3; // @[executor.scala 518:26]
  assign pipe5_io_field_in_0 = pipe4_io_field_out_0; // @[executor.scala 519:26]
  assign pipe5_io_field_in_1 = pipe4_io_field_out_1; // @[executor.scala 519:26]
  assign pipe5_io_field_in_2 = pipe4_io_field_out_2; // @[executor.scala 519:26]
  assign pipe5_io_field_in_3 = pipe4_io_field_out_3; // @[executor.scala 519:26]
  assign pipe5_io_mask_in_0 = pipe4_io_mask_out_0; // @[executor.scala 520:26]
  assign pipe5_io_mask_in_1 = pipe4_io_mask_out_1; // @[executor.scala 520:26]
  assign pipe5_io_mask_in_2 = pipe4_io_mask_out_2; // @[executor.scala 520:26]
  assign pipe5_io_mask_in_3 = pipe4_io_mask_out_3; // @[executor.scala 520:26]
  assign pipe5_io_bias_in_0 = pipe4_io_bias_out_0; // @[executor.scala 521:26]
  assign pipe5_io_bias_in_1 = pipe4_io_bias_out_1; // @[executor.scala 521:26]
  assign pipe5_io_bias_in_2 = pipe4_io_bias_out_2; // @[executor.scala 521:26]
  assign pipe5_io_bias_in_3 = pipe4_io_bias_out_3; // @[executor.scala 521:26]
  assign pipe5_io_dst_offset_in_0 = pipe4_io_dst_offset_out_0; // @[executor.scala 522:28]
  assign pipe5_io_dst_offset_in_1 = pipe4_io_dst_offset_out_1; // @[executor.scala 522:28]
  assign pipe5_io_dst_offset_in_2 = pipe4_io_dst_offset_out_2; // @[executor.scala 522:28]
  assign pipe5_io_dst_offset_in_3 = pipe4_io_dst_offset_out_3; // @[executor.scala 522:28]
  assign pipe6_clock = clock;
  assign pipe6_io_pipe_phv_in_data_0 = pipe5_io_pipe_phv_out_data_0; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_1 = pipe5_io_pipe_phv_out_data_1; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_2 = pipe5_io_pipe_phv_out_data_2; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_3 = pipe5_io_pipe_phv_out_data_3; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_4 = pipe5_io_pipe_phv_out_data_4; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_5 = pipe5_io_pipe_phv_out_data_5; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_6 = pipe5_io_pipe_phv_out_data_6; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_7 = pipe5_io_pipe_phv_out_data_7; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_8 = pipe5_io_pipe_phv_out_data_8; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_9 = pipe5_io_pipe_phv_out_data_9; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_10 = pipe5_io_pipe_phv_out_data_10; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_11 = pipe5_io_pipe_phv_out_data_11; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_12 = pipe5_io_pipe_phv_out_data_12; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_13 = pipe5_io_pipe_phv_out_data_13; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_14 = pipe5_io_pipe_phv_out_data_14; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_15 = pipe5_io_pipe_phv_out_data_15; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_16 = pipe5_io_pipe_phv_out_data_16; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_17 = pipe5_io_pipe_phv_out_data_17; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_18 = pipe5_io_pipe_phv_out_data_18; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_19 = pipe5_io_pipe_phv_out_data_19; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_20 = pipe5_io_pipe_phv_out_data_20; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_21 = pipe5_io_pipe_phv_out_data_21; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_22 = pipe5_io_pipe_phv_out_data_22; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_23 = pipe5_io_pipe_phv_out_data_23; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_24 = pipe5_io_pipe_phv_out_data_24; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_25 = pipe5_io_pipe_phv_out_data_25; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_26 = pipe5_io_pipe_phv_out_data_26; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_27 = pipe5_io_pipe_phv_out_data_27; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_28 = pipe5_io_pipe_phv_out_data_28; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_29 = pipe5_io_pipe_phv_out_data_29; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_30 = pipe5_io_pipe_phv_out_data_30; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_31 = pipe5_io_pipe_phv_out_data_31; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_32 = pipe5_io_pipe_phv_out_data_32; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_33 = pipe5_io_pipe_phv_out_data_33; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_34 = pipe5_io_pipe_phv_out_data_34; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_35 = pipe5_io_pipe_phv_out_data_35; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_36 = pipe5_io_pipe_phv_out_data_36; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_37 = pipe5_io_pipe_phv_out_data_37; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_38 = pipe5_io_pipe_phv_out_data_38; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_39 = pipe5_io_pipe_phv_out_data_39; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_40 = pipe5_io_pipe_phv_out_data_40; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_41 = pipe5_io_pipe_phv_out_data_41; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_42 = pipe5_io_pipe_phv_out_data_42; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_43 = pipe5_io_pipe_phv_out_data_43; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_44 = pipe5_io_pipe_phv_out_data_44; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_45 = pipe5_io_pipe_phv_out_data_45; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_46 = pipe5_io_pipe_phv_out_data_46; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_47 = pipe5_io_pipe_phv_out_data_47; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_48 = pipe5_io_pipe_phv_out_data_48; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_49 = pipe5_io_pipe_phv_out_data_49; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_50 = pipe5_io_pipe_phv_out_data_50; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_51 = pipe5_io_pipe_phv_out_data_51; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_52 = pipe5_io_pipe_phv_out_data_52; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_53 = pipe5_io_pipe_phv_out_data_53; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_54 = pipe5_io_pipe_phv_out_data_54; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_55 = pipe5_io_pipe_phv_out_data_55; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_56 = pipe5_io_pipe_phv_out_data_56; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_57 = pipe5_io_pipe_phv_out_data_57; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_58 = pipe5_io_pipe_phv_out_data_58; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_59 = pipe5_io_pipe_phv_out_data_59; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_60 = pipe5_io_pipe_phv_out_data_60; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_61 = pipe5_io_pipe_phv_out_data_61; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_62 = pipe5_io_pipe_phv_out_data_62; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_63 = pipe5_io_pipe_phv_out_data_63; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_64 = pipe5_io_pipe_phv_out_data_64; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_65 = pipe5_io_pipe_phv_out_data_65; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_66 = pipe5_io_pipe_phv_out_data_66; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_67 = pipe5_io_pipe_phv_out_data_67; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_68 = pipe5_io_pipe_phv_out_data_68; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_69 = pipe5_io_pipe_phv_out_data_69; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_70 = pipe5_io_pipe_phv_out_data_70; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_71 = pipe5_io_pipe_phv_out_data_71; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_72 = pipe5_io_pipe_phv_out_data_72; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_73 = pipe5_io_pipe_phv_out_data_73; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_74 = pipe5_io_pipe_phv_out_data_74; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_75 = pipe5_io_pipe_phv_out_data_75; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_76 = pipe5_io_pipe_phv_out_data_76; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_77 = pipe5_io_pipe_phv_out_data_77; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_78 = pipe5_io_pipe_phv_out_data_78; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_79 = pipe5_io_pipe_phv_out_data_79; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_80 = pipe5_io_pipe_phv_out_data_80; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_81 = pipe5_io_pipe_phv_out_data_81; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_82 = pipe5_io_pipe_phv_out_data_82; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_83 = pipe5_io_pipe_phv_out_data_83; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_84 = pipe5_io_pipe_phv_out_data_84; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_85 = pipe5_io_pipe_phv_out_data_85; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_86 = pipe5_io_pipe_phv_out_data_86; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_87 = pipe5_io_pipe_phv_out_data_87; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_88 = pipe5_io_pipe_phv_out_data_88; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_89 = pipe5_io_pipe_phv_out_data_89; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_90 = pipe5_io_pipe_phv_out_data_90; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_91 = pipe5_io_pipe_phv_out_data_91; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_92 = pipe5_io_pipe_phv_out_data_92; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_93 = pipe5_io_pipe_phv_out_data_93; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_94 = pipe5_io_pipe_phv_out_data_94; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_95 = pipe5_io_pipe_phv_out_data_95; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_96 = pipe5_io_pipe_phv_out_data_96; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_97 = pipe5_io_pipe_phv_out_data_97; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_98 = pipe5_io_pipe_phv_out_data_98; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_99 = pipe5_io_pipe_phv_out_data_99; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_100 = pipe5_io_pipe_phv_out_data_100; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_101 = pipe5_io_pipe_phv_out_data_101; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_102 = pipe5_io_pipe_phv_out_data_102; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_103 = pipe5_io_pipe_phv_out_data_103; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_104 = pipe5_io_pipe_phv_out_data_104; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_105 = pipe5_io_pipe_phv_out_data_105; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_106 = pipe5_io_pipe_phv_out_data_106; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_107 = pipe5_io_pipe_phv_out_data_107; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_108 = pipe5_io_pipe_phv_out_data_108; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_109 = pipe5_io_pipe_phv_out_data_109; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_110 = pipe5_io_pipe_phv_out_data_110; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_111 = pipe5_io_pipe_phv_out_data_111; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_112 = pipe5_io_pipe_phv_out_data_112; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_113 = pipe5_io_pipe_phv_out_data_113; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_114 = pipe5_io_pipe_phv_out_data_114; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_115 = pipe5_io_pipe_phv_out_data_115; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_116 = pipe5_io_pipe_phv_out_data_116; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_117 = pipe5_io_pipe_phv_out_data_117; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_118 = pipe5_io_pipe_phv_out_data_118; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_119 = pipe5_io_pipe_phv_out_data_119; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_120 = pipe5_io_pipe_phv_out_data_120; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_121 = pipe5_io_pipe_phv_out_data_121; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_122 = pipe5_io_pipe_phv_out_data_122; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_123 = pipe5_io_pipe_phv_out_data_123; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_124 = pipe5_io_pipe_phv_out_data_124; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_125 = pipe5_io_pipe_phv_out_data_125; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_126 = pipe5_io_pipe_phv_out_data_126; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_127 = pipe5_io_pipe_phv_out_data_127; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_128 = pipe5_io_pipe_phv_out_data_128; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_129 = pipe5_io_pipe_phv_out_data_129; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_130 = pipe5_io_pipe_phv_out_data_130; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_131 = pipe5_io_pipe_phv_out_data_131; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_132 = pipe5_io_pipe_phv_out_data_132; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_133 = pipe5_io_pipe_phv_out_data_133; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_134 = pipe5_io_pipe_phv_out_data_134; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_135 = pipe5_io_pipe_phv_out_data_135; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_136 = pipe5_io_pipe_phv_out_data_136; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_137 = pipe5_io_pipe_phv_out_data_137; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_138 = pipe5_io_pipe_phv_out_data_138; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_139 = pipe5_io_pipe_phv_out_data_139; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_140 = pipe5_io_pipe_phv_out_data_140; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_141 = pipe5_io_pipe_phv_out_data_141; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_142 = pipe5_io_pipe_phv_out_data_142; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_143 = pipe5_io_pipe_phv_out_data_143; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_144 = pipe5_io_pipe_phv_out_data_144; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_145 = pipe5_io_pipe_phv_out_data_145; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_146 = pipe5_io_pipe_phv_out_data_146; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_147 = pipe5_io_pipe_phv_out_data_147; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_148 = pipe5_io_pipe_phv_out_data_148; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_149 = pipe5_io_pipe_phv_out_data_149; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_150 = pipe5_io_pipe_phv_out_data_150; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_151 = pipe5_io_pipe_phv_out_data_151; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_152 = pipe5_io_pipe_phv_out_data_152; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_153 = pipe5_io_pipe_phv_out_data_153; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_154 = pipe5_io_pipe_phv_out_data_154; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_155 = pipe5_io_pipe_phv_out_data_155; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_156 = pipe5_io_pipe_phv_out_data_156; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_157 = pipe5_io_pipe_phv_out_data_157; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_158 = pipe5_io_pipe_phv_out_data_158; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_159 = pipe5_io_pipe_phv_out_data_159; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_160 = pipe5_io_pipe_phv_out_data_160; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_161 = pipe5_io_pipe_phv_out_data_161; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_162 = pipe5_io_pipe_phv_out_data_162; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_163 = pipe5_io_pipe_phv_out_data_163; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_164 = pipe5_io_pipe_phv_out_data_164; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_165 = pipe5_io_pipe_phv_out_data_165; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_166 = pipe5_io_pipe_phv_out_data_166; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_167 = pipe5_io_pipe_phv_out_data_167; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_168 = pipe5_io_pipe_phv_out_data_168; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_169 = pipe5_io_pipe_phv_out_data_169; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_170 = pipe5_io_pipe_phv_out_data_170; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_171 = pipe5_io_pipe_phv_out_data_171; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_172 = pipe5_io_pipe_phv_out_data_172; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_173 = pipe5_io_pipe_phv_out_data_173; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_174 = pipe5_io_pipe_phv_out_data_174; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_175 = pipe5_io_pipe_phv_out_data_175; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_176 = pipe5_io_pipe_phv_out_data_176; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_177 = pipe5_io_pipe_phv_out_data_177; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_178 = pipe5_io_pipe_phv_out_data_178; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_179 = pipe5_io_pipe_phv_out_data_179; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_180 = pipe5_io_pipe_phv_out_data_180; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_181 = pipe5_io_pipe_phv_out_data_181; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_182 = pipe5_io_pipe_phv_out_data_182; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_183 = pipe5_io_pipe_phv_out_data_183; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_184 = pipe5_io_pipe_phv_out_data_184; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_185 = pipe5_io_pipe_phv_out_data_185; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_186 = pipe5_io_pipe_phv_out_data_186; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_187 = pipe5_io_pipe_phv_out_data_187; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_188 = pipe5_io_pipe_phv_out_data_188; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_189 = pipe5_io_pipe_phv_out_data_189; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_190 = pipe5_io_pipe_phv_out_data_190; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_191 = pipe5_io_pipe_phv_out_data_191; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_192 = pipe5_io_pipe_phv_out_data_192; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_193 = pipe5_io_pipe_phv_out_data_193; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_194 = pipe5_io_pipe_phv_out_data_194; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_195 = pipe5_io_pipe_phv_out_data_195; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_196 = pipe5_io_pipe_phv_out_data_196; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_197 = pipe5_io_pipe_phv_out_data_197; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_198 = pipe5_io_pipe_phv_out_data_198; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_199 = pipe5_io_pipe_phv_out_data_199; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_200 = pipe5_io_pipe_phv_out_data_200; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_201 = pipe5_io_pipe_phv_out_data_201; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_202 = pipe5_io_pipe_phv_out_data_202; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_203 = pipe5_io_pipe_phv_out_data_203; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_204 = pipe5_io_pipe_phv_out_data_204; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_205 = pipe5_io_pipe_phv_out_data_205; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_206 = pipe5_io_pipe_phv_out_data_206; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_207 = pipe5_io_pipe_phv_out_data_207; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_208 = pipe5_io_pipe_phv_out_data_208; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_209 = pipe5_io_pipe_phv_out_data_209; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_210 = pipe5_io_pipe_phv_out_data_210; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_211 = pipe5_io_pipe_phv_out_data_211; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_212 = pipe5_io_pipe_phv_out_data_212; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_213 = pipe5_io_pipe_phv_out_data_213; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_214 = pipe5_io_pipe_phv_out_data_214; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_215 = pipe5_io_pipe_phv_out_data_215; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_216 = pipe5_io_pipe_phv_out_data_216; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_217 = pipe5_io_pipe_phv_out_data_217; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_218 = pipe5_io_pipe_phv_out_data_218; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_219 = pipe5_io_pipe_phv_out_data_219; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_220 = pipe5_io_pipe_phv_out_data_220; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_221 = pipe5_io_pipe_phv_out_data_221; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_222 = pipe5_io_pipe_phv_out_data_222; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_223 = pipe5_io_pipe_phv_out_data_223; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_224 = pipe5_io_pipe_phv_out_data_224; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_225 = pipe5_io_pipe_phv_out_data_225; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_226 = pipe5_io_pipe_phv_out_data_226; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_227 = pipe5_io_pipe_phv_out_data_227; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_228 = pipe5_io_pipe_phv_out_data_228; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_229 = pipe5_io_pipe_phv_out_data_229; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_230 = pipe5_io_pipe_phv_out_data_230; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_231 = pipe5_io_pipe_phv_out_data_231; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_232 = pipe5_io_pipe_phv_out_data_232; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_233 = pipe5_io_pipe_phv_out_data_233; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_234 = pipe5_io_pipe_phv_out_data_234; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_235 = pipe5_io_pipe_phv_out_data_235; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_236 = pipe5_io_pipe_phv_out_data_236; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_237 = pipe5_io_pipe_phv_out_data_237; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_238 = pipe5_io_pipe_phv_out_data_238; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_239 = pipe5_io_pipe_phv_out_data_239; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_240 = pipe5_io_pipe_phv_out_data_240; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_241 = pipe5_io_pipe_phv_out_data_241; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_242 = pipe5_io_pipe_phv_out_data_242; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_243 = pipe5_io_pipe_phv_out_data_243; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_244 = pipe5_io_pipe_phv_out_data_244; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_245 = pipe5_io_pipe_phv_out_data_245; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_246 = pipe5_io_pipe_phv_out_data_246; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_247 = pipe5_io_pipe_phv_out_data_247; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_248 = pipe5_io_pipe_phv_out_data_248; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_249 = pipe5_io_pipe_phv_out_data_249; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_250 = pipe5_io_pipe_phv_out_data_250; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_251 = pipe5_io_pipe_phv_out_data_251; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_252 = pipe5_io_pipe_phv_out_data_252; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_253 = pipe5_io_pipe_phv_out_data_253; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_254 = pipe5_io_pipe_phv_out_data_254; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_255 = pipe5_io_pipe_phv_out_data_255; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_256 = pipe5_io_pipe_phv_out_data_256; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_257 = pipe5_io_pipe_phv_out_data_257; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_258 = pipe5_io_pipe_phv_out_data_258; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_259 = pipe5_io_pipe_phv_out_data_259; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_260 = pipe5_io_pipe_phv_out_data_260; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_261 = pipe5_io_pipe_phv_out_data_261; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_262 = pipe5_io_pipe_phv_out_data_262; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_263 = pipe5_io_pipe_phv_out_data_263; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_264 = pipe5_io_pipe_phv_out_data_264; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_265 = pipe5_io_pipe_phv_out_data_265; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_266 = pipe5_io_pipe_phv_out_data_266; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_267 = pipe5_io_pipe_phv_out_data_267; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_268 = pipe5_io_pipe_phv_out_data_268; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_269 = pipe5_io_pipe_phv_out_data_269; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_270 = pipe5_io_pipe_phv_out_data_270; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_271 = pipe5_io_pipe_phv_out_data_271; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_272 = pipe5_io_pipe_phv_out_data_272; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_273 = pipe5_io_pipe_phv_out_data_273; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_274 = pipe5_io_pipe_phv_out_data_274; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_275 = pipe5_io_pipe_phv_out_data_275; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_276 = pipe5_io_pipe_phv_out_data_276; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_277 = pipe5_io_pipe_phv_out_data_277; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_278 = pipe5_io_pipe_phv_out_data_278; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_279 = pipe5_io_pipe_phv_out_data_279; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_280 = pipe5_io_pipe_phv_out_data_280; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_281 = pipe5_io_pipe_phv_out_data_281; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_282 = pipe5_io_pipe_phv_out_data_282; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_283 = pipe5_io_pipe_phv_out_data_283; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_284 = pipe5_io_pipe_phv_out_data_284; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_285 = pipe5_io_pipe_phv_out_data_285; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_286 = pipe5_io_pipe_phv_out_data_286; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_287 = pipe5_io_pipe_phv_out_data_287; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_288 = pipe5_io_pipe_phv_out_data_288; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_289 = pipe5_io_pipe_phv_out_data_289; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_290 = pipe5_io_pipe_phv_out_data_290; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_291 = pipe5_io_pipe_phv_out_data_291; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_292 = pipe5_io_pipe_phv_out_data_292; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_293 = pipe5_io_pipe_phv_out_data_293; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_294 = pipe5_io_pipe_phv_out_data_294; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_295 = pipe5_io_pipe_phv_out_data_295; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_296 = pipe5_io_pipe_phv_out_data_296; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_297 = pipe5_io_pipe_phv_out_data_297; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_298 = pipe5_io_pipe_phv_out_data_298; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_299 = pipe5_io_pipe_phv_out_data_299; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_300 = pipe5_io_pipe_phv_out_data_300; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_301 = pipe5_io_pipe_phv_out_data_301; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_302 = pipe5_io_pipe_phv_out_data_302; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_303 = pipe5_io_pipe_phv_out_data_303; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_304 = pipe5_io_pipe_phv_out_data_304; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_305 = pipe5_io_pipe_phv_out_data_305; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_306 = pipe5_io_pipe_phv_out_data_306; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_307 = pipe5_io_pipe_phv_out_data_307; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_308 = pipe5_io_pipe_phv_out_data_308; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_309 = pipe5_io_pipe_phv_out_data_309; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_310 = pipe5_io_pipe_phv_out_data_310; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_311 = pipe5_io_pipe_phv_out_data_311; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_312 = pipe5_io_pipe_phv_out_data_312; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_313 = pipe5_io_pipe_phv_out_data_313; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_314 = pipe5_io_pipe_phv_out_data_314; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_315 = pipe5_io_pipe_phv_out_data_315; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_316 = pipe5_io_pipe_phv_out_data_316; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_317 = pipe5_io_pipe_phv_out_data_317; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_318 = pipe5_io_pipe_phv_out_data_318; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_319 = pipe5_io_pipe_phv_out_data_319; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_320 = pipe5_io_pipe_phv_out_data_320; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_321 = pipe5_io_pipe_phv_out_data_321; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_322 = pipe5_io_pipe_phv_out_data_322; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_323 = pipe5_io_pipe_phv_out_data_323; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_324 = pipe5_io_pipe_phv_out_data_324; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_325 = pipe5_io_pipe_phv_out_data_325; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_326 = pipe5_io_pipe_phv_out_data_326; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_327 = pipe5_io_pipe_phv_out_data_327; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_328 = pipe5_io_pipe_phv_out_data_328; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_329 = pipe5_io_pipe_phv_out_data_329; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_330 = pipe5_io_pipe_phv_out_data_330; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_331 = pipe5_io_pipe_phv_out_data_331; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_332 = pipe5_io_pipe_phv_out_data_332; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_333 = pipe5_io_pipe_phv_out_data_333; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_334 = pipe5_io_pipe_phv_out_data_334; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_335 = pipe5_io_pipe_phv_out_data_335; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_336 = pipe5_io_pipe_phv_out_data_336; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_337 = pipe5_io_pipe_phv_out_data_337; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_338 = pipe5_io_pipe_phv_out_data_338; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_339 = pipe5_io_pipe_phv_out_data_339; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_340 = pipe5_io_pipe_phv_out_data_340; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_341 = pipe5_io_pipe_phv_out_data_341; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_342 = pipe5_io_pipe_phv_out_data_342; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_343 = pipe5_io_pipe_phv_out_data_343; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_344 = pipe5_io_pipe_phv_out_data_344; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_345 = pipe5_io_pipe_phv_out_data_345; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_346 = pipe5_io_pipe_phv_out_data_346; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_347 = pipe5_io_pipe_phv_out_data_347; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_348 = pipe5_io_pipe_phv_out_data_348; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_349 = pipe5_io_pipe_phv_out_data_349; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_350 = pipe5_io_pipe_phv_out_data_350; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_351 = pipe5_io_pipe_phv_out_data_351; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_352 = pipe5_io_pipe_phv_out_data_352; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_353 = pipe5_io_pipe_phv_out_data_353; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_354 = pipe5_io_pipe_phv_out_data_354; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_355 = pipe5_io_pipe_phv_out_data_355; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_356 = pipe5_io_pipe_phv_out_data_356; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_357 = pipe5_io_pipe_phv_out_data_357; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_358 = pipe5_io_pipe_phv_out_data_358; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_359 = pipe5_io_pipe_phv_out_data_359; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_360 = pipe5_io_pipe_phv_out_data_360; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_361 = pipe5_io_pipe_phv_out_data_361; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_362 = pipe5_io_pipe_phv_out_data_362; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_363 = pipe5_io_pipe_phv_out_data_363; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_364 = pipe5_io_pipe_phv_out_data_364; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_365 = pipe5_io_pipe_phv_out_data_365; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_366 = pipe5_io_pipe_phv_out_data_366; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_367 = pipe5_io_pipe_phv_out_data_367; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_368 = pipe5_io_pipe_phv_out_data_368; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_369 = pipe5_io_pipe_phv_out_data_369; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_370 = pipe5_io_pipe_phv_out_data_370; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_371 = pipe5_io_pipe_phv_out_data_371; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_372 = pipe5_io_pipe_phv_out_data_372; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_373 = pipe5_io_pipe_phv_out_data_373; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_374 = pipe5_io_pipe_phv_out_data_374; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_375 = pipe5_io_pipe_phv_out_data_375; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_376 = pipe5_io_pipe_phv_out_data_376; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_377 = pipe5_io_pipe_phv_out_data_377; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_378 = pipe5_io_pipe_phv_out_data_378; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_379 = pipe5_io_pipe_phv_out_data_379; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_380 = pipe5_io_pipe_phv_out_data_380; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_381 = pipe5_io_pipe_phv_out_data_381; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_382 = pipe5_io_pipe_phv_out_data_382; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_383 = pipe5_io_pipe_phv_out_data_383; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_384 = pipe5_io_pipe_phv_out_data_384; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_385 = pipe5_io_pipe_phv_out_data_385; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_386 = pipe5_io_pipe_phv_out_data_386; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_387 = pipe5_io_pipe_phv_out_data_387; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_388 = pipe5_io_pipe_phv_out_data_388; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_389 = pipe5_io_pipe_phv_out_data_389; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_390 = pipe5_io_pipe_phv_out_data_390; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_391 = pipe5_io_pipe_phv_out_data_391; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_392 = pipe5_io_pipe_phv_out_data_392; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_393 = pipe5_io_pipe_phv_out_data_393; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_394 = pipe5_io_pipe_phv_out_data_394; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_395 = pipe5_io_pipe_phv_out_data_395; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_396 = pipe5_io_pipe_phv_out_data_396; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_397 = pipe5_io_pipe_phv_out_data_397; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_398 = pipe5_io_pipe_phv_out_data_398; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_399 = pipe5_io_pipe_phv_out_data_399; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_400 = pipe5_io_pipe_phv_out_data_400; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_401 = pipe5_io_pipe_phv_out_data_401; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_402 = pipe5_io_pipe_phv_out_data_402; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_403 = pipe5_io_pipe_phv_out_data_403; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_404 = pipe5_io_pipe_phv_out_data_404; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_405 = pipe5_io_pipe_phv_out_data_405; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_406 = pipe5_io_pipe_phv_out_data_406; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_407 = pipe5_io_pipe_phv_out_data_407; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_408 = pipe5_io_pipe_phv_out_data_408; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_409 = pipe5_io_pipe_phv_out_data_409; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_410 = pipe5_io_pipe_phv_out_data_410; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_411 = pipe5_io_pipe_phv_out_data_411; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_412 = pipe5_io_pipe_phv_out_data_412; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_413 = pipe5_io_pipe_phv_out_data_413; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_414 = pipe5_io_pipe_phv_out_data_414; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_415 = pipe5_io_pipe_phv_out_data_415; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_416 = pipe5_io_pipe_phv_out_data_416; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_417 = pipe5_io_pipe_phv_out_data_417; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_418 = pipe5_io_pipe_phv_out_data_418; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_419 = pipe5_io_pipe_phv_out_data_419; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_420 = pipe5_io_pipe_phv_out_data_420; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_421 = pipe5_io_pipe_phv_out_data_421; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_422 = pipe5_io_pipe_phv_out_data_422; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_423 = pipe5_io_pipe_phv_out_data_423; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_424 = pipe5_io_pipe_phv_out_data_424; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_425 = pipe5_io_pipe_phv_out_data_425; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_426 = pipe5_io_pipe_phv_out_data_426; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_427 = pipe5_io_pipe_phv_out_data_427; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_428 = pipe5_io_pipe_phv_out_data_428; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_429 = pipe5_io_pipe_phv_out_data_429; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_430 = pipe5_io_pipe_phv_out_data_430; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_431 = pipe5_io_pipe_phv_out_data_431; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_432 = pipe5_io_pipe_phv_out_data_432; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_433 = pipe5_io_pipe_phv_out_data_433; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_434 = pipe5_io_pipe_phv_out_data_434; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_435 = pipe5_io_pipe_phv_out_data_435; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_436 = pipe5_io_pipe_phv_out_data_436; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_437 = pipe5_io_pipe_phv_out_data_437; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_438 = pipe5_io_pipe_phv_out_data_438; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_439 = pipe5_io_pipe_phv_out_data_439; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_440 = pipe5_io_pipe_phv_out_data_440; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_441 = pipe5_io_pipe_phv_out_data_441; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_442 = pipe5_io_pipe_phv_out_data_442; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_443 = pipe5_io_pipe_phv_out_data_443; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_444 = pipe5_io_pipe_phv_out_data_444; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_445 = pipe5_io_pipe_phv_out_data_445; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_446 = pipe5_io_pipe_phv_out_data_446; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_447 = pipe5_io_pipe_phv_out_data_447; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_448 = pipe5_io_pipe_phv_out_data_448; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_449 = pipe5_io_pipe_phv_out_data_449; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_450 = pipe5_io_pipe_phv_out_data_450; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_451 = pipe5_io_pipe_phv_out_data_451; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_452 = pipe5_io_pipe_phv_out_data_452; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_453 = pipe5_io_pipe_phv_out_data_453; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_454 = pipe5_io_pipe_phv_out_data_454; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_455 = pipe5_io_pipe_phv_out_data_455; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_456 = pipe5_io_pipe_phv_out_data_456; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_457 = pipe5_io_pipe_phv_out_data_457; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_458 = pipe5_io_pipe_phv_out_data_458; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_459 = pipe5_io_pipe_phv_out_data_459; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_460 = pipe5_io_pipe_phv_out_data_460; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_461 = pipe5_io_pipe_phv_out_data_461; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_462 = pipe5_io_pipe_phv_out_data_462; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_463 = pipe5_io_pipe_phv_out_data_463; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_464 = pipe5_io_pipe_phv_out_data_464; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_465 = pipe5_io_pipe_phv_out_data_465; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_466 = pipe5_io_pipe_phv_out_data_466; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_467 = pipe5_io_pipe_phv_out_data_467; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_468 = pipe5_io_pipe_phv_out_data_468; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_469 = pipe5_io_pipe_phv_out_data_469; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_470 = pipe5_io_pipe_phv_out_data_470; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_471 = pipe5_io_pipe_phv_out_data_471; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_472 = pipe5_io_pipe_phv_out_data_472; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_473 = pipe5_io_pipe_phv_out_data_473; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_474 = pipe5_io_pipe_phv_out_data_474; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_475 = pipe5_io_pipe_phv_out_data_475; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_476 = pipe5_io_pipe_phv_out_data_476; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_477 = pipe5_io_pipe_phv_out_data_477; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_478 = pipe5_io_pipe_phv_out_data_478; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_479 = pipe5_io_pipe_phv_out_data_479; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_480 = pipe5_io_pipe_phv_out_data_480; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_481 = pipe5_io_pipe_phv_out_data_481; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_482 = pipe5_io_pipe_phv_out_data_482; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_483 = pipe5_io_pipe_phv_out_data_483; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_484 = pipe5_io_pipe_phv_out_data_484; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_485 = pipe5_io_pipe_phv_out_data_485; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_486 = pipe5_io_pipe_phv_out_data_486; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_487 = pipe5_io_pipe_phv_out_data_487; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_488 = pipe5_io_pipe_phv_out_data_488; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_489 = pipe5_io_pipe_phv_out_data_489; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_490 = pipe5_io_pipe_phv_out_data_490; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_491 = pipe5_io_pipe_phv_out_data_491; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_492 = pipe5_io_pipe_phv_out_data_492; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_493 = pipe5_io_pipe_phv_out_data_493; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_494 = pipe5_io_pipe_phv_out_data_494; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_495 = pipe5_io_pipe_phv_out_data_495; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_496 = pipe5_io_pipe_phv_out_data_496; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_497 = pipe5_io_pipe_phv_out_data_497; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_498 = pipe5_io_pipe_phv_out_data_498; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_499 = pipe5_io_pipe_phv_out_data_499; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_500 = pipe5_io_pipe_phv_out_data_500; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_501 = pipe5_io_pipe_phv_out_data_501; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_502 = pipe5_io_pipe_phv_out_data_502; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_503 = pipe5_io_pipe_phv_out_data_503; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_504 = pipe5_io_pipe_phv_out_data_504; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_505 = pipe5_io_pipe_phv_out_data_505; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_506 = pipe5_io_pipe_phv_out_data_506; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_507 = pipe5_io_pipe_phv_out_data_507; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_508 = pipe5_io_pipe_phv_out_data_508; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_509 = pipe5_io_pipe_phv_out_data_509; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_510 = pipe5_io_pipe_phv_out_data_510; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_data_511 = pipe5_io_pipe_phv_out_data_511; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_0 = pipe5_io_pipe_phv_out_header_0; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_1 = pipe5_io_pipe_phv_out_header_1; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_2 = pipe5_io_pipe_phv_out_header_2; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_3 = pipe5_io_pipe_phv_out_header_3; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_4 = pipe5_io_pipe_phv_out_header_4; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_5 = pipe5_io_pipe_phv_out_header_5; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_6 = pipe5_io_pipe_phv_out_header_6; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_7 = pipe5_io_pipe_phv_out_header_7; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_8 = pipe5_io_pipe_phv_out_header_8; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_9 = pipe5_io_pipe_phv_out_header_9; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_10 = pipe5_io_pipe_phv_out_header_10; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_11 = pipe5_io_pipe_phv_out_header_11; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_12 = pipe5_io_pipe_phv_out_header_12; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_13 = pipe5_io_pipe_phv_out_header_13; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_14 = pipe5_io_pipe_phv_out_header_14; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_header_15 = pipe5_io_pipe_phv_out_header_15; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_parse_current_state = pipe5_io_pipe_phv_out_parse_current_state; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_parse_current_offset = pipe5_io_pipe_phv_out_parse_current_offset; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_parse_transition_field = pipe5_io_pipe_phv_out_parse_transition_field; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_next_processor_id = pipe5_io_pipe_phv_out_next_processor_id; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_next_config_id = pipe5_io_pipe_phv_out_next_config_id; // @[executor.scala 524:26]
  assign pipe6_io_pipe_phv_in_is_valid_processor = pipe5_io_pipe_phv_out_is_valid_processor; // @[executor.scala 524:26]
  assign pipe6_io_vliw_in_0 = pipe5_io_vliw_out_0; // @[executor.scala 525:26]
  assign pipe6_io_vliw_in_1 = pipe5_io_vliw_out_1; // @[executor.scala 525:26]
  assign pipe6_io_vliw_in_2 = pipe5_io_vliw_out_2; // @[executor.scala 525:26]
  assign pipe6_io_vliw_in_3 = pipe5_io_vliw_out_3; // @[executor.scala 525:26]
  assign pipe6_io_field_in_0 = pipe5_io_field_out_0; // @[executor.scala 526:26]
  assign pipe6_io_field_in_1 = pipe5_io_field_out_1; // @[executor.scala 526:26]
  assign pipe6_io_field_in_2 = pipe5_io_field_out_2; // @[executor.scala 526:26]
  assign pipe6_io_field_in_3 = pipe5_io_field_out_3; // @[executor.scala 526:26]
  assign pipe6_io_mask_in_0 = pipe5_io_mask_out_0; // @[executor.scala 527:26]
  assign pipe6_io_mask_in_1 = pipe5_io_mask_out_1; // @[executor.scala 527:26]
  assign pipe6_io_mask_in_2 = pipe5_io_mask_out_2; // @[executor.scala 527:26]
  assign pipe6_io_mask_in_3 = pipe5_io_mask_out_3; // @[executor.scala 527:26]
  assign pipe6_io_dst_offset_in_0 = pipe5_io_dst_offset_out_0; // @[executor.scala 528:28]
  assign pipe6_io_dst_offset_in_1 = pipe5_io_dst_offset_out_1; // @[executor.scala 528:28]
  assign pipe6_io_dst_offset_in_2 = pipe5_io_dst_offset_out_2; // @[executor.scala 528:28]
  assign pipe6_io_dst_offset_in_3 = pipe5_io_dst_offset_out_3; // @[executor.scala 528:28]
endmodule
